`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CPn2I7daMOzItXm7j1790g307K6Yt5pMCMq2gFTK6TWPH/ZCgmcYzKDh0OPB2sof1fOvV/L3GNPa
e+NeTQIdnQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XEyadwQlZVZDQz58rBwoYtrEJbuiVzcvx7utG8/V6HHIVBXjppJrhJ++Mx9FyhPioR2ZWmc/JopB
eqWsi/SxMVFjgPKe+2HPp8+IgJoPUB/AGQLIhrfziikFMRJ98TflqbdFI18QMQq2TDNSQZm1HXSs
/8e45G+lfb3IRc/5vhk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HWbHLMENc4OlrcumquBeAzrrc5NxXEFu+/K38d1FtWtJaBkmwWp/VZDDeNnZuiS5WD5ap4DKyU5+
m8R+vhqY6YRIjl48Kx1+5i2z6frEHdSRdCZjfEPkB9B2L7A8pvyS9/YyWL1vdDc//YDOCBz1zMCD
nJsdH9uKFdwbmiAxG4soYmQ7r1KWxVsZMOtX4bheD+fy9IkcjhPd1iZlC1iH975LThUkBw9eu+Qp
BJ+7kBSSqTFc38f2yS0umi6umNwpDq/jU1ovHlyp/pXwmFZwg0ov1Zvxc4gi0yHEtBnXaSklxXDF
Hb0FZlgAgCSKoTqUPczKmE76JH9NEGOrxxTH6g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YgAVLyEpHxfYCuul1W3qErkqxVZmzQD1JfSViVpa33W39pYP5H1d2EZp/YoO671Pcr0OHtYjq6gh
0vqRu5QJ+eW4oFnkbQmqLIWgXbBRi8OjDoZctCw9JB9O6sGi70eJy/idfMIcrnQyGSjfjaBUcKJ3
idJ7/2oXcgUBumYSdBTDg9f394SpXZjZnfi7WNTBxFTHTwySMYoT/BdYKWzAlpcvnhvGm2TuIUrR
kYnQ6VRdATLSk76P31pf8b7wPv9fW7+y5W5wsmRnjkeY9WsFvzy52Og+8TGPNWIXDBgyrhXkQ1uc
iAGGtp3qdJ1vXfQO2+stF/t9twP66uJv63hU5A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LK8Y9agL7deL0rWLeZpe9CTnMl/nD/BCX7vzQUQ9T3bt3P6yr26pebmSshl9Lwt/Xok4IGSCyMHV
VnOOeyHaZHvKsYBeD1Egn7pZ1V66aXhzXzaoKL/A7h0m9680xq3duJhz1KT3QpxnQe9EhtOvpeOi
FcjjOdsMtwvx5a7PJTgLYnLqG9ul4NbzkJzU8BMj9f0u5k2ajognJ0slOHN2EyOAIMhdw8Ead8J8
y591pJtRZTxu5ZLONzv9mFLOryH3AEBrctJu05PqzUZ3uj+3yGYqRm/K6fA40HC0urNlj1L5G28h
hcD5fsTOsx/SWpkFEzsaPWX4gdsKL2ufi8lWZA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CO7gH/890LuOMaBYzwXTF8Z+4q/08Hd2Z6bHo3hUab7ak07zXpU+iDHgxck7iMmmsk7o6ZqFlyAP
F04kDiP1ll6s35aw2YJnPxE8A+OMJEiJEII4L22offm5wtttzAw4ajmqXOfdTJr25HgmVrnhP85U
wE8Jwh97mnNgPa25RI0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CEvFR3i951wRDLIlqQnkCMH9+k+npBmQSlTonlqasYMOYGTlpiRZ89TxNR3uXFrBvzInIJ+lI5CM
2IH4iqDiJanGDlnns2fXzD+8OERjePv4Tokb+8CiEFQ0UShldf5PuVRbGgxEZzblc0zU5IYIp/Px
ttvCoPc3o2rhHibcVppeeWDgUJJ5alBq9rOtzfN/wzn7iCrc7AnR2W0cRKoDhuROp5XgCglweg+2
CxaggvdhNR3lt2CK+WCO0i9HDSx4hkF8/WIkZkwfE12pdeBiOcZuz1T39Tj12eG7i6QsfgGJU+YT
yRgl8ag9MQzUnOBoAmI3RgTtJk4q+EqtdwqIBg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211312)
`protect data_block
rvQ5x0gCrZlGQmNKzc0g0jCeua7KOeaKWu0KVH08xd0fNBg8dCk6wIlKC41DTqQtkNWYRqoRZTi+
Ke77MJj+65GsM1SBvKvj2EfG2fhsdyXGf2fIcaSOst6HTYrxy5KupSwkP6h6Xwwml7MVH0JgroKa
g09QlAQJ0NI0UlR4Y5e+jWx2Y2f4/mxMzVAlylju0A+OMHnpyRBt3zhS1DPm2t2kX2xJ26HsYppM
CKXedU/p6eVICYzCY7pnaZNIXJowNpHx/C6NhlQSLUW68wiw3AtpCN35vLchPkN/8rV/e/gMaqzf
T2pZXA3dBoIfFXEkikw0KrmytK9EHA7NmySYAZuMGAQ8H+rdbBAZWWMzh3hpFUhkT0Pcgf39VvVU
tmLx3PVsM7U9wq4miI7MyBaV9CB9lRplKFvoq9i2Npau5Jd6K9uQHCdNY+RnCDyvWlLmGuunIGQ8
rSgITSkGytleveE5kCaVwqZQymsK9BrhWQnJR6UXzl9cloAJws8a7d74hXOJJ7eljIIC8oKP7aiz
zki1yDBtsKxaKtlqUcOW1aL0wp5JKwpOZjxVFs56s7zM138y4u8Bm7M7Qj643mzuV0qRSPWjrAi9
qkQVmNgDtduoryMjBBnCpFeyLKhVTo2U2iNiIJHlrIPe6t48kqew4gKhtj5MPUeUXBAsCiJAg8XD
zDytot3+eQAi6z2LrvLGCo2s0l5O5mSOw2q/DZkk0BDgmPRTeFapTc58NyojHP2oCp0lcDlF0JdG
VEQUQtWHMj+XMvsj71GjJ39BfBjAkfmgPgGXEqiXRf+1JAznUZiWqVuvzAv1w27/bQJjAzlgidrC
N0tEC+0JcR9Lkf78vFFPawGJCbuCImzltcJ56CcjV+rdJMp4BDx5r+S5DBWJk1dSj6Zaksakzmqw
nsbt5ATHy60RmPMBy4PFb70Db03REGC5bMQT64udVZkX4DMOpvMBJIV9HDQeyjHoWsI3aWuG7MOk
cma0JjxkY1l6BwSowGzXfzJb708gG6T31T0HJEAAx+NXXjMAP0SJaq8E8l6RIiDIIncJwSGRBUe3
La5R2Ha83dvyalpVftNnMvGrLtkblUaVNEbUg11TeiJIIHeR9Xgp8impcY98nRe9VhstBHzK1wS+
PVAGuaBI6W3FfWp86uuDlvQYbCFfGlPnv0Dh0TXA17S7q2TWO0HGKKrlhHzXjD5uwuvLBBu73E/7
r1AnPUqChMD7FV54R3m1pE7iHOEzn0x8y9CYL+J+D0QinaVlPS65LUFmdNeNZZNpyGgnri3rT+Cv
PF/OgaS9/zddZEQnn92NlBlZGw8AZOSUvIwKIlXadXme4r47/dwd8AFNohE2aw5ZZ6vzZgH4MtVi
GpDiBeRnA5eVIRMH0iEAb5DPvWg1vMZOmk2N0wkeBvVp/oY66tedENA4ygL4CP7VSZLqjQ8tsc8I
kIIkcbekG09vYYjPYE8MYWTsjFp9REzgnza4IsknOnFCL15t+f5/rnsnMNZEMMfjOuC+CxN5pW+h
GSFWWBjjqcGukfzVJMYwNZFp/GxayM5PEb3Mbyh2MHvhnpOv+NsPgqrG9DFJHRoIero+nDOcdQMb
SzRFzy0++CbqF83nAfgRRJ5i52E7knQsoVmUGn2Zw2TfxQRkdMLpG2qJpTqrt0jNYODak9WeYbyX
Gw22xHuxbIR8xgZuQgeQ/YkAXa15IPdmswstsROh33vTMNPMQEopijlDyy8Sr8zFZ0fpHTM5fWbA
LFGE+3Q3Lexu2dH3Mj3axjMU0O4mctBzjGQfVripSB1YtarEKrEiwQBXd9TOkq+P3PErTKwSyK1Y
xoNdDPGvuwCghULX/fPRlX8jTWMZidZ66uJdEXmkmTbeLcKbFIJz7dF122xz+ggHS2q5NYKsE8hu
KjeYMXL/FYkt3Zv+IKgmw327ShZBxyOjkt6ALZSO0RRXr3LyQqfTiqtZGBvGZTC+yeHkb2nqOzWf
3MdU6Kb5XYRp19PdJ/lMOPJvQwonLFLvU3He9ATViCP8lg9c4h/wUXic0z0ibCQ+eelBIEpW5w+R
vjaBv+m98x3sfJHHCwlWlZt9jbT9MJvHmAcA0YoCSHIE1i0wOxzuNy+8JCXWlbYDdl/iCTTPnY9O
ql1NjUotIahW8jBGkfoZERffe9WLKHI8tLpjJZrzYIjYIjzDIjUO81MRse5kg+OumFLq2SteCvzv
bbbD7mWBl6Vu6ngmW8HjvIgPpMTvPGeX5H4S2Xo4NN0I5vNl36wlId0rEcc3YZYaJVWJOGxHrb5/
d0H5Og1DB3ndiT/PZdVfa3LsFD3Z06yJvPD0n2PIfFnSe7Wfee8fUuGuDZLQvcpiutVWEG0ZoJEU
YZggr3h6/4wkHZgRx+Tadu5TOSCP51oZMpGyPfbSlw87Gg9KX0DHGjieCfTj+nFWiftlg/x51o0I
Kcs81jS/jhMliFiDa6Zpo7ZNEx0/H5sSvFSrB6n/Klsu1Ed9oE3rcwmmgaxqIJGwxvIQuw6u4T6i
hukgQ4+TjyBj5DVSbz3PP0UTblbZeup63n/hbepQWtar5ew8hjYDyBBEpQp3/FiDeIhOXuFtsTEg
Cff/eUck/uN0jYs66OVuvCjLFkoxxv4L8AuTqs6vIyKSGtMVgu9QfttDDqu+s06PIyjM8ea8bA55
e5WoI7OrmeaKczssHBOnTksVKRIwxGFm64V+OOu7QlbrvsVxutSzLrCuGFbeli8otHE9P2kFAIec
hq2ISKfFCosZUsksI2GnECmtey64Nl5eyConilETU9qZ/11pNFqxxBp7eU083Puqi/aeT/zfO2Qj
VsyeGWCo6/fglFWzevIvGlXW5i+wYnSGbd62/GrV5yqX1z2FrMI1iEEx2tqMuk5zmx/xl+NoGyTf
6xfyQkGXMgikj0EKDUK/snqNFyfdC0rLg4dAOxX/F4ep+AuAY5dqzFmwkiTml8bQ0dijmG/xt0Jd
BQayPDHflnhwunlhCHwqsqJ4/R912Rsmar9KRS2zG2Yyv/iL6S2HPk2zpHu1lu8Lux7VCjBc9iEV
ZGOoOy91jwV3VDcUt7vKk6lvIErRtao8Xbsl33JfiTh0x7ojjsFb5GxGfIz57PFX0w22EUECTaqX
JiObcWIzwJGA3gJ9DO9HmXFqT1ADmDy9C/CSJjEI7bczT83vKkiLD5KGUCeHdSeJ5rhcnc88op4P
Kd3dN+rR7CrAqqc8xQPbFCwNV2LoGOvVnrsizD/UvKAtv5USemgzzXbVa6llW61NH0N8K1BdhKFZ
muPfFABhxBklvYcElhViDOM/mofJoGZjAIYhtk5/S98Nx9HBuGtZGSvhx0utT8pFaUPo+r8lBEaC
QbTEa8wpUQp6FdnwPGCHaRdSMaG0UMXYkNM2DtP0hKNvsRJsraAxn/XkWRuN8MqkkLhMh5f+l90S
d7rLRn1H40Va0dlmvctRnljD7DWEjmZ0ofLgInDLa+lt20pCZjyP75SCv78gktql88e2OfDE7Tjy
UfDtfX45TZk6Ym6XwFCEX2m+vNIkmUHSTn2leRW1Ew1kBnmluJM82exyjMovtE/eAjAfbGqATziQ
ueCVuST3kkgETKtRPCSNfr9YrjgzPrOOWX0MGT/qEbp33cKNUSNxxAnqq2+Ndd9+uruc3yfcnSmW
k/7/9aJz2GAs9zwYhzD3QAqNiHLqIN8RqJVPfDOpQZYUCxF3uSdW54+JR2kGsujelZaVhvI+p6cE
NKaGuIKZrqSIma2ATfXt6gRyp1TXpBJfe5K8rAsJ55TNnglTkX1xH2hfICbRN1RAXmzOlnXVhfBn
YNhoGxfGx/xYg5fXprZJspyZ3QJmhe0arL3wyx+rpKdceviGp8iI1kRYh+GHbkD2ao3QffXrrkzA
037dGKKiVBL7DYhbSIYTeaeY0SRGMSB70RK7j2uxpeSpTHQJWRDR4gQh4TETgjfpZSqkHY5MG77h
z6fwsFEIcAgKKRYKD6x3JQLiyRWMhGVt5VkyWuhwEKxsHJcECBYvYRn1hFtabUs4aj6JhtL6UzaI
1S4Gu0p6ARexcKuI844yXmxTluOLzJgTf6LCLWF9Af0rtJ+eoeDIfxfHe5r66XVphJJWYdQzKBhc
jh/IIgUgccKrnoDNjhrv3K9fO69J6QCn2Z4ZqlbyQLdnJhJAynmni73LepdZaVd7zrBQtOH+uNNG
dZ29cgO4n3E1AJZLJ5SPw2+6f0rDM7GNp0pNv7TzrVZLS+L82o0VUJ3tu/i6YIgPzS84lhm3vlxG
SxjPVmUM1/6YFT/b9Vp0ux4It325IopoknISTNsB0/q4xgfKwlSVIwhavVeGrsi23ZEgHeqn1sjw
Ml0tVfEqJ4MjBTZRa/pT04KmhahkvcsWH/j8wxSilpsIddAZmVBOvyaLLE6qjQ1gX39v4nQLFzv2
SIsWL0yDXDF7kPhgE0IUM2K7zgaGoHs0tRIhNb9Mxf0WplAEzivTDJohdk+mxxNkbtuBDrJmSA8I
yoiodZSuB9hbFFbM4xxB3I2jbKRKkjKm4OKN7wivT1lCSPwJ/qIj0tPccaWkeVoau/3b70ydVzFR
04hinVD5+nKGFrFlDL39Ti5+TqlXzEjHqfhCc2BaHen4FX+mVLbI58HvVrOgOxU+GnN0Bsiiztp0
QJ5cwLpPxP0/x2wKQnMBcHKJsEv2J25bT3AwGXg4NkhjVmCBtV6GwiCATdEt2AIqrUT88YDI2iw0
qyusb1xjANvbkJ85FIfdfdwNFHhLbLPCcbv0OVcJCohpgMDUM/3BKnMFYOjp/CwhF0P2kGittV1j
t9+cigJ9jTvFSVGN8f6ZvX299wVRkJU12Os2JSKbohWHj1aOOuPa/hRJliXDaMw7hyIC+Vbn5mAN
lWPIm5S3Awky+ckXtyqkDEuA6ix0bNDw6+HGfQt42rN2/DSVWKuOGkzGyixcZqcsCtp8o3koz0H3
I4rFEDXsMEq3U7N61SL4YL6NrmopZVdWYzt00MKRMw+vyiKWijP+Q6tMmohnVapX/TD0/kz1hWw6
4ShWrZLVUAaCbmCTL0Lb6ndJDw465bt7bzL+JwOXGMNN05vkMzhEJD5w3H/udwkmBUDO+GVW/qzf
sqQV8QNQAxrxZOlzLR274BXXrJhsxEGDNnN3G8YWGkce/drXueA8WfWf4vG+mm9T4fb5fxnFy71W
sSYTlF6cafvTMa3FkLNziNyK5etV/TARjgPzxt5+w8D8ZKlqLHM3qWOEZ5NRvm6ZTUANFBraFPEg
fafw2AbBaORSxpJQGJ1IV186LVI8qte0EO9LJJ90h2P6FK6EtEs4kAO7mD3Tq7SQSDTlQIfQK/4k
L1yEWFrj/C+bFCM6DkFA17rjlw6K9XGAJyuvgcR3JFsqrcYSWLj6aQyr0gPh96YUYEM55TEtsbal
jZh9qIqdPKwY1CgIQg39bic/qJkEMnNw0TYrOvvrz69Z6MgTnTVvZ8l2MWqdL4rBzRk/wOTocnLW
fZT5UWIcIuk6KPN3VHl5/63ImackbqPcrM58gEZgmWE7uQJ53ltMfX4RYvt7HZxyP2w6VNnxFmFf
y9AK/GPwY2TMohk1BFH5GQ9scyCQ1dfeVKSfJncXsZyLwIKcD67ndEFaehC0Rt0xJ8GcHU0blZdb
dQJDy6Ce8uepGn/JzSG8klBSgBujpTHgcksk1EXPCLf9xYbFPoKWuZ1B+NHntpMxgahPSjhmRs6k
rusX3Bdjy3H2fsdjT5W+F4Cf6Q9jAEQXKxw5FBEkij/fKBd1LcmUZDu4ESAgL5tegtAwgjzYz1Iz
EHKiWQG71lgVyXoYJBIsPstOF05Y4/thvPG9B7VCHRhNZVHzahAJfu9K2mHyEqJRfMTLjYZc9b1A
GSdl6n/TOrXv2jaE0yMrqzYgxCog9fe6iNy3ShHIz/1Ei1mcOVQConIDB3qaNovVP9rO5evSChBv
mdmQWj5FAepmRHrb8iWz9PcrtqishlaI/XPj5zkbC/hthiFJCfifYX2y2zqlRwzK+meC00QHPGj1
9oXLCHaayZIZNM/TvV/o0/Q6f0ST3lAqFi+tcT1s3ggaWH/gl8ZdLPYNDnAxNkhc99n7WKcWkeK2
x1fy4hVhY/9s/Ut14pyDtiNKq/n1A33/X+wwAHXpBmwE5aUWBmjK2tTvzHbs58fUbuMUnW8dfVGl
SZ/GpBTgjPdcWEl7Xb6QcBORXNj0XSfOJLygNmk5nf8lFhJWCBcmx6EN95ERgO+nsLkYViNy0+dF
TIIYGt/vK7bjoD9Uryj1+skt6+Hr7eFl31GQwy5BtvPxJpxLiIjKpwoe+Hsf/B6samYPg3hqUnZ7
ySW+HoHV+ekUftTzvt9bSnslGUgOLVpf6ivr6Aj1RVHtg8iZxAY86jxBOlStE3ZUiRVozxkkLIsE
lLGx5I8iKLpaHd3lVo9tHgQ+Y/y9HVDLxUqbWUsCL/oQQveXvELOoA20Mdn1GsZInecF9KLkIkHR
3BXysNpxpSk9rxGOUD+3W/hdRsVfXZekW4pSF7CnWSQNyW/l9goi/uh0aq0dYWGHEWL4SN3Pc5LL
I+Bpn0o2L/MbNJfoI0hi+8qya33mf2xwyUUxoDU3NQq7hwMyZEe+84cYrnKhylyXxOWV2VfqHQIF
7hX4oDRD+ahcXB5AMr+iOi34XJThwvI9DN1/J95AJldHAqJ/8ffemrs7wxoNQm1+EucEwyOPoDA5
FYn8cyoqRIC5iF+8Ff8Ok30NuzriuKItS6kF6zjQg1LhCFQWbM8XHIynjguD1z62LDBl8eMDmwk2
VQO026TffV9Eb1inFq2paTYRHcI4alEK85/53PgO162ml0kJ79dtkwC2zGR0y1V6nLpnGEqxWCM7
GlE22NJEgMz+2yLKXahGer6QdqXEwwsnGm8IfjHdQNfrTXQgtZYnpOGUX+BMfG5FKrs/zXN8sfb3
swJNALXVFmRvXD67nJVmOS6qNwlvoGuWejt7pgWUSRIT6flNG6zbQvUB0vWhnlZAVAa6pagbCMp0
6aAf/H40eRQ20KQzqcFuMu7TBt3/Sl1ERn14yzQBOAIjYvmv/kbc0iB+jTe93W5JD41tpuq/ND9n
VgMmEaNhF+Qjjyaalo/Odr7oC+XDWmGn2LUjhOkQ/9qewCaitJyG66dtivCXNClrE6DsNNA5CNKA
ZxcFKc7JEnNlE/qw+btVdCphmTqESJqsh+zWigQ0gYkUFd+9vy8q0/n1TvYUkpnpv7+XF6kycv53
YAeEwrLpxNNfbbywhxVUFPKHw6cm++1RiPOwMwdSOT0hN95aWybF3q1+N2xQVaEQ3J2BWg5GLiNQ
uN3CJM6qc6CZuGd+T9HbcZUiGJVKj9mOtPdTOML9+pHoO1nZgqFKDIqIIv65Cs3GiyocpHEYjnrN
flg60eUuFxBaV1wpg5Ern+TtuxNMuGibAzJ0vdRjZe0RD4lNQKVq2Z8E9s0bZ7wdthaRgKMm5YUX
RHJZEjYo5Js7vUYpXEjkiupXI/2nGajUypk2lcA0UfuEnGs0KmBgEuX6mZLgCHzEbC+f+U4jtyOe
fxUbxzKSoxAl+UX+eDI/LwPIsfqvqTMXlucBjCTHPCsxfn+fyDfoJbJH8WdKFZR8FuY5VMahpTCs
0g8nhISDMNTDkCKhXdMKXP2fBJ/TO6MI+qHdER2hBJlAPLSaTeo8XzW6WjsxQsXVqRcn6rjeqPb9
TyfVoh3KhZtAPT+ch99H35/D98N/BIiuananuyahfwAsLpUi0Ipt/mda+RQFuZQ/n/dvcRfbQxf7
janduASQEEuSDuFbvNyrEt4UxI02MEQ8kEut/7EvGx4GetXp+3gQ+p6pBs+hhmcyv5s1tpgINupG
ZaLPBVb96OIUtCcOzLCk53aRrZXNomuc2+/0EouxafX/YX1CRRWsG+USTQSSCb8f4q9Lb+8G1rt6
khZxqvAieGZdaukMlNYMFwOmQ9jiruLyW00S5HMpERgwBMbM3lO1bFmgCLyuf9f23n1UYtg1bQv1
InUPOYiLgTFMddpszWLGViUovhI2gfV7xJkKHbvRuEwXZwqY4NI8HjwSHZfFo5UUPrpMIBNBVFgk
xbWjOxdQv9QK3qgdE2sbP51Dn7Y1NAPDbrRDrc3vQDHIJSEH0hu0vFHLUL6gZh/b5C76zY6Byr3D
ecKS/jjJhz0CV850dPWJGHZPdq+rwrDLRqrspVScpG3z/Xm3gth7R9zpj6PY2xQxnh2WaD8QZLTA
3JC7TF4ZB475A9V/QYVz09nmo84i3XzNiNvRmIqB2L01MIsac4fVjzQLa4ns10gfaoCwJYi8VOEf
Osszf/55kQV3LcuhqlFkoITbaIlwj1k6LIsHFX2VmPr11KMn2buirADIGCAbDuTFaJv+x1mnPtau
1RgH5XCx3m9jtJiicQeoF8a0DgEC9wFuTxm4yXegTnG9aQ80prmcAjL11YazzWYLfTv9ikTQpCjY
2y6sbZq+sdgZw4hbKZGDBw/RJ67Qp0cCcf5Cm3+cGl6zrKIeIQPk3XUb053OdFZhRLMqaiCknQJY
SSd1BN7s2tGx3k+Vxxso+epL70Aqs0yGr9l1FT4V06nLvBR4YWa7MJJsaN38EBfZizAMZgwPpiEi
wqlG9m4Tx0y3HXv8WLDggIIOR/Iu0gocGw7oVNXvErh2SGfhFbiPUqbOkrEOoiTjJjK2l4e9lD+B
termptcSvel2bsVnXd9xfCSpJlDcWpLF0x9iFFSHov+0cJUXbpAzZn2mBiCmk9v+oypnbiR6Zrft
AmZopevktjZymLwtM8Mru+xTuaJdzNkA43xN5V7dRC5TF4zxH4PSkeXpIcCCdjXYbr3iDKWZsBBf
hUYh2k7uLq+FY3LkvAXSLlfZs/GDDMyKhzbbE/juekyNXzWkFcckkD26keGDXZV0GrvIM1twE9OQ
YFbYsBFN3lGcIDwGl7xKG2SzY+7yELjKc0NlJ13T4H/Gk9eGaZJDkaDXR6STRJLVb7yT63hyU6tY
Xf8x45IiJjpW4Cbt9zawmJqZ6kFr6MPvjgFea4PAqpIzT0tqxK46xaUVXUBJ+tPl7o5dgJs1m1Cz
NRKFhQr6rccW1F0VRRtzNIASubg3XlI6r2c1VNnZUj6vSBxsMt4ormyCgulN5olobT9tReMTSA72
L8b7BcJRTwdpyKuSnKiwxJtfywughHiJphikjmOEgVgwxgdK7Qw+hHT+ZQDjXzac/oVmiK0V2pAA
tv7RRR/nZsKTN2opj58wJO2ixru4TMckIGgmDFI350tdgkQTF1axh2j0j2tPMP13GWjZWgAEGM8N
xjgtslPUxSyr2t/6NPiAdPWrKt1K04Kjx1UGksjC74vRdyv3CF4SGVmbcLnZZlDQAttdWuvdbQjG
Q4/YTPSxGR0OJhtg9yGdLyplT47k/jrpH+KdiW8DcboMcOb9cJ5/kVBOphoG5hIOn6rstwf4Ybld
Fw7AOBDcKuoJB5dlWYdmhkKzQL3eYoQ9F1YJXdte8UnxusICKZ4hOIaLxYe/jDCMVzKcB+8W5O2C
bMTxqE7Lvq2KZ4OdOU3jEccxiFkaa8gmXSSididW8EPcQgZ/rJmhPOOsyyapAz8LV2Ltm+hty6+m
JrwS+gOx6pEDEYfxx06Sl4tgdw6dgLmEt2e9cFUlEL8bsHwi3YsleEgnPLk9SEkU6rSwL5NmBneN
2vl9jFz8a1DMQKQkgwe7tyoddg6gCoar/e7RTsRiDXSwtNpxE5o9WJUiwyIRg0koz4vywqLjNJqk
GPsR7bJj6DJox23/QIrHGxIf3pK7osj4tVLTbgIEOUDuLrInbkAdnYAtpPwAMzLxP75R020bzosm
QTpcdz5hKGKsDQSlr1SRH96ywZs+7m1BCHdFH+t/QfbYpX5WDIHAxUQ1KgwyvrEwsRdPyU5N8xF/
qqkZXnPnNfb8nIuRMbf77ReyB08WR9aMAFe0hmMb/5DYG6MnikY9aZk7DKOiJzrSfA4s4Om1DBAB
wf7Msr37DD9BrNlrF0l/kdQiAJg3wnKZnTVv2C7RPNtuSEz0h1lBliB7oC7Arc4R6WaobmCDBhar
JpDABod4qbJ3oYCEbIchmhBmi6WnyQdONrr0/0kxU7JBQWwGjtZ58g+VKalRBkuJ7/hy8M4Ik7rW
MM2/DKLYfb191lxWyLRgaKyZJow3zLBnXAUV5C0/ilqe/RNJm9HnvGtFZIWAm+GE3OBLKAfsoAGW
TJCdt8m884lOGT3gvXpnTdmqdQCYEvlhTXCDCwvC8LdN9P8liFH9kIqnID/YRnga8jHi+kgfK4MH
RGRGw6A9CtIwQvEdfrbCrAfdvXzEs/LlfCVU6Go5j9WWPbTEB7Gx1Rqnz7eX7TcDCOmSc65SZqdz
2iU9WVQ1ZOomaKJYNCHE6avgmZ8GHLxqN85iRZxvwMiFz8muoYLMt95ZUIHCumX5MtKd4evLyxMr
UaOQaTbZLmChubDBFuoCqRcNSSVizYDyh41wuzrr1WleXu4ekWoqPR8M3+12Tbe2vypvv7S5tLcf
j3+sm3+L/sH3y+hmS9j0YTlL+3RMJgm0oacXd84a76AEgksUeN0aHEn3IzBRuiUccJ6Q2R6K+FQP
FMoU+Vmet/mc8dpksNPgIw0HO43MjG6ufsDCWhFwPbv81w9FLvEjbDdkcphTJGu/awTJhhPXojvN
VxoXdPVSzYnlbsuo9As4G1OVfZhHpoQbOUaKZShT+wJrwU6rE3f9cgM568dTOBpfw1o8aFuVcwNP
K6U+STjobxEwpYg1bvIC4+4zh3JDYwih4FjbRytE0GmXbcTBO/mVWa4AlfeQfj2tAdcXUZAlDHqc
vh2Zu0YVy7dfqSNIQhaWLn7roc3xhmcn2hZG3mcCu0u6sKxd+uYGEvmBQJk+BDscNOEotTIXFAjJ
xTXeWp9EJ4sKApJZFqr+ghnselbKmxNGqDpZngj1m0ZrzrHI2EyrPGuIuAQpw7FUCza7pyV5QslJ
V7Gqzgvt+k6F4ou3ryAqNTueF3NJXewnrnVLzl2tGR2zfBdoVTEbrOWFuMj1L8B5ykeGTrNYif3E
jjpVNH9NRoj1tKm5dI52frtZDrf8vTViFydethhX2d5L9R02Oq2FH/z2zYW1dcyfeHC7ezz1tgIb
AgTlLKYL3zpaZam5KuA6teJMXzXT4XcINtu76zfgSxHDZ2bzKMVjQ8xz8eGmL5w2jNTihIZCHDZZ
3jHzuCjXncwTVsZqkxkJJlV4s0626tcmQGVVy8glqjydFEHxi+tiFqQkk5ytSvpfzTa/Irutu+gA
WDdcSdTnG1aql3vkpqEXzzmuKelLcw35j00whgsJSJYN4F21qqi4uimT148ye9GmvPam6bB56l34
S/e1q2/DysDE/QsFBeI275TAF+6Ke7iI2HqoCZ0s3BA9a24PBVOz+NH+8YEaaRJpYlQMQMP0VW/W
1eKqwhL7j09XMuSMJetXfTrxLT7B/IJihVOVW/Q8AqpxA4taRkqD3CWGyDqx/jVFTOgxNTbIt4pL
YOtYMUWUDi85P+LDpbUTwAxL5qiioMGeu55H0cZpWYk+1MGuz5wYrYx1Qtf0XlfZtxrxYwQed8ZB
A7K/L+z6flDUigAF3qJrOHZvUKMz1CKDVdQ2/ACfwVD6wWYDV2EAgTSPgRYxnq3sfL4yblI4cnGe
Nzkq+GFvv/zyh8cS7KhJ4c+YdBmh/SrD97qksuw9KWTDR6xZlCCcSwgcDZ/CbwWRk9yNj7rVzHAp
Rf+xHH1xlfqi4z477/4VGbMeHr7CFQZguFeD2IuHdiV04sIvMBXN2aZLaz6Ud2DXy0+yxH42uM79
3O3OWoCd0M+8mDerSk57/R+muK51IvKIqJlmRd1WxUGQK/Tf99iYigBjtA5BBFf5w0qWyk24PaCE
kXvps8t2HwJpf6101vd4H8oMHt8QxYaesybC4bDKbjHZnW96lU2FCpXP0QlGnaweFgw92aQbmvoh
DVfjs3rNREB/0wlRpnpZgQaCcKC8PxBHLTlRCkFyOYea4c7Kftwb+as83NbzqiP1pePVZQivS5S8
R/z4txWa0gLWyo+Cjxh9yYRWqOKJTUdsgphQ7Ly0hZ3Pd2PbD0+uGcU0SvBIOTeDInFGvjuW++Vz
qvTLjeQ8+cwzr4ZMoXgMaLZE30nqFjzDICJ7iH3MsN1A57kia4t8F8LVTYciOtf5VfTCKBCcctES
AZp15GElknFjGqtcwINlYvOYuUO3N3uZPrnTkiXGMeSSwRe3BDPXjbHl7mBJtwNBFmtRJVbKeDV9
yEdyMrlWLe2mnq/RP0WjdHCHauOR8pgRXj267kjKnsX0UMg26VLst41eHZw0uMDscOMrxOu5kdpb
t0rRkhlMOa2P5z8KqbcfYm3MzIuJJb0Q1LY92NhefLEjVd/E/5NyhR9MzDIJeVrPuq6fPfd9CpjW
k07Wa4T4WUhLC7UiqegM9rU3KET5iM4b6FSrXeMF8IwiDZkw+86sU/XWFHK8oEHOUJn4w+dIklQ+
uBIrWSW/z7dVDkewU4KU1OVhLANa6OjPnGwV3WhXEck6ob2SUpQvjmDO/rcTCdmPt2XP0pyuSfEu
Qybr93dbWZviSQMHWO7ul/yugbJDi/+44oLVtjEi6/NkiU36+uxWB+yirzdipT0c1SOR6Txpg6pR
snpSpIgIJlp6HSpnur6PFtP+iEv4SZXWiLXRA4ChLNIBdpJRMakCV3m+OG8748oI2ataausjjNd7
skqrcrEr8U++c3Bs9P8gzcb0pUdJVParcoQUicFiELlexyxd1hgc1qzhPuKPqnnlszBmjaJbE06a
hwSx71xzhK/k5jelWon753arqgR3Rw4He4GTArtta0RBtR5pijntpF/v3DQ0a0hjmVFvt6/AJVC7
XKvs1EMzrosLMlDk0Sakmho+44j6njJFrAPjkQcG73TutNtPGE07kw4751aAFo+64s/eO8Sn0sTb
IImHP+JnW8H7iZSBSEfr43GbeN7kcIadRnEg72JLYi3qbRxbnPRFTzzC3cdFyOuAej9mGxTDvam7
7HT5tCBt+0fvV5+yoLChOJAgM5tmGrLjeWHwijRdVYs8jK1AD2jUJxkrhbIXU20emdn9vqMFC1RI
ZAQMUJ5EHKTgfEhW6FNh6XuPqxA3o1xvSyK4Ch1nWS7JAb892VOqDbQs4CyVyIbccnLga9r0ho3d
Xu9bnLZWZCNpP0Hr0LpKA058l379pPZKA3xQNOE4GY89eLeraj8Iq25kx9d/GSqS3ytf5CkuUXAG
JEt0G3ApRiYRJhdzEsh2XUDa2qiZGj8Xb/eDITfkG7sIZ3XNBn1PfqnUH2k9T/+8aLgXbVm1xypq
sk4aiAlH+1t/6p25B1pg1eqk8wkhMXT1yOblTT0UhYL2k73Np026MsgERPnuJ881wmzN67P+Ecjx
mVpai6aL9jpWxZEEYqZ+YdIjn09dB2JpUOIxLNMv8odCIHQOMwnGM2tJF6SiTj73Dp/sBo42Iok+
Gbeo5w1yUvUcYcI9BcvIN8pVvhDmM2BP51ur9iaqvMtLPFzBvY3+i4tF2eAXni/VV+TyRlca9F22
gZLWf4XHtdpm1ws8UMWFihxjq6eA9QDtnqPOVkAvPwigsnlTwfTDHdxaClNToK2Gs6Cz9ju5/nUJ
psRVAJh/MrHXw0NbOpCiEUZQQbd9Yt8vMirlsi0SdimUBg3AoEJxaPUR3rBsbJroOnG/auXYDqCi
lO017VluOprtcCLWTUgEu4yxLxPkgygnLmJwVwCm1rfOmtMmdIDm2eVwjG8NQFx0qIPqzMNyNcNH
+N3IJVWoPwIGR/SvNswjw0xznAlEhXXHhE3vFIreq22cGh5K5Bx2Xpod3bfiLyckaOLOhC3/xeIQ
MrEzGUxGHKgA1PplhI4vV4I/KS7E95xhhwgG7JD1X0WicWUAsCRSsmWPlfWnv+JHd0FeGY+RTo/7
Xp2MXR0z1dOGFD5BalNI/A9sheWA7I/OgsCwPjKfpS0p/pb4HtargrYAmFFTDh5M/kxZ/Bn4lavu
kBBo2hee2J5rUXArr+bkT1m98f3GUE2lO3DxJAofTWLg/0AzAB9trH9cuDuAHsaRMVjtY2LE+htZ
6drZ8CryymGSzVBjyAhEYfU+v4bs3Ktd/wGyCg0z6CzsLhdZK4iXOe6zXyUJtLJ8FV+u8QAcvNui
nGKl5VvVsPDhybu89abHT0r60RIpYtFx4GxnYNt4XYIC8o4+Ewdh3/ICfRHIAknUEmitc01h3BPt
NqiggJjWfUekf0b8j5JVx9f0NCaVmvUf+PyfrE/SiH3PHamg6i/UHCCwVphFopYbGr3wijfbROwg
xBR8ak2T6Y6AcCvMPQNcUMEmJcRPIjt2MAv3Or9v7ERW4SfwlwgtACSKt69Kh+EU+3uo82M75ZWt
CE4ffZyLLONkHS+NBIoDTIfrWSGxRBuEguO05GhNX5vCHLskVtFMRZdJew3nE1jUo6UnSD6rlNYL
Jft1618PglwiFoVWzfkFu9S50jHftYSUs1VJAWdLKa4IB77M57KKJ9fRPzhMdv96vHEE1ybf9qsd
C3FRvi3it+mSwv2d2QgyzwU7vUaLNgYc5Oylz99mplErnfXN9DzOl2AEzhsqmHmu2cwNQXhIRB/h
Wk47Sxtx39NNzeWxPMklcddyUobApDtzJ7qO1xrt6xN8e1I5pFCR9Z+PBhQDOEmkFSk32B7RMzK3
NiSeb0w+yJcTEY52cijvGBT5j9uDj7HmHCUVu6jDr8nmLdNjhNjjEUqBUVxOnt+AluXnQjex5zRt
dA2sTlFIVuufV1U53pDGquuSWzQ12AClJigN/g3sFFLFHJEzvBztHXJgdKYyEFTkb20G01t8GURu
OunK9XcU0zymmIyOg8o180kfWMX3kyZGWDYGj3Ri+lRhBCULsOnmbsTZ3LtcIKysXuW9uZtezr6a
ASOAIGJJHyDl1MH5IkYO9qdYGMbPF2sCknTEGzeqXgIM+COzVPc5R9UjzpohSI4L/HX//VM1sUBY
gRGu0vuWXMZTzIjBT0VHfGSrSfSBUBUDrygsD4filp2Uqe7H/G4f3LMyzcnh2b+l127mCPojFTSz
6JGH9IL0wbF5ikLkKR5SQayRv6tQCPWN7J+EhbUTmPlH99Yb+/4nbxhpcAVcBzzHY/0idEi/5GwR
voia1GG8n/xeyQ+Shi59/uQh9JKGhOxEKcomuzpefoxmv0FmXMHBgZKxLQd/RMFSRAhI/m3l2G3l
rOgl1ZmlOdxJcwufp9ZQK1Z4NQRWKXOqqB2r8FsgL+CHf2htMISiAVZMHdEVss0GaD89cXkMuHJ6
V2tpv/snPnBoC4kSKhpC8iLiKJ+SMOA7/wEdiFmRphfM7IeurMVhP40I26ZVkrxHhl7gx0j5Dxt+
UUZ/a1QLjN/HPWN529CLYBkzSS34kZDQ5sthz82t5sgr3hS/4awcSnaAgJwyzqiC6S93XNpCiq/3
dcwaSn3tnwfbXkT/cfmiKVBqvbLIQ1z8DKBiTrBI4mWcgRllW7KrKmXSog6mjQdQOpsB9bwcMhHc
tJClgAeO1sSR0k8scVDrTaTHXoaf+pf8znH6UHB9QDdpjKdZOAVmuFVv/QaafAdZLexRAJdNoTS2
LaiPiNZIcF1eReFABs2gEU8lv8AlNOWz3E5Ks0AnMoCnHzhjua+UVetM4QXZPqJ7D88nckxDWMjm
WCkpXScZL4t/4qI6uyWf+krMDQKsGleIjvBWbJAfI+zWch1bnLsuN2KxpjJxLcoWunLJElHq2cgu
2tNX0ewutXgT6p9kXrzLxRv9G7bcy2sjKs21DfzFpVKS8AeNAE+EsLOZnzb7Vnbcz/o9gkPr04pY
IqudbaIt+z+Qe6nSvUNITWtIahmx/08Mo2xljXcV2bp/EJF/rUagrBqNBcd0tTyz9IqNuhFoIiOP
2yGJNj8CF5omIkkZL0F/KM8h1oTo9AH7z3AA3efc9Ra+hzA4wS6y5QIWO/of7z+gqsGSlF8MkE6Y
ljp5+9r3KrUcIEs1TkltQnPYDgfd4p86kYNINB9H7sjP5utk75V9RVU1QVkZXuyu/D8boNcLbbN5
izeuBL9u5XxOck0u8KFyxgHHSaBAYuVXQDOz54XKS8EYgdfonX1On6bZlWyhR369gyLnrG+ZlAkN
6IuT3PL+owirWM7s3hsPrkeuzYc8LmthrSV0RN9pIINGS9yzAy2nsu/lyB6GuUkhXpH2vyYYQ9e5
/1dBdtgXrEnBSqUJyM/6jtnNw48rpphVvTMXfreuN4takn+gJ0lbvMQKQUKF+/spbv1Ete7ZZNaK
0aWM8AWAyhK1psI4JnRsSzy+cpBkxh0/Dh9SwlHvwOTfJH7OfqpJih2cJCWwi1md/fkFbjyPARYp
b0TYnzMGmIgHRBwJPis8LLv7AoAj2Hz6yYmEozoSD7tw0EQ8FmUW+XBOJrXyIENkGOWL3lZCjnuw
aMbbF8F9hKnxXVHsoXJcSnihgEp+xrMdKxhzMU77m4tHeuJAlgXVeWwl0Cmt/e5lTdNOtgrFI/JK
cM78pzbILd4DMkcalEEjZMoszzhPuJj/ZHKIn18v1+DUtj67TsDzZyjMxv6/AhUjXLxG8zSioC0a
6EsCMjPP2/VwAa6NVmZIX4Kr+WpiUgH6ycZG6u89NPy1Gb6ZBlGgn2pObFAacFdiqqzkQ7COqMkE
MDI2lUxeRiTxUOq0je5nIqUaL2hbh643ppBQCVsUNjxmyxUT/58YEmbrRtWd5fJjP5+SMJlFTPwh
oxive31NBkdZl8k7M6Ij2MOVYC+nV2zF8pdJmOHniFCq9uBY1RYFb3YDoUVuTiRpZ8cuCkNh7soN
LryKItIyrHQxKxoBEjm4B+MhNA//mdKGn8myQCfEsMkF0fQ6d7bShwmAtRlbk9gzTCk39MnERXtn
F1DWAFGLbQCR9lMUQjq/GoMPk+WDMjkB7LqtAlV30lvQv4o94FhtKbVqgFy+YnarvXVFFOVQuiKb
qmbzjrKswY0pNxNQPmtGcgWcYZetVtege6HK2pf1pbkZr4fcB3ge9MopLHnIYTx01XlkLlOgW5+Z
3GgiWgXgAlKi9BxmkVqn+6dWYbuOjFjt6NxNG5jm7wQn3dMeM12LvTVPm+vPlSUqppjxtxBNwoQ1
3rQwHMvsNOw9zp4ZL/CWAbXLVjK22Ama5/vC49kh7LNeLv8QiCDV4rMeVm41b12zCeL7TRPNBzqv
M9O0BlSAGKslCEiDkyl416RDVoowjlDOj0GGnpcq6SHVLeFqpg+ucgTHmVnaPUALgmliRTIaBohX
bECMPfBauwUMxW4qUvHugXTuQdA+ipizJ12Aaged5BoAZs2rCKFUYMgN2hYBHnaoGp4nqie4dv4W
oyzCFAaKLAZ1hYpdGssMNlh4/8/cUpaaam+7FU+a+dAeE5LfLaVslkBTxilkQs8xoXvmrCw16i7X
PhjKZIJDzvKU88yJN+2TL4BXD0Q1pGcUA7heDAsdkfWNUxi6Urz8vJhy4jEcFp101ndP23mM2w9P
eExfcINqJ0tYVKiZSo2E36S56mtahEdTlFRTxhcgrIGIorzXEfX8psDZkM14sShlwpM2Vir05Qzs
LXfBnRiSvcSOUo0vJJj6N/43b+e76Gbf3G6/+PRtdAwnOZsk4Nsxmeg6kBBDkgyXgZWiX17mYKnX
VYcgpkBrQf/Dbqhzj1JmQLjuM50anI9MHVZZ9g8StjSc6ArwKI0WIvGpgSm+zLz+n3PTLBgfUJlR
hE7usq10iVRwMTQszRGjOn8Vwz7PyKDfHv0tEcSTjhzM6DRNB12o7mR5oo+CXyU8tuAF/hXDGZFc
TZB/7jM4EwL3PKGBBRanmDJn435PRkaiyAkuan9Wu+5A5dY0Ie2Zdcx/08NT92UFmlfcYQ8sB6g1
nNgbLqlOfbVWN9G5IM0+fjD8m7OjxGVJcozIVxTMUXt4VcMavUI5f22oVRE00GmMwOvQV/xo+M17
k3F8wvciunDvwjHjcwW96YmrRBl5TOcnPg4HaSDeUPi2vcyWnm8fpIZBLDHhw4UI9rfe7WULnaOB
YDwLg4YuRtH4q9rUsIv3j5ptNcAFFrATe2Y+UGzJ0pCvpwa8EoUxLMNh+sgsluWjqPfKAwpUaUHo
FKGFERNFxwthQja48vQTsyj0ObMKFNZVZ1/2bZHJ0pkSqGO8egcODXlmPAeev0mh30h4luuPbXVL
z/WlJGvbHX8x9BZGVgwN0D8DezN58tSUV1EswF1+oEG81wOJrXv9HLq8FwmJb/UMtRdESb6vIrWY
DlI1nX8yy1r2SKFwJ31SCilD0SBjsl6Rl1uJhhpyWFavS8rVcVZyy2Z7kOzMbfUfe2pky4QO3Zg6
k3J7tF3LY9mvDEYpnGVGHfc6+dzTJgB04Jp+UcB4fS4Yz0fMW7QZx8Ox22tl2+yDmWfx4y2KObmm
Lar7FqMZ73Y/mlnZMHg7fEY9FGsEce+ZyPOj84hW0CMlpu8UjpJb1PkXDdq/vEUL7n+15gc4pIOK
F+bQFwWWYpgy0hHtQlSZkPJIm0PGleG5GyK32BwTMmAqgnLDyGhFGN2rvJNE3yKz0CLJgAX/HYon
hkbw2jj4Ui/Qs60zGAfBCxB5LxfGM3/ehFwqM92wC/D+V+vnYvzaQfBtFBPUBJBEXhONGcaUna2g
cgyVogeq2+x53glBQuej6+K3yd6wuiYzw3snuHs3K9mP1zRrLNZ5Fd3xNQ8n3RkuUyWSonj9BRry
siaOdxzyY16VWbSqVA5OSu1VJhggMENLuYyGiOdmAA1Oy4fFko2IdpaHz/WzxllZgPaTiZvrKzWE
kk2Sy3q8whdYO18vUNlR5lMJNv/O/5Ga27pxw9994th0RlG9eGdDtolHiWFAJuvUq1jBB/3yHjGl
KGJIzngsUBbxunT2xqdMdVJ2U5DGbmdyCwVL0LxFPm3YhCLRi0xFZ7VZX+kuQYEShxy2q5yGu6KQ
zrZMWPOGerw7ibyyHqHRoAx7BjuVGorh/WhXyF3aPI5Nl77139co/to7jM6LQAiRnrhnfk8u3weZ
bGfnjYXMC3q2yqqhuZFeh9A3QLh6A2kbCWm0YpSiUOcup8G5iR6wmQ9oGthCi1dxXD6T6VMFyTGC
f7deboy5hOb1HRNLcWnNL4eoA4JBQUR/1WgHX+bgC1ylreK5lYW0kOZLO7Yvqx5+KuRAyGxwt5Pm
RrAl4tlN9gYVd6dA6D2bVZqFn9uS6clUjPu7atAT/bf3CS58PexY7q3Mp6nnR9C6Y9Bf4qOLX6K7
R8JXgzDnmMzCZCpnS2FEhATFLQAlhKe+gKzkYiKaJPpqG9/VDnKSVNBgyIp5xiTXWRXFcE3Jellw
V+QXSxUiqmoh6PQf6xcJYd3dATbQkZ3FMrg0zJ3Hrwj0KBQJRd5xe3euQJnjW8/GGZT4uD8IE5Yw
aTKiNC5+JQiIK6FkUcK5btcm1A8O19LKBIVRn9vXIcFWp5E1KU0cseq2HmaZIFQglp7hBxPXLPa3
TlaLOuSct9U8cp2T95YIYjZyKqnbQ+jRe/9j1CB5cg/DezKlPIBZpuPaZkr/3tEsBYUKNYEdpkdx
b/6kxVnTge9y3b5eRHx07r70I4Qw0RHmymrciwkj1+az9QTdurhtCVxmAlCrjAz2Z6Zst/36UFaV
mN4XwA4COpNqmwFVnAvmiihuaLkoBshdTSPVOujhByK/1NY717qrLlWIGBIeWpUU8Iv+q87oxaHw
FYdh160GDlEmimB1E2fBg7kS3eES9C8G5oSsfNxZoc5/nruPhKibdFHe62sOnLbKuhvlzNMeAPk/
UJ+qrnRgXuXNYQYq6+CSMif4wXV6lLy3Fly3gfBjvMnb555YeHwHHqYai7SuuXRLzQm6JvrcAVIH
A7q8S0XjzvPC9cPGJskxukF12Q9AwvldVfLg1tQrI0ukOKRXkJSDjgFi2LJzKuGIBS9JIdA5XSm3
4q6Vn+WU8NEsays34iS/AstTzCiIe1Lds3kcnVrN6up6tvJoDQeLueppjWuE/7fM+cCQvWXtZbxW
MMDe4DkncaKr0ttv7X4Z1KD0cvrDy7S1Bf5oZ8Cn+tYfGtnkqyuwEEgkzFLdIx2ZG+2AcvYId/qJ
fUsqKCD/qxheP96snK5OJfZIUPotarDn5fXb914zeIud8JUj+G5FIrdC86E73sTJx3RZ10k0/Tka
E6265Pp+fh6PpEx1iuyhHyiltfGf+CGPM0Q8T88tD4XWhWRWis8nL/GhWvW9TeRLbzRcSZvF8Bgc
aNdjsoUy6hVCe0EZW5wVfhw3J2dcAzNphOUU5cMqb2IErHx73yCy9xzCTFMoN+8dl4X0xYl39t8E
QqIUNwJzecis7ysmSKEgV+zmtzgCEzGoUxm7ZkjiigHV38Hy/goV9LCx4ZOvHd22aePJGzLH8vaG
tUXaXTNyg6BjRFmgXHLQ0uqSPhENZ5nqcUyEGOlcqe73Q0wqeO0jGxAvV4GtWvADl+93Tqbwnge6
0G6rbU1JxKwzBX9Uuq6x2XXhRWB3KifcZLOTQOA3vKErNcvqvIHpMrchI2ayQ79jEzwdio/HN4N9
2yJM3/pmqLnboWRL9Q6HBlsvy9eMwTg6qdw7JgLlMVqxMGIMEivhbxw/rpRdqarHxmYwR3694hbe
R2moXRRQWYpsOurtL6+TAGRRl5j3R3KTsLWVlciErJXXl3heTY3CPVG/vACVU6ZShTqZp1n/ap0D
8wh+8YRvfso63HVMoZT3yldwecuXZu4rN8kYsh4uI5l9If+6UR8IctXmL+GF+66YAfQANIbxihh1
QVCv5c5wYhFZCmwHhoMuu6joYRs0LW8rE6hfN92HujITzjTgjzy4A0VUG8gluT8Qcp7p+Bkj+fI9
PhwQab2uKVORFNz8auUnUNoBuM+RQmR06RlrSreW1xprCZo4JvWr4PScmjtwxLjSitElNHZcQ3bZ
STg+1Ms1nYgFga3EA2ctnTnvxws19FGaqB/hjlWXcXsgSt0uMu9Etjzz8X9aRmloFFkyFuVd0OEt
2WABIVglZ94A01Ha5nJC882cNPJl7sGcpDtWjb+bEUIZMddi1bSvXuFR4KIxKEDVE3/HtVd+p/JQ
s4BXzDnaFuYrzYEvCc2DLjuLWzMnNg7Ils6+lwc8jkHHwEyKqARiWV3D/bMA7zi8E0wFe4KWTClS
I/fgd03udQwTQ4YxEhSDW5Ahv9tGX5juDMyjZLHM4Sk7BoCrBD63oDherDUk84mqmvXpOUBT1ZaI
4Ldxt2kb50NBbA3+Igp13mlk+krHD68cG5duSZUQ6hADRdQK+OWH9PZrBtw7w0SZy3WOrg3TeB6h
3eK4MXlZSlMoQBqlMEUqDwRo/SEl3QxVEbBvzcDqHpEt1+emS/NDeO2KuWzty9nW9kt3B0Unc4bs
DqBZGagi/dB+qllIhTXF+RC+JntuS/Qm8LuPEyvgxMOx7NrBtJBfUXAQfNAzT674qPH3bVROCMyg
lmwmPacu57+tLOoCEeRzYRt09l9dRU2dCLptKSo6L+WVY3ka9kdkz39sboOo97fkXhlV3gitwgHN
CReUjgq0S6Se9XjPobUC+vmcpNsPf7+kjjccHk81hUbM0XurzIadbXOGpPGwhWBhXZXr862Hc1Mj
SOztEEeyCLNyT1xsqlSpMPDxRBkU0jzxFNDpjRvqvAMyidYb3K55rARNT99V2lzEpkCJabKtnz3m
xNp6Ku6mg53ZSOGG9tIRi5IXhzRsnmGD1VHuPmPgJ4fCjd7G98F2Rs3NgkTBt1hlzzMq1gq26Sel
GBWZsEyvEAGV6IutnSkplBim+7Ru5eCmKP0isxAJb5MtvET2Zdj+4Vm2uUf8jqRYHIVTeo5A3gjT
UVHj6m3p5dva7bYfFQoioyZxCfgxOVWHvRQhjFBKTYe0HZZ/fJImKQOx6U/BG+xBqSrN+qLAYDKI
vgBTJO7YHBvxLZWVIkZA2ipc2OeUtpNy4LwvE0i+7PpsJUxRwsYblDYJuwsrMmrvDrkLAOo+0EWz
SU9MKODD1YRGnIpqhCh4UICwGhPU4xAk6zKIcNs0kYjL4Yb2TqZBC6cu3orTPVnifXFCuvxTJ1+B
/tRhhIgqEUrVfkHb0lQkPkVDZ1L3zz+t98UQ2YcGoReEGljklY7Ity4KFVpN7pRpHZInv9lnOruF
cOq4xiV0ntzV8TQ2eb+L8ms2w+m6TJaK8tvLJa/y4tVZftVn+wjlOYIxyn4a+1+enFR8671EBht2
B8B6VGcHnvMLCoA0hzTOdqu3/ls9AcQYXXMSsuTrph/9KjTiEge3R/hibiqcjYiXT5vfInmATdCp
RD+TW2qhJ22AF4TiQrZT5cGDuyY/obo2hCArXFVg6GIAqH7FDYjBx/Z+uSZGawRed5hRMpU2MElQ
WOREpwuNKIj3anRYvlNXDxeaHDVFrY+tYMgXaCnq1OlGNzmV52dCL9PdK+vZi6sD5+AWeVTPQ84l
SUqp2+xfMV3BpRRzP7VPrQSuoPr6nF8PKPH8upwnscbg5A3a/+Rcl14XvZSXD9HrkAL4mtsEZr34
g/WEiLni92wQLCP43ZC9rg/2v/54h76y4U3rWXw0gekZnsBdoLVVrzD64ezWJsR2ATtpN5NZHzjr
OBuUbazu91xlomQwnbko31ejZhPENKFEDCuuALNb+s9R5x8KyHqLFrkaE2MDvzziVAINfG7JhqWF
ep5R8IQYSqoe9JKwOR1eOWf1pSpJRXhx/IaTjwGIDRHh7y3GCHXde+Kl2hppjCv7vbmfFlqmPOl2
csGkMI3aaIe4Ccw2mrEeQNzsgHKHdenGQwLflN7fgOqYMO+eHbPyMi20MEYqs1TZAY9wWODu0EJc
ednRUbHVGuyouqSPyDQG85u226SgTkoBNzrGFyMTQVHq8zs3Jqbh7QFonclcLHyOobnaM1X9I0Pk
MUdCMtdk7P25ESuIiQ1boKMScTOfpoDMEF9ctKqW6Q6cmKvzdoJ9pdhTgskY3IPFir8enSDv+pA7
x/A6iKsdX9k4+NQB85TYfdgYAXLriQxpzhgzk0elbLYVU7HO+B4/rSU+Y0M4Q1gRftCKV6Cfdggb
tSdzUah7hAbWeYYFiMkozYpelNMj84vIUOzWYsWa2NNadIdFfehN5xSmqL+4a+Os1g2jV0Y/eDvO
HI0uu7cw/EKXegUm3M4UlgQ0q6yFJppGwB5S6tiO6K3R5WG28TpXwd5U3cDthD0AwKaHDjVhomrx
2+zIT3nEJwxIAjSZmKBvY0/VWJNZl/c+Re0KRA7zbfxbox9JTZmFpd31abVrL18ll2q7WpZIXMsk
v9ettb0kGh1PTSOQ/NKMytFibNIgBYy8dp40Ea712RaP9n31vzkrj4uNDOqOUHTItCFrdBMt/PcA
li1hJJhEtaDYPgKrdmihEpGWOFQheAaYbrRJmQfeB7s/MCRU3+te6VAurrHYuunXxVGgzW8UE50w
ZX7BpcCCzi2ggJLsckGwKM6KwesCiREmyuM3kGAArxwjayAtvCgJ+WoEmVPHosoGoT2OVbGtJJZx
UsBcXEQ0eQdp93WA7mEg4detk9jF1ajELwPOIsKKvkHsYbvt3idTQRqKsPCL54BfYY/IA47EPyE3
tpZpXAaTsPE25kZdAhbsjPjMSQIzHsfdXsK5nt678vpHjIpgEcvsgTcfn74T7wzJbsZMxa1oIQA+
bLs4WD/4f+hoI79m2gTJVvWTVxjrUsrPSnpvPPshZjnwiFvb/sN8tz5c8yTUm1+zCrsh2SPxl61i
X5dfgWNpyDmMAj9/oSGuctZUj9Dz9J+zG/cGnnaHwfcaopRflwIyTR6NgsV5a9w5ddlsipNeQ0R3
6yBqxKnzkaRWwPydoV1iRAXv7tZHGGk3T7JQ1hqIlM69of9ZvblxHzFnAV+qm0oBFC+DGEV1BICP
0u1lFYtuA70DAQwu3CfT+eSMDnEv07fRMDq8MUgQCNuf26jps24k7Cfye9wr2MiAeO9k/0LWJpau
ZSBDhRQWvnoXT6WUVWjyBi4OmLZIvkE+Skqf0EWZyqnNOGDzdsatcCYd9iQ5vXSZIkh5/4DxRrT5
Sogt/5ds9pG+qFelpedSEVuMoSlwmL6MD5nQKGw4lWmBqiifR5Edd4phvKbiPGSHC5dCns5GhL62
6IFuayPSduGYsquaTflyZL3nxJaONv1c4hX1gOq8oe3vYvZJsaxTKhYdsldw1Gpqq8A6JBMSkGVR
GvOC5vLIAFehdglIZ1tsyBkP2exMbP/n+HeGsMjmrZ4Ymju4xBBYIgjqtwt8UbEjyyBzzLEEoaZt
q0xxykSjuo9hGKXfwdeRBpI5tTw+ariTqkW+LKFGQVD8Cq2ZgCdVbr7+mhPk72JzjPYDcYLBV+L2
KISvLm2mWK4M07cu1Z7KzFYSwMfRoORReb2/LIGLi0ww0ahbe+RqKu8ERPQe8EJHHQM2NZBtss2u
EJsN3HHLxUCRJNEIeXxPje5fG+yb9A7oUzvNiZA5MVPyYKnfz7/8TVFeoB4H1uzEv6M2GqqJiZFr
QQcxS7NxQ+R/UmkQofW47onfbc8ag4ijLBSJjJAwVWCnIX17jWIu7PJmsqTSSjYK7WQAqrcthCvH
ORXoHsGgGg3Zgr53fA8+VJjPurQo9vZrNHk7SGzzBUbzP8+iwkM1H7GP6gSIw4cZIXuKSqh/9AxZ
LLH+D82voc70hHq9iIfjI0DNnRt2q67fIEXtgRJMol1DdEDqn0IVpj2W5mwKvs4YJLVZwldoosN4
touZY9vZ/YVKMnvzC//O7k3tpbrEh9KlhxkVserQaA3m/3qlSnJ7oYJ7NXYg9ztWTO1ghBiwALZP
wwRi3wqHKP5jzq4hzArvbs/P9bQlij9k5z7dsLUKET5iPlD/RtQ6UULBbc5v+UESy4cFhlLs129b
ioj7UODcEGEEY1Guj5+y6wvkWPhQk29BKZHWIgYuresdY/IHztWlPBWU65yqtF4tCSnO2DslI6Jd
zjwJCF44q6ur2aqj8CwtZOCMvYLT5PT1vbBE/4xCczqNuBDAiJ9+wBgxRSjLfqkEzl3IColro/Pu
4n3LJFXxB/ji7b6Bco3QNOjjwgu3pSnxjvEbgKFl/JeYmt791vWL/IN6kAUZF+yRGmZed9TQUBdG
sPyGMUcnlw7JMyC1NLIwT2JhDfD0JDa4g6dq3a64noJ9mbLDQn269u+YQy9csUg3NlUhU7ynh9it
dQ7cWtCLvy5u6Ck7RlQqDA5bZE/Ob/DCeqAe068Wtasvg2ST2/BNCFBNh1qguOOnp4hAgu073kCa
2dGOLIyWf6+DVyrY/fJMcj2R7ojLOpSyJA6kuuVIc8JHfnCTNtyrwlRCUqGM0oQpN36B8fBHpRsO
iGgFRtvRxytnv/DNmNGm/zgsxW2yBm6sj4tLbF3pvsAdqKY2VPBqbqOSeQZ3S5af/o5OW0fbaA5o
D5q/Wewnhn21BTbWDU4zsTpAdYAOb4QydsFyROcS1xVChy3BRWHMIbh75X4xwClUYL/Jigk1B57y
PScPfIV56x+3+FTp73/ZJgoq8HxLJqlqiDwdO/aTjCLNB/BPzFBozkvjhHGYURdBMmEDqlbI//9p
IM5+5nhn5UrfKCLU7POfh6L0JoLk2yXTQ1thk171LFUWoPK7j12ZdFy6O+CPH2zixJPIFBhYVL/Y
+0n6ksPWtDs4HN59IBG7G7R3kSi3RwlMB6PbgfZkyv/eYxWuvjIhj0JQeh62EFlJtONIG9tQeHCP
mXkS+nVcreepAHosnLwaBi3l7e3D8M90vfJq49E9FFfHhFDRFgXAUQtf49zIQhOUQ87wO5DIiDNw
CH5m/75UZ/ne+pkTJQHhgSP4AfDoXBHyUDEHmW8KJ2KMjmjrRL031u9HuLRhuJuCnJWDYHB9h6MI
xdkBplnz2sqwIIIE+7MqYZjZsB6Fuk0JBpPKlsD6pZ84MtvK7p9PQ/AynBY1JHhJfLbeIv0J1U74
77TYoycs8bx9xi5UofRqMwKfwdhKFEvz6XG7qKR3vzncvjdf/DUOjcw5lr3jfvC7zbFIqLvbnche
x1aI3dtbrq/KiHLFmIK76ykMxzZ/nWadI1vaXZ4tc3I1jtARfLvOo1jQCSpZz7O+RhEw+/gTGKXe
skm46d3C7SWtXt2VEui/vFqCbJLm8uJOAzQ+PLZLkkM+OAGex+QVbpZ9ny2HJj2Z/6lHS04OiDPI
kSSoosXXJwd4PT+IYx0TUvqUeDs7KrQHh0WmP88av7KsrCga5Uqcf2MZJKJQq9hGDHGZ+gqmXXn/
fBn5Vnbr9Uljx0gN1XrfibqwfMVrDi825nvfHhyOwd2jHlw9LW21W24JLeOQAIdSHbnWeiDWyLv7
U5bcDJxi9WWNU+74VSZlSp9PLiCKMQuaSbmUT15DZFhuJGkYtJO4AnOFq6AD93FzdYVuSpxy12u9
xBokieRi1Dky30lI3Tin7/zWdD2ChIoDhCosVpVj5sW1AuDQE55fsN7wcI3bsO6kn1WEb5TwnGMb
l3nxiTLIFMLn8R2UrLnSJMgji5dJLga8tciR1s9TBbizpXri8MsRZs6qIGd7stR8GirJ7x2PVjug
b6dtoGoon9UstbuulRuKRw6SxsRYFZa75TzZhJWzFpc+qzAiAMEkVDAvbX8yqfQwDuunTOhJE5gE
iMPTomOqoD1tRzQQWGzM3QT5uBvdT5lRWcxLv/y4ALpl7bjdOen+06d4YHu9NXdMXWV8C0ZICa66
wUgNOCqkjnTVL3g7w50Y6+ruA+3Fjj6dqDwL6KhAf0k410ApU+GHR4iZBspiPfA524IIoF8c8rYg
BYuHPNv6XbqCEIpZfm2w8R0RfT7lXTnYzespYi5m61+z50/V1SgCetSVr/l7N7XiuAY4wn7mpXXE
dN7RbJkrlpz0gw4p72V1eLDUQLabKgxH4JI9qsJzjIHH+aS4aWHALVeJO4KBMbc98tbEaLgH75uS
hQKc2MwQbUYCanaMBxDec35EFZCI+qr5qctOk9qOULOYaQZDhQSVkdbswwumqs2ZmJaU/1HYETHS
ecp+U4pRBZDhbFASK+gaHrXfkO35+b/m8aQ5LMoCha28aDZCr4jpYwD9yZ7AuovNFrllnIy0sv0A
0XHdsUs+gq7i4Y+Pv0N0HGcjwQBucSMMkkSL6DRasS9w6Tj9+ndJ7Z7ofxDUdB0fRwh8Prv1/Vlb
H6UR8yWIachdi60w1vrAZ6orrUvCB1g7wAAl+tApQzzh2+CVGX4hfbW8azUPIKPvd9/INXEvlPmp
mxVvsT8+yCwYCuem7Zuhl3K9MsxlMHuyC6Jt43BSA4mcwCf1iXJe8gkt3FJaCptwACeDGQ+qUEqN
3SGzYMQZWVw/MwL7AMFLvMIcQE/BtTIkXjT7kPdDTFWQPh4acFG7UgJufaNENCvMARR3QvAeFxNf
YrlZD06cXlsKOvI89j0LNWhWRuEkOBy5pl5rTPhIZx188jM8ZCQxEW0pKDxhjIm6pcnV2aqthKbK
tCspyvoPRV/vJV2xa1BCXM6qZSOm61Gr2KcM4HQndtoTzuYevHbw6Q2IPQ0pZm9+O+MGjyt8JNBN
c0Omkwrp/gDzlU45EmswOhjYLmIziC1yy8jRe4mG3FGgWtAs2v2jSNtJ+GjWKKpE2p3Qcv3Qerob
85+HJc96XnpVZ4uBdEGtOc2+0DwXxarnNyAMEepqelykTQseBgJfzZVZwInPKJ9ZwK543lNP8Jgn
KvFo3T/nO8e9YN+xLdYKPHkiZFiRnk3/YazQXVKAAMfYCfWm3CKwkc2QcPUzuCCP1fRJal+t17gk
cWMSXZ9HEywOFacnLOQ6ehneYpH8NkEPWS5uv21n8QgTWtk1+hiuJQojq0I0gMSNIU8H9W53BCz1
XAMcnIahNGJjTZyTqSwJrFfjuYAP/4thBC7ZJdng5mAKrtIXnVDhPw9gO5i9O+vnw5R0OwZwUTI9
hUKLxJP0pIaa4UjdG5RRqSNpV9ZOt3t8uSrNinwzgWbMA6nH19OcOlZBM7FK7G13BK1BL71Sxpqg
8Ljio180v5p80PXv9XVyT1zBOTqGQDcBH8NCyxksusZcpQOVRJo7FZftQMyk8HLyGHfvvJCnqA7X
B708yUWlIsVm+HnRPEd/uZ3AmJk25i+wGf23fawQLfqg4wNU2zlOdlm+Wyx4ykKS/GZtV5dmUETD
kssfThqfPZVrctoUGOLzVlZdnbT/wIqAgYB8/iDotgX7YXtnpjlp22G6xDOtpPYU6ft10C2T03f7
1YdO3yb680MoQsyxkHlsmDkeKjWP9H7XNlMFMBokjIOkfix/vqJJ0mtxBXr6lRmNH09qBFDont+w
mJmIG2mKaXpf6HySwtgkqQvBAA1zxwpamsx0IWWALJx1/iBPTs98Es5Hj9aBwXX8+ZkjCksKS+Po
yXRHlgWp6GZEOw+dqGLXIu2J73uCQ2swLX4ojLZMFjAB/Rdd5+/Wbs+pl5e66wG+t2yrqKbjg6RQ
MfUHIJq1DngNvGSAfrVA7NHZWjn8U9kV0leaxMuR59EmYzpr8OCcuOqu6DVqPGqQxvnGjJFHYeO0
vx6QX0f533MeFbf0g6hcyEOlrqY4r2kFv5hXquAd6H7HRWbsNckSxSHy38VE0EAqoBsf4ql0AQYn
OQepQIyvWr2KAK3RGXQQCevo9LqV2xEsOXLbkWnVzf+f46srMuUimuj2omYNWbVQ4bidmQhqQBjI
AYGLpEnapY/jSLInKf3lJWPZd+9797W8qYaXXrc+s8epUfQzMLRwxsiA7X9fb6jD9Aen6uQ/4qL0
4V3/XI9CpP8tc2wA2K/g8vgbo8pZpMe16eRt9+yVl1h3auuYeDqVo9nS7VdxXvkhcNlficDPpFSh
4XtC9PCTT+96yUKqBEPG41eGT+WDEUoBixsLVPU0QILCZnuQUXSsefc77iNvptxYck5EG6tXm1NB
eZ+F0Vppynh743pPO3z918C7MYalyH6oIHUX+/X8KljnP9ZphMWbfKbw/5G16U8M1PIaASyxTxRp
Aaz0wWUNdzJpXPVAS7fjac0Fs+cilclhcMgL8jWtV6FMNTOtGLqhoUKu4iiudPAC1tmTeVLwZ6ZG
d8kblTmpKzFCXAn/rEdHuVJvZiqX9qu1vRrxaIIdhWAwu/RF9UtVY+IhlqdIdKhosWF1OkZ+GYlx
KBaAH6kBRZHX0Us4KnOM6cAaPjCB2PaqGEfKof4GKiZgc/TGAozGEkebi38Gt+hOcFaGhd+SYD8X
n9yismX2GRj473RM3VnirUMt6wYgmadzlUcDSGgEF9F9p2QC8qAeUct7rDWHFkjBXr1waHuxj+/Z
AVprUCxWYaErG7e+FukhkzE7aa/+K6K06c3r3097SY1m75AVRqVYXskvcZAVAuPA/k7AD2Krk5d+
bJQtZPiUt6iW829MMqS99/8QIHFpazEg+/UJO9QS/aCC27amT0sJgmShtV1LUxkKeMuOaVF5A9nZ
dAp2U6XTZLNPjs8rTrAr3AUd729NQF9dUakK8mzpd0jln8NSv4cdGXWsMuA9vgDgGL5l95t6PvEk
NHFvucNGQ59XIix7rqp8pCXVzJjySbl3mf4+/C8Z9ymq5KOXL6DIZN7TgflQUK/Pv257pLHH0U8K
QXYrFVEMP4VPdIZII+bYF+BbCBI5ENiUSVeLGdoCCeMay5AZQcbmw/Mh6sUOvnbP6PJJEPsADPL8
BVNOFSDVsVKYQazjpMqgBEjdF3vKFoc5RvyvGju2vGyARmP2AAp/cDunzKqJHpLd0fdPtYrPl3n5
37suELi+CSGMJUhlxKo8kSJvN6ICXd1FamIAZhSKmMHDnn3rBtPmUNbHW7lGzRQDn87EBMUsO/8U
UeGfPyb6Zxb6v8ZWvKGbTUmk0XxFx0unX/1GBelmoBKlkqgcJTYsHai/ayw40nelsZf8hw69vgyw
JJG7CdTJ4UtV1nf3ReDkpIilCKAQ4oM5CFUM13Hg1pc4bbtqc/VtyUO+kxYm0TuFbLThtPfuVwCM
6A5zQLgXFXI9SKWXKsu4Ii8K/5/skKsFfIW1j/jUTofjNPqrMZww2bj6dj36x/V0IspsGtleaW2W
XMkefisB1YqQ+onIGCg1va3H5TkRoJr3X8jaTqELjnhZ+YBHM4fY0XRz4JJVD6ec7/ZpdofoYPze
0TdNWJVG/GAe5PlJORZqjBZi7e9A7NntOXgNyZ3eOyt8D2UU4aImiZ+hLv2fpXf5SmmXZt8eMgiF
4AETxfSDDkCnfXt/hmEJJMB2QTv40p5ybeCkVI6WwaexeL63jSWWnZ+9ezeDh5YuXBK+goox74VP
+AP6r13PJb+fSLDj/5nrwD/4Bc8UDOLuceWr1F7BvZZcBps7wXuOl8jrz/gbYKZTRO/9Bj/UlHXc
8Z5wDt7L6+81wOlP4RZh+JviWTgeUZnlDoBKN2ZkGFhD4w28htEbG2zoRTh/Hz31YH22jQc6bVFv
IzX7vc8sQpFRlHqwEBq24wVhc3iWKa2JZUg0Gh3q/msVvFnChi4f14/uXqe4gR/KTD4M1JNSDGwO
m69Qaw4/zrHPcN3JGPLzRkMHYtyg37WkVr0pKzPFRkeeob1jAwDs2eGM5FTx0Ix4heG88dGJE4sQ
HbiMbyLeqiVrzvNjtX8upP0ytw0z48Amiqw9zjNOuPkWr5I6fFwD/DFMINzsi3+4LcqZRtRascWL
PLFX41evqFGSUEvugB/kqS4dDlH8KE8qvvW7KSRLbsalikXX0AabcrpwdG1I+wYJw0BfrNY8SwwY
Vfn/XFNWUdiWyAnL/RdZRCZc1HlBsnfW3ma26kvU0SIYp/rugbNk1sQhJgPIDgL0jIyrOjgSweiY
YuIeHcKR4U3qfCAQlIRwgSAZUb3tCjAbkDJz3z4aus+WXckXr9P4/R2Sti4paQ034aWp0Tl8hQ+G
jshw3h1TKhgxxeTr+jil7JcF+yHbK5PcKSV1xqxcTmX+HURtPjzs0DKzgJf1D5bVzT2v2TY8OHvZ
OHzM/aX5Oob3dCE+gVUOCTtdLUJ3SNt675xJkIBtT94gXSCvo/ivuZcr6xcurGrpu7z070uv3syx
wFpcW9hVosMTU8iq4NvsrnmoIcU5t0M3A3hZ2jL0fBu0fCSEf85Jk0FImuj+Apg6C8w8m8DZGRYM
q31dMJkt8o3LCkFTiRVf+xEaz71PvO7NWzCBIXNlY6n8p0eDO7hJtTei99Hoaue+PCUIGnZV/hM8
JEBkNqoqif/ps+ra0zWnUSbqy5AauwMo1vZStGB/5Xy6RpH5GJr/DJVBEB8kyYi8ZCgSI/T5g11v
wdq5SFuZzvTN6xi1H6Ohu/eBx+4zvhBmVN3o1j8T+SO+1HFPT4bsRzwPKgHD+wWRCvm/t4xrdjFM
7xmqUHfAcwjBIGf3vUiqeoFQJvWRqR9MPM/gP3QWHg2krvE5oAleUxWvYKa0Gc+J9N8ZK+4egNAj
eG3SRloV/cpGi7MV+QUsX5Kt1JW/eEpDPEGLbZGAWr+1A5JP8oIPjQP12YbFhx1a2q1i0Cij3joP
lye/tSimG8NWE1hUNwit1PW1BcE44t7AZTA43n/U85YwcBBN7TSScm6a3znlUzhBjSvrBoYc0UIA
z2tYCVmEibjJWAxAvHGBZppQW5zwVyTxCAIHwLmncwwSJSlBRCNfZTuLFZSxyBUHyguQSIAxT4vg
OtW/zfuxdvYZxvnSYLy6GYYN8Pxnd3i138eRitWCFdrx+6rj9efvdxa+g25ZcrBx8EQoxzsfvx4M
zGQqLyqiN0QDJoVBLPiOLsCsdGkKFnQik3Uys0RBsEzEcDNxI4t9cn0lAgQrXkBWMycNEatWwO55
Vg3Ulzt8URqW0Nk4zjy/R/scGdOlER1XAOW4Evzza9MM2DTSF6AOXJus1vXOp4Gu3NSwuAwN5V/B
mUjO3RY56F7Hew6uConyfJR1ihF5A6uFuKm0xepNgOeUCyQZwgo/SdnQBsebC4JeVkmdYYIdJviz
gpx5d5YjP3rNhQnQ+byITuvWz9ejbg/wkDVrhg4hLnFMgzfRs7fVn8RPlotP7+ape7GFn4XlAqkg
f8HbYmEUzo2VzAVgbGCGI71kcxvJhv+Jtgm7vD8S5pV2umPqWEF7Bb7jWx35xeUCbj7pECkBQV15
taer18+jyhC5ERGcrhVaG6Vvuu2MLACcwLsaQibyQCWu+JYtrTxkWHposQhMwhm8p0y4WMX/M/Xc
z8tdMqpe/AYy48eF6AZsoTnMWO98zmH6+6YsgMZmP4UeWZVeMMkylnuh2tgzmF8I8LxcZf+wdmpV
Isat5vxB/c/Gjq/uALtFbQa3yZfhDg3juCUzPX/qkWVMOuA6fECyiJpxSIJJ7VXLDvqUCKlzlM9s
0eSHIvzq0OfTpO5gLSXIRPjM+pomM5IvQ4Xlk3FEJN8MHOTBOhB01i48T94GWozGe5Lu8RFK+t9w
v97C03HuDmJrkJRE8c71sq7Jm0tQPR0ldyDktLlI/JJTHdbPcFvuawj1B5agb4Y8aqR3QB6+KT+I
PFB6B8P4fmFeqggob9gpxQRqmymPC3XGZXjOWl1rMuYNcbVZii6CmBRdogjPcXzG/o9Xjf/qO6M7
oTjEFaG5WKzC7VpXD6f3o4BjZmLNESgecQ60qevWQZlfqcxDMmPA+s0R2iFXSqjGUvQnfqJSpnaY
c4QxrH2akOP/v2VjhE1UVW1aONSAVhWOUFBx1kuK/yeCEw246qqyZv/pw7K+eh3nTfJhqaIy20R5
GHyzfA2M46sGQI4x9mCNPtPZk8HdJLusafqEZTso5NYAzlIlDhXcZ67wFjuzq/7+E5M5b/SjkoVf
MhnivEEoa3xerPMSNWgXHThNC9V6wkSBKcqu9GyFDtjgZ+trSm/7UjfaFw+KlSmkaKA4FHHtqMvQ
88MKodb2WLRNnMeVMPJJZ0qRrj+GfKCED0inEuF+AhznqrWcWSY6ntdpzUlwCsPWpG6gKMy0uEo8
X3THw2eH2GF+5SXhLdQVzXRzlWI4+t3H5NNr5yON6weNGt8ZxBTh1zw+TFHQZ6fe7gAZYbDISJd6
XPs800niZQDQaMgOSPZuEksP2CzGQoA1jF8NaA2M4V0HI1autDzSmr2ZNfvsIpYociap8gNP7h3k
QNCGVjH+8A2ETnT8GbaPbcWkm4FMcLk6fHbC/BCtmpLaFQhNRl0NB1vRN8dLLmlfqV3sE7xuWyKo
1K/WVw68mFSIqKT5gapyGGFa9BN1xg3xcH5zLLLdVdp4aZSOE8DBweODbx9SNhbd9T2i+VME70E5
ckhuyKJYVf7LRnMY232aBkzv8Cc7+hOQItengcef1LZOQs2PGZetwcZO4MAHXXaxT0rxXKMfZz9s
a5yIIxNMWk+U4tso9A4UZmlRm4Gz1b5cIlVOjow/LCHJOVoBmAhM3oQ7fWpezNGqbVr5oGCs1nNv
lZd1q1t60O5krRZkIPkqatawjAa60lCBTG01m3gc0+4BQf/o8KgD7id0gIWLBBNaNC/wFnYDK8EU
QSbm2GAbKfZJjLsUtFqgoVjJhoeqCoFSWh7pEdLttnqKwED539sviJYp4CLCU+anpSi8S4PN5dAk
EAsgGZX0PeG3Fbc7n5Cgoqv5XhKvVX5rHNRYfyxrDRpk1WaNw7sobZmceBJ9HfhiDnvJGPmt0UIP
Pwqe8EsK7GyFUslmSPOlQbKgvRZgXm38Uc5iz10ZBCWh7Tge4TpS15Rn8v+0/FrOmSmakrk8ftwO
QrYVsQKpMpXYiCeOmsgP0BsDyyYT9OU4JOJ5IdTpFe4Uot8EH5bfaiaJuNOwBMbIheU/VgNnwCTF
FJP4xhgfwdPNCjg8VGVk8ADOnQzL153Y8moQ/ug5WntAFu2cE8QKSrcOXa0AU4ncWRTRcDHTgyer
t+qqoUsGKRd2FXT5FbomaEUzC1cVamUFilgqBvdoA+AOuUoCmXcG0lakRMaeJzYz61MnTdq3YVzM
ha/45DWYyORs8Otnat8Qnv84+XHGah6wzY+gEVHQwG+4YR+8Pw0uuAKhNC1yahKMAhsQuaEc1aGH
SANd5KZ3NUhzTjWW9ERVbaPD+eSid68EH4B2skbRmSldsoO5ZW/c6b7dc5VBljHfhK3n/qOPIt5G
RkyFtWfcFUB1Qujsa09iKhkaUCVIzVwxMgCJxnGRMWFvG8Ju7643ctOEPA8O5VOU10zUg7Ka55r1
fKaMlhK2MN7/0Zpf0TWJ8O7onhVipeYGnP5AcUPC7NbGd6mTY2IQ3oSOf7oahI6rAQPEdgnZr/uB
3+S/s0WYAMiUWasfPL+SUeL96qWdLmfwkuxydWxTlQkqltymWNv4r65Kzz1nJ+FZSQsGavKDJIGM
6K9/FhJH/bAOjpcrije0mVTSuUJctdBBGXwE7V20TcDUzp0h7ZBiY07+ZSjbhtwYvWmb5nO/9LGS
cGC6P6KN+RTOc++P/fXKsgYgfPSMo+Ya3uh1ZJN7aJcJ/z+hc5w8uW2KKEtZyG6KVBN0R/SyXyML
bbKMcKYHqPcAzIo3VbPoMP7tGu/QFHnNgpN2Zd0D+zZSkwozW0Uxe7YWsoCA+ugIvW8K8OY9jVgU
J6CvZbmhbgnUQ9pM7CAq8Pw2c7pIdWJva0eOGzhyxMhSj3evzWwk79f0PObaAuhD0Y7YssdMIrkz
2ixlZddpJOd4F0oyw42zEjWOhAvwaK5/g+b93r97dWOXBchf9UFFEQj1QvuWbpUwK4FI9WkjJTRV
4m9nFWuMdhRhMXXA2bzv/yp5aauy9wCDurec/wZPx3xItbS0HvuTLZvPbSZX1GFm+9ifZm34oZeM
xUkNhaP+/XrOm72LIDb7An9wL9XfzLVVgAnjyL+Qjon+32gfKf3P3x5P7T27I8bRMHeiVBdq94Mm
+t7tDqq/For1ubGHPHSvItcldddzXtUdag67R9mskikMieGfFVnXUpcpxWimzooVR977K8mkQuRk
dnl+IYAYJVlH1x00VoFeLCeGtXKgeYDDK2oLjWBWhUfhFRmv5dEamw5QTra9RD1Zp23c4Cj7HCqN
zRhk2Zi3+Q/IYFH2nnBVDb6gw2nWjfxbAO91D6Rn2fxKrGAXuxtrSEOYjAi9WwEx6VKUqa5gTs38
t7shRH286aSXwkv9rcOVeoS0bIAxoAkrS4jaRe408o16Jptnw8Vd4YZyytB4DD2ZDDOCIuFRtzEQ
IfeUOKopMvekDEe0zgZAxWgILf8nAsZ7QvdxGgdb+YSouXEVS6QXEyg9rlE3zYpfZ9cwkL+Lv0q5
SKEZkQvBmtffgzv57NNrU7Uem9aIt0Oipk9wN4yl2S3IUm6aM1Z85zuk92fTcQqbPGIIxtYJy/EZ
RiFYolkmr4dipzA+TMYCqrbyXNFNzPDCHK6W9O1eAC7XZArrsybPbPjJdjsLWxatj/xpMDVUMSu7
hOr7dhln8yFpCHEJT1CQdq6Zh+5I1vyuHm9Ulg8hjlR2WlhVjE1c4AlU92aCkKVCBxUMc/5C/+Cc
H9mNjoM+TZeNNriCxcFqqksxzKRDZJV6KE8l3gUerVMCYhRaAEV9OyVgr2Zf1/wXalMBPEZQt71K
FftbXBGCB5Td26xT+0d0cYbF0ic0QX9W4WZ7EdAxE2uJBJErZLoulzICGtIZfQ2eB305WzEZpmH/
RkkiUG2y8bRrpTpYzZ1RJSlZwqEZOta3Wn43bS7X09qqizyi16KrkU7ZjHqnLoOzBQY2MyZIKY7U
kdB2hyJ6Jvk8aNt91LfYrfRudbzMLFtNasIqkgObTTvBj2JFEEixt8PDdOWGzGW0T8xxrRiXTQcR
poHWHqwiT4TE0wgmEkjPfmtk+pPQ8Nh2T5Q76eJHXCPmMCVRu5gqwNomfJgY3RH2w5VgKM+4CxGN
LrKfXcn3O8Ldyhe0lVBmBTPYA3wHHsJof61lCfKf+f2s4hoI5i5aig38MIx9SxHyDdqhX1KBCh1R
ln79NocdCKlUVpLe2PN9ySCWelywG6pdtg9IIVUQUa0u6KsyPMaA0thIfhAso+0CdseZqTszZjJw
3Gae3/f4w1dovEZ6h8MTrTS5lREGNgwZaeyHdHHJX5l4agwQEsOZ8ftRt+YlcDsaYQqND9EDYhZp
BHAu3cmbB3hjwyhy7h+5eb0soIStOaqD0esrPtu0dNbZVNJ5K4vKHgPep0vh9iJpCejZO1ZntMOS
tnOcnaNYmXCUx1tkEJ/guraiakXKMv+bQR11NkaHglIaOUEdD7cjAy6iEgiHbR/0SZmjlKb2zILW
baLleyVYp2f7dasoqK62DzPX9gVygs72I1Sijk0+vpW8I+01KNXxXebT4zobid84LJU9/biLqYSG
lOoqzZaVbA17WZiz1eXJJ3Cd0nJZM/MgypG0w6D/sBuO3bvDy0bnFz/VDqdYXykALPFdGtKb9nPq
tB4fq22osPMNvjQdNtzbi0qDrwYoxNxUOAkjgiIO9RHtzRG6KGYE4fyD/6sH2BDQjs6Yj4mAuE+A
zjvumUxOHFWGXX88IWivyZsARDcRm7TqFAUHnQA1cPrwFW0mk7QaGPifbJi1YN+37sCi/jI7h8Q8
bFSi8WvYsqfqkcVOjx71ID6GMTkkvIE2vtCAYQ9PABneULI6ZQTD8zACZD/y64YFSvYYeXhtr/X5
/eAi48NYWtz6HuV6MAXhwCM3EcFilbzmJAPOLIJyOJjWXiZi54TySVRvJy1jyTlo98kp0JbvyzTR
iRbm2QCe4oG9G5y2f5tSz9L2Ph2XQr8fvqgP2CVkrkubhsUHQx3wcCzISd5MLUOobdR1k40Q0rFD
6hz3FQGDGwapoNwu0fEMgtT68hQL09Af7p/fVZdR8JnCqn5DfejnF87YjYEsUvXx6OM5U+oS525x
F6WyLFWBwhK9VIEzsn2D45TWwnF+b+EF+f1ADyYd+fWMR6szZb1+KwK5YHP9lN42z+/g6zXXfG43
mneRg4QdFe5C7scLGMBX8jJmdLiT2SqYViy/GnhwxQDv43QDsN+J/jbgDrFSYhK97/2fXwU8morr
/oL94N3Mk+v/POnorYwsR+eBKbcHMXlSlNgoHOQ/LK49hQFUl973gatb+cmwigLYZzLudSRE+cOx
YgzyoDJ46xhp2SyM9QqIfnkIaflvaT/Wj//uLBCj6tub1WU8c33p6HInIwmEH9jGhmMW76u9SWaG
bxnvDGkFJm5X3MDhuCuyoodJHkB02+1d/rpQYZh5Iz9uvv03IVY+QVFvWd+mcT35QIiGaJbitlx5
pjruH70dMgnmI5Q99AupOtwX8oCyTfj5hIkRAiTMvZ5Ali5hKdbN9PdZ5fuagNJhPybO+4nxdvKB
a4uiHYBla+LcibLoq9X+lpq25f7SzD0t5SnqvKzAbz44R7Zu9XIBOtpwRiLq5LkHikOwug3hEvNm
hr4jn/4jNtMw5HcA0IBn+Gj0XyQFOX4KLFEVtKsEfb/ByFlf67XDhqgjrO451QwB0CFlifT0FLXZ
yHxOlVANdxbFoZ6/z0ru5n8COr7d3NDY3MAOyZkvcdJHf2MAYUruPbSygFmrPfGd3BmL/A6fz45e
yR/6+BDj11vjTGO1SooSK8l/HeT6hSkPBFNFlsFpWL8mQjLDGbyo4w86Zm6vPSmbZNy9xhHl9n3l
fCm8VwGTG2bvS25IjL5LHOVg4zpgQBqgvZDlPe8scQlDbRxIU9nHkwZPUsR1zrwabmGUDHt9V8bg
HHwYZWuTDnzYc8BS4MztJwB8x4U7hUSlqni8/3UIs0+ZEXS3O9QMkTbMMh3iVfxpgCbcueX5tJPq
nBpID1d/2psob5lnt334CCMLpVp0Gw8phXTEalpZFr9MsEr7bzmWxvDP4cGTzOV9cpbOyoBe2MQv
vHci8SpgWRsZd24f5Wm+OC1INW1Zy0aLq13eZHlAdLfzZ2f/IINqQY1phikUmznhKjdtO2HB4ETG
aZZqPZDb5oyneeTrD4DTRhT95FJdnccmZc91gxax/MlnZn4PYazRimlaoBfCp8jzcltkQaYJfqbM
HGH1gAHpUU++61bjtPP0kRAUDpyZqOpQXOiXEFmbfqp84022onh+xj5mUCc4Nq4IM4GMiihplKWM
m4xQ/kJGxPsTTEs3koWFtX6L2Fak7g/fUab0dKEhbFSUzQ+PsaqwztUHwWUehEPUQI+hIWtxwB9I
P2ztiwknn8TS3hxnOy9ud3jCiwutKq85DbtjiXQhRnDHBYhldYTvPoN/Ahw+wsxftRz7fl/eCc85
/3kdrq7yyJA666WivY1HksriEkCaU6C+M4yeLrdCweOMyIPkWnjREehkT5+ZtlPBOV2JLRSwT3Wy
S1//mvE16n4IAG2ks0fU4gchSwpBr9IpgcH/P+/jyJ5T6sOXnoVyBu+IgUnL95SMmV7+BXIvCbVM
TH0lkHzAwRqtemXKmBT3DIj3G9gEHbcTg5SKA/NwwPmtRCL2sLQPd/dhlr8X/lYsHl2OTNvAVS3z
vS2fcJhZc1gK4IVpkL53Ro6GkKQJAAGsHv2U+Qb7MiIP4eHqEZS8IBE9nckiMJJoujNEX+WAuJMX
9C5dHh6CVZHnXXIEdeyYErD8H15qJcbX4y9GVWap5ds5tDd7varMX171FRwO4IuiofcP9YM13pKl
Rdv22WrcBtWwTnx81z8Gl1i5FgIQQLjlLbcZFDwaBrM2Lmn4rGS8UHzad2a526OUTzzIS/CP+Hms
wWFucjm8bY+Cpz/u81VHmo7c/PHtNnLhHcWCcMTNzkHI/Blg3YMlQGhI8AMrZdP0YNkU+FzHcSmv
cKdjJwSWv/frBuImOXgb2/j/bNVQGyEzsoxsaeC82TlGusHUbY8tmsNb6Ckv2Qrnsc7xjiqagoQB
QwNCggbtYQUm+gt/hiNnHJehNlb02SSpoVxZfUt1nqnLKYUCSvlPAk1tijhC7DHf99x/yGjG8IoX
VilKQQCHS2dTsocsMpcuz60gVYVFvv0sGnW5jhsVXR2uIi1vNkUpqzyhlHvXr0nxw93lm+PlLmYy
9jOMHO58m6c7Sh+14nyntU7lMKo+3j17skVdrPSfX8Z6tDSRbOt0AVQMVZiun1L5j+tMVFEXAcV7
IMI8UYb543dfWWBcm0I39G/Er6WUjQEI/AxAi94+SV/jDiEhKgN/ddNLARmSo2pKw5JpxsAud08B
XlY8EYnaakXSED3woXCzWuxlmANFmVuH+chrDvqI16Nr6m1CaRF+pQF9yj1+oCzXbPg6W5XiXicK
CgBX/YwRE0qOAgxGqr3pF13S+AwS62Oh7fOzIxGf6Ycw2/I5Qgd70qqrkPnjWrlZrciBs+K3DTwv
p9FFPWwncMOrmY7Gy/rW7dKU62XtdK0k+p9HY6g6Atpi3qYgvO77Kjybnslp0oXbznJOBtp/G+UK
m0ubGVRRnjlb+7HzEvbFH+A2Qq7/ieoUV1t45SPknULfF3W9M+G8Cgku2uvNwNJLFwoFJO8tBeEg
k6/aG0LUPq4XbiuIEXvyVjsoA0+Gl6fJ66E0/Ky7IhBdMhAnFydigISwCKr/wAvObOyjKjzVx/Ga
ny/Y3t0tJK9OYODlPNDypR/PV+omq0gVrHq78e1sPBAe336hOfS5e560sWSsgMzC2ydG4o/HplJs
0f6tIhI/TJfZd3SJP3EUTxzBZ5wVSPTukkW5899AlzyfHWONkc9aWiLSTsoxCsywYLATos8d0laL
qJFVp0JOY/iyiK7q7jp01GpR7Razh9L7cuIAt3p8doQ3mZ3Q+Wd8x1XvGzHmh4FnIWkWPE3c/+14
edv9Celj9i8nilzsZ68sLUY220pyAEiVla0qHY1px94+ngBE5zii96BEnpoRAKGWxUsp2ie/YZoB
kyLuluzC6YEd4subOiJMR5GeK+ah0uaTrnbD8okhVeWsre2ytdgu9NDeAAgLYDVPrq6OceWMrKB/
O5UN2EOGHrzWL1Wa+UA8wZwq+kPm1VmG8QrjOrQtAk8RRcp65W8sehVG++X4eycNyw9EFR5lDqvO
Q80WDSQtgdjI0ntOA3nU/jhfMC+POL/aCTf4v6rVOXL+3pHKmSObgY1aqxg4nnxLWCkwHskHs2aO
TvYsdNQb2qlhFl71kNb+2zbOZaauJS+EShWoeRFRECnu6eoP98RtPdj9Sl6Uve7IQX2YVJsBXAP3
d4AJpQDkyVHiO57pTpiueYnh62FXfG4s4G9C350W5kCIrMce1rpy82bDfW0zg4AMsNqz8nxZwx4Q
PtbY+ul5vK5wu5tp5hgXzYWHa5tPu9hcRt5XuSK6w3mqfkR/7ddgvMM7DmcJZNRoU0Mct9iHTvEe
AcjExhNSZe5D4VyCN+HxLqi6UYSBoMvLm0nq2JrcLhYewAGygXJdKIZ3bCd/wSb+9lNSidgYzwIr
u/l2ZZceJhA+itPVG9NrHPDxXIZDUto+ysVcM3M4e/tPpI96K3HtQ/XpNACCizmlf4REWPAbeDnn
i709bKiMU9JB93y/GgqfElb3uX4Y4ipqFjQMjRsGUoww0yU8fLFEikQToRHmfp//lmivnzzPd0c4
YZv9Ow18yOPEvGnVAj3vWd9PxZnSRqEl961pYSTXduLcb/sMvcSt9H12z+VYwPVsrNFCCyg0ob1k
3FxyNaD+OsLLKuo1dldMsIcBl34DPatTxgVoFkeW8hIE/1mAPRUBTcKmmj/tGQ5eJTTStx3qNKys
wCdk0w+fFZo2sNVU07FmHzC4ptmgRph/YWCGBCC3Xrk3kcgIRGmYTkcB8wpln894N7OC2kTLeJzJ
zZQkXbCy6XXBb6MevEVMdxe4WzBXYIMTm6MwjR1O6Q6nEbbLF1seZPjfLCMgET70H3RcbkDZKXuL
l+xqX2a+yiA/BXxjDA/torMyhowGNen3cm6XWaVzQADMJUtChjSISmf78Xkl6jTTGIyqU7CNPFkc
xM+/q7CWNlDrO+czL6bgfpp2D/A2msojpl0jaDWFvxaUna+V4mwYFwP9ZFvA5uxw1KZY0f0scc8y
Jj2AgaQ+/teB8Wq+whrPQmfKvy0lUYOEk3y9Gz9rsB2KZMBMHJLkJVJyhw8zL2T6mitb05QUEPD7
VKks4FjDoaoffGPDOzaYzz37cVvmKxb1r0Y0Hmu89vzGLMN6J1FNeHghC3rejqYNvh36HjFrqDh0
Bv1QfgeB02pHDHfnIX+oJWKW/fTpdlj2CgDb4YkCocukHD4qr5WHLaELtKtspFNjWO4NdGf5P/no
XYx2XRQttaBIDsGKIWNT4edmAknZP9TiqmcQCvZc4xWzU5+Xrrm6cW/pZWvprDTv+zaUXqfOBdey
71S9qRS14vd/bOj2K8m0+vJG3SMnhIpk+bGtnFfL5IHSVQecaBjLG1la0KOL4i/Y/9z6b3T+WmWz
4v+9A3bpbbaiZYw3QCzdoWs9SsFBGrqRGslEUIu7teMXhULKA4beG+y/9ACk5d87QOl9MBBl7itr
SC9R7Nd/ynFr7+WO8o9PNsNOyklNKdENw36SbXTu1duLuQkB1IcVPYlpwEI/dUagGSZpkAB1J474
/bthVKXw1PKbOpjiVnWNuOMgH2PM2CQYR5tG7aZzEBNhRQBKzMtQN/vZEJd1fqLLqo1L3FFTtBA5
malrZ6XOeejdWiwgLLjYXc3jgUiiZoAAPVkKyV6uAbA6UKAq81oV8thXqtxrieshGmAS/mBQCQLx
7meS126j6Z3vG2bnYuSvHlm6oNTAohXju2b7EFbFTjF+s98Xw851EgVG2fBAfO6PGGWT8q9vZAst
wtY6MHkYI3jTrBwZUAMUEAPvcab+0LMqhrDvTc64oC67QZb2xRAaFsPGketsRechw0CKyWKZzW0z
UJYGwIq5SzASTc/MX/Ap6A6eDdkOU/bQtBEeRCakKZe8bGGW/+jYNkm5l1tZ4nRfA07mtDWIflHg
WEcFhpzNnyjzEiTqJMGIcmGvtven/TgnhUpl5IWdSvboNWR+zRcayCbWjUD0QeQdtxnu+c2RHn1T
qLK2NXjJQg7Iukpf5i7OOltXVaEUnRRJ+NiyOIZyJ2wIX9rN7EWS1zo4aqoSsT+TpcI5SscZ1tYk
jcmcIxkavaMQDhYpJSS5bWVTKiGLos43NZq42alaYO0vbaQslS2qOf75Y9BCnEaACmgDkcmwIor1
NBrklYmCbzCieVigKL2VA4oVvGkq2IHv80GsEtScdMaALtNzbq2jZvI6lpFePbD2H4T2dxe6eQjr
/9kVxx80PeIpCrOTC+AY28KBda8OvQc9Fb1lghFxBfDyenqPKy5fFWSaVq3cVVCNvIyB12Y2Eges
njQciLBzx4hoUCcd6KAOGpueidcBGkfIPLTrP0B+PDhlppOPRh7Pm/aJEYdGqs3tKs5NnaouFtTk
5j2wmeWUZ90E9i+guj92j3s6HoO8ED2JJXbqO/vp2wo2cNbC45GgGqwYBE5Xk85WCeOmL8oFWCMU
v2jKLTLInzOspnpXoss8pquwji0Ms215dyC42MXmZfl3zW2EO+q1BPOaOykvO1BpGdzLT5dlCaYT
v5L5XsvJO7Qu4q/NTO6MZa9kID+CBXsGih6KaDcKBKMbeqwHyzBbtTPzaGBaxpzFC0calNgrqPF/
PjAfKrm57RO2+hJ3IRJ4lDp70jzq7155lAaNdg6JLN74mJ+zl3fTsULLJtVaCN7uS/YYYxdy7dGp
i8svF7TClTCHE8sU1shKX6ThheI1tvDoiByN93iNnEr2s+KUaY9TLfWLdr5dQT6dfLqF1E7LbRbP
fjKugwF/M9IhdsK/C6fjMvAiuZcRru1TorefC7677CbIXiRzXa1WbZMS9paoFDNt1iJB1CLjQjXL
Khd5pZtgKi9x991vJmwXeooYF5N12SfXTx7ybAUQobN4XQBS9nqKzs9BtDhGhJ2cAlLSux1CHy5V
0MolEqC/UO2elyUhBLt1GKPit+HiofcH22U6k+7brTkd33eHC+ChiqGorjM4k9c0IYQY/LoZvL9k
7MAkg0gpgCi35ZNmILwv6Ziz4WaboBETuxKFDBlSZR4Aqt/BiQYOS+qyNQ+FsrW75NdBjdq24kvC
mfmpw4K7RWSqal3nfQooD5bTkWrn3cpYZ2cHmsCcI3R3syuOaiGgAaEvJ/ZpsMAkMOfDEXLhZVGy
5wtiE+eOIlXRV1E6HsWWn0w2epaOIkDIa2JJhm2CGF7NU3o8amVF9tXMCj/v3yDPZ/cr14O/jgxx
5BJwmutLUAHdrrWOKamtJ32Ky4oXFsRfEfVqlPby6EjWjE7GfR82nwfFvq85ikvbJBhqeAG/TktQ
P1/tPSZhYlAsom4sCsGaU/mFA92R9fp2pdAHHiwmonpRrGPMJAm+6PPYylE5fJOTHom1WCnp6PcH
zmlvueNMqCGuip0EQVWM3lHWmzr6VJjOFGHMhj/pYvvOQRqtuG1dBn30b44jA0ipNt1VX517EaO6
7sHYUVWHTNTHveaTVmYd4DYcrZOF65TFRkIMqiT9mUID8dw/7H7YfSHpKVUPziQNiq+gvSh7jJBz
8Cpi0Zdf+4aQDlItL3DxbLzAnitfljPbbWnEz3MspPrn6MNy92J2gD8IEZXPb2Arzi6zKaSVzPx9
ClfDqOokaPJeVAWOZrIwvy1CLc0TwI13hK8Gbi8qRcrZrKc67Crszp5xHH8dhpV9OLCEjztORgNK
8T3q+/PaOn1P9tEbQwIQPuKa60GHwj2U5fj/wtQsRcYzYW4t70WDJ3fX6eSx24afRGOXoyYn27YY
dSRZsyanYnUKWN9Xvo3VJqO4I4aIzk5LvM7WzF5+nqjOaREUv/xWhYJ3tyRv0zsDz4VAQCuW301F
BtropUmnKFL9vLofUQAieAr4eDTw6qZLaCfAIRT4m92hi204+f6reYGDf0hJyCzaQOXHsJMRh0CU
B2PFiNdDJwZOkKOA5ZBtpqX4ZSr1K6BHuYCpYGYFr1DURDP+NbwIZQ83gfZ8JAMmk92zCZTSEgdL
CnWzE9mxwm2shFtISxp3y9uZrclLfSP6Xw2HdDPagfADydkJeo1Ui3HZlkUCbRGCSemUi9FJ03D0
kPmCzmtbL98gJl70HBYqb/V8bxckFN/BsCj9tY1VpfNdN9KXrRbtshcrhcKFhbqOaxnal75MSok2
bKomZJ8Vhzr/9D4BcOQWoAXcBNGvoJowl/Na9GLE3erEtQ2lGX97DNsa05UO3z25Zs7YCI4Hfbn6
cj+oAP20q3PqvMGKBHavlgIC5vRTvj7UjshafnRWo7zB3DB+HuxWlb7t1Uw129UHYq7VEc4dlX76
ErSlHKHpSpLkQf+PpQzJESXXYGwRp9wK4O0k4xTi7k794mDAAWcljb8N0ZEVujEwS6yXXAoQfWf+
H6yHFSImW50ne7fp61ZUWa4k/P7un2XdX9DzznFTol371EjrxRkx/F3vxYDaEQnmZ0CTcFra05Ab
AIzn/EUBfhrnZVYZU7V/hLeVTQO7VgBkNOSm9k56p3HDjZ1snPM0UuwJwKF+a905E/xP9vRLAEVO
IKgKP2sCn0oWIOfGrcwElqsdbRNIBsyTaeiO94wk8jRKCLMOBJEi93Wccx1lr2wU/6n970+9GBLg
zWqF2tJFr4OJYYF8yFmdOrsddFKxc/gCvd1JLXpDPA9dVBur9YZdKPzvKJiwzb6GL5dmMu3w6Bw2
AdL3rQH0Jbd4lAIH5aGO340bOvX1KOMK8alwSr+YfxCvFNrmgVzPlRfZPGvpzpAh7yZ1pdkK2jeZ
Ab4t+bZlLoWLrqAGJ/DH57UNfTvcAI5gXhLnY8XptW7Lq/IJ6RyjlWGiNUM4+J6VIIvGbbXhQyYg
MKEPlarKJkJqPKoyAfIFnM9UIRbCILtrMHG5Vx+fQXqAx9Wr3fb3zd7VuPeHaWkcowg277jX5vmE
ky6e3Ma2s269jFCKxDaHWB8HVw8ikAlDEZwNO7j+ZEClF9EdGhvYOIXctGPitbiMobcnFn4MT3br
WAyvWa4JGdXITsKG9arAgcmC3obuHFhzeC8az4noNn8myNWPZ19hxxlBPwglsLYB97qEHbO0By2H
uu+m7StiplcKGSPaNPlF7Rf/SNsqBeEijLbv5QNigkntSMK4JpVDBzUq4S6rhmvXs6gsQgQuC9T0
bUvAbKZ5ERa96PW+M/7Q94cBwQOulul7uK15xJaY35W/4tw/BhOwoXycTF9k4n9bDxnW6Rlj7MjB
ca3JZvpQlKLE2Uzf3oCzyp4p02sGTToOFwt2iNdR4O1Bundvn8W6PaW3Mw6C9lWP4Vbvbb64T1RB
f0PbujDnkYI5e/9etZzZ/+w9t5nQvctzpx9/aOV8UGEhR8upUw86ChDBQF3Q1TlqZTfsExhLXw+v
FCyo4HELh8wLHLKLekit0hVthEMgg4dBl3XK/fIPSjKAko0kCdareYRf/gYBSv9XuTgT2txT6WYk
ro5Bsyx9euUhDe3+I0xdrdbLRbfYFQH5NB39PEmsV7SVtk6DZjYRrgECgqZr/9+EQ7diXKEed9PN
n1DVYGiQNaNhY2euAE9WLpDAZoKS+PAKciiq81vPYSw6M+tFFl79knyNyaWHrzsXEvKhGK8E0mkO
O08fv3wJGO0qoEVHIvxwLOO0yLhcpPAXBZqPPynhL1gy4D3j1tWjAb48U6bRGdALacK+WN+SgD+6
3JneI05Cc6rWdU6bN1m+Lf7zKSzAuKUW22Y89XmMD3F2RvYKnZ8CcOcjXqBL1h/oiukuwkigr6SU
zwqqKDlztIK4g1jrS+t1KbqWSfRBHiOWI/D6ayq0kmG0BjzCjHABo5IyxXsC+exEe9fNhINZl8Z9
TxRzARXB8gBjZBXIStZYzPAJu40ATaDltsxCHoinlyjtPPpJTJ1ihkaDgD/KgHZoYDwAaPZIwgb7
NktSBA1bk2dESIqO2aM3IIpTY5hXGP5XQG3MMub/7YXHdl06tgyC+3GPJ0bfu4P7Ut+vH+RK+aXN
SzxxrDafakE6w8NS0iYV/r33beWCajOn/DkMBeEYmRBTzId3zpKteg7aHTkZpV7tj/aCu2fCshfD
AL5Mcigv6SR0cWmqdJWSOv36p6IhrIPZ9SbhAI5dIFcM/ZMNRyZ0SEC9iHZM1PXyMS1LIRS69O7U
581ex2oBAKozfCZXnp8/1/iDnuOuSUr9hG8jml5twN6fLwzREg4t1sdnx/X9BHF+niznQxpoYGf2
SpsXr+l3xaifsBiTCe5Jt4L10xW9g7z1K5EdBJAzrEGwhxzumk0QO/J/yAyYZE4mNgWOvIYmzSHt
a3DgGcBvV7y79RsZvZ4168+QkbGvQgO7DTB8lkN0Sb2W4kDz465y8W+bIEGsVTbOYsIuDqt4hHM+
XpgQRuTk5uLFEaShn+z6Z3ZnIjX7fdxA8BjueJvjK/cmH4GHkiKx79/1mLYPe44I+3mDlOaePIy9
hHD5txXVcb9lk/5V+K3+ZOv9V5jSxf5QaZJu2pKWg+udFDF8U6GZvW8zHhe85OH+u4E9V4W+ZwlG
u2shr2dmc6zVByu6QE7AODyZf7YtWuuZuNjN83a6wzcnurXdjn2iKSOtGrvt/6adngDpn4PVgrMT
22z1Dr8pBAws9y8eFgs3gNtwiQlaMF9Y/68MuXBO/Ta9hxu8tScPmum+ZyRhdTO1YOK+EWPmVX3K
qqUt41KJsrUafscLTsWgZ8dn8zRfbK2Lxf3HGsn7kxd990dQlD/PRcqvBcraxvgzmXAqE9mVb7QD
VNucGjDFmy64OVsdPbZoJD7DXhlpUqr2LmlVDrgA6yMB0TaMSuYa5ahPG0udGSX2UnIApwPDKYCr
Ip2FCwppHeMMIdpDyUP179dBCnB6jXPyuSO6ktvSNMl7+UDHliMT1lM4nRokZMF8//Nqi2fS/3fL
CEXN1t+bX8WLmcKwvv8XI+Guk0ZNkGbzNo4/5FMBuXko/iAsR7ZLiBLmkRpv5NMFqK415i2EfwAT
fSTAK57e4cHts/n99ljJIRHdVnGY2aPb9PPhL8wQLIb3UoIuYTVw4qds3XSOSXmLQmrOrYP4s9Qp
Byf+VdJgzhF4fEN6olP4O1/L5ULY0Fb05tnraHJHm31YU37YpPPeViVv0YChVuejDJiDfyjZwYK7
f8QhxoMfJskIEioUMNoF1RyGqedp6V0KWcsb8nJcxig91Fy4FAnYkm3ZKN1nAeoeKhptQcVEELQX
HSkw2WiD7c73bmVuynxIgEwnaYJRhlHPK+rjx/yJjh9Cb+2ep+HH5VPxxkM5lb10qpzAbpoAnL0M
YoJapnpJ7ANCWB5vQoDJTEP1GNJBFlZZtTuJ8AkMqM62XQU2QvhkWBKA/ehJ0J9US6X6pnnc3j1m
MydD9EgUv4R7HxU+DA1A8bJ+bVxrVEojq42Fv7G7vfrFQirLAD0MroA4n6NYEnMWyP311gBsqux0
Hd4jAmj5SyourwXcRkSqyhGgypG2zbXzO28PLiOf6csmmO9WgPyiNvto39NJqVHwMBUI+ZI8ggIX
p0jObHgCUMkKRyWZlJat8bqwuYQTr/EEubt9nbtedB07lHPAlUsGE1D+H4vWxS+qfevHpy3L8+pO
GabHikeaDdD6p2FSmRV/8deKRaF8Dacnzachg9emHtgVgdL8DF3bL/Da0s8024BUclRZjKN10afC
nxbj3lslZ4yGCAR2fOBMGMaPodz6NLbBlL/QKwcQWsed3zSTiu9RMs75N5kZmiA6E31UxukKqvYa
6bL5RPSMWcNe9obTagvoq3xnjY2A1UCY+N3MXmPQZ8QxtbdSiAMecsVXsepzxeSQhcEnRuD6qrvu
8rtfycvckMAoejjtAHIqodVgGLQU/h8jSs4+KeyaVqkbltoC+eal2WpvTC+t4pP6BrQ+C4tL7IYh
hTuYlGgbAFB9rK0AAz2HILdRwwL/BjxKH7BpNwAqV4EJy9HbacPKXKgct/dsq/7zB1lWeFwNnnHU
UOKwn534DD9KQ6Wdb9Lejx+WV/FUmorxXWTGIIGaZD6r1FWI3UMiusufjfCM8e5s/asiD/4tYvxz
3HMiP0XwsopfoshGo1d5DBjKyAFvPcVErUBqN1D9zWDy9bZHfwTigO3Lts20o91kkU6KCBXIKOrm
8cbkSQ64fo2eHRejUmQ+pxn9wKnPJ+ldUJ+M1qJFjoCIM/yt5gtN6QTEoWC/2ArcvG+ahkmWeRGp
2mu5plIkkIbraY33TLnOpCkYQmFCVsR3L4ke6X6U6gHlP/YT3k7x8TLN432MxdRKgjFlyCouVHnA
CAl5Nw8Blawn/5oNLrRYveF7U2ZwmbDnbrUgwNeqN8//8ytHOkOzaLBOBVmeCzYhL1BBtjsuCqci
4DgjY6w7iXES/T7/I3OEs//LeiSEWKxlzHNyGCUBnUYN53gs8008JHp6PPCX+l6HRLxI8U1nuLDJ
lNP2D1/qNZhDO//m6psk1bytdcAioh6D6zd94L3H+NtL5c+yoz+aIF2K/+Vs8uVHbpclrKzKMdb0
rUUH076FaUFg/q9vzaMaKLr2v8tVwynEaKSIJfDR2k723O4guW/lzi/4DaCmpIa7crQerDB6H4um
XN2v6TaTqjbWW9QeEZVjZ+Coli+kenNB2MOAEKr5+3CRqLWcHKb51S7MLibiV2+gHYUDox65VQkO
1mTYG2QujszCk0xatuHP4e+ciKvoTHKJTqynklSH0GVQPMSVOahjg4AXgZsDk4hW2eVEWTcV9FSv
Mk63WSv5nj/4/wGIWJFkh0iaJ5UE8QrF2ryDo4LhSTa68YoEcHXHvg0YqBlU00DJ0YKsa9Bvhm7+
LXZEWHvizBecu9VAAkHwy5CErY/P6JL6hw8WVprq5jy1cD7NQEem1cEAILJyz5PlZSygd/IgHQas
Z4myPYlY6GXJPNiGGJDVQQu6v0HafL4FEWk0Ov6ZeAYVoo/zfRIIdmbcwzmDRWaHXhnktkXaOgRm
N51OB8uluZBclgbs6pDmyyjkPnK0BIPfwWnTuRDhq5LqerGVoTVt2qk9xp7s3Fc4wke/s51HuAbP
yqqVLFXFaB78ImOIMWbzpKn+lYq3/eQ48C2d0n1OrNnkLVes/FIRtGOKd2nOX+ufNqdB265WoXNj
Itdf64Y7bdaxoTHzYY8CEP7UGySMdkTKQscXMhsDCd2bAKm7pJnooa5xJP1Jwsd6JctBslkZj0PP
rpYCv1x4S/7FTM9LUGrgXVHN+3L0lK/2LXfV1DvjIcjb+7ZSYPF2p8szNK+qxI9orgYKorZcmpj/
GdQ1CkIdQI1rQQ7SLkm2HlVXdlC+QgFZ2lskmsOkXYo1VQXR8Y0VcmZ9CEajH01xPVjsztKmOX0A
oszfejPrcFhm0SWnIgu4IUXgZ2XlYRjSVNXu0g8cSbvhvjWyck5vKy8dVVZfKb1MZdtcPD97eiyd
JO+/pVAsI3yjZIlVcimL/Lf0M2rhRufXDPoXubEizcnHiFMZEHSOuKNGZ60j7f4tjQ5Z7ySp2pgN
2PCGKsiD8gFmxljfCnGKQYEQJPKmFJYb3stmYkk54e2tjx8S+1+hPRq9fTZtBGfZl7QJ+OiB3gwe
+/p1XWHBrtoAglEx3sJoAVLSFW8LxSVtrzOB7PoBQ7HAADuLEY3vdjta9Ta3KgKdqBQYwXssoSVT
fCQXLV1IsYpBW6nfCYQS5yyQrxop7od7OKdTnbQfkHIitGcL98i48m+UuZyutAmBy26xVq2sK4hj
ZDPVcVonxAdvox0bG3EMuj6xqjFqaFa98YMoe17UFzmIAZFphd4HXp54cRyg7A/43ssvXBbt7oxI
qHJxuLqwW0wUrw7uOafj3e9+aQC0Ce6LAUtsrBXqTQzNYCKfPI+kKGIdR+MkbpLKWwwK7TG6HLXB
fZPDO7vtLiX0HX0ycIADBlNbT+q45ocIYw/Cc8DQh85UExBPCJiq/1fMBZbH9ch5iafnvKHpD+At
HKrZGtMCqPKQHjrpUxM2cDh7TD4/NdgvN5EK4fMzQX1lv9Uc9enQLCHnkx7S/EJ/WTYMASS/T0br
O4f22CFEcw9BuKSRc4Xz2PRnLu1Es/kC6WGRrTidLUSxooXps0pho+Bs4+yt6Vc7wbKVppxAHrPm
vsH0UNdlMWMrmriMiON0VcAQs8M98EbWz8TpnYiwtZJMiVzAqU95pxsVBJG1KLCc/NZHHY5lxfAZ
7wzYOOEzyA1bMSx0AQV0pBxjRe58rc27sTunS1xYpbgTr2oTo8ZF/czqM0H2V53RDduOZV63Gz75
76U29Lj1vhOxs1BDgowWxr0rJ2RPPNguKJNBa3JSlW/Xuqhji6gPYXpcV17D1TesusxPogGhBtdo
o2us8n20pY9LTBzYY6xSfs7P7Tl4rB1jCRKl7fOcU+IU0he2k/tS8SwzbhX/t/edPWAtrTwfAyPQ
sqMbnqk4f+xwWfJU5qE+Q+EFc2IhHGBHBjZiwOh5JN6XI6TzKATnQr44AmOXkod+r4Yfsp7UPApl
5bwXiOwxiv8qRHHHgxI5d7dHG+KIVH7r6Xgd3VaDTgO3tpIJSq3SicG22NaSsyfqc1Cpt5c/39bq
9MjjNZgwJxk17B9xc4MTQEabQNydpUsqAfx965Zx39NLAiD53xkC2IImObDAHvtowleWq4g5wy7B
b+FIbwzQnNUkkGoIw7nNXZHBR2HY4RheXIr0o4JRSAh1Klz6Z+BwpoZjPVhugZPxYtxPdwN4eZkU
GyiQtnoNk9W3ANQLD1sCnNjT2Ylqk+S2WSy+rlfKsiol5VuaM44sHI7dn8vCoV3xBjn2vgeem6QZ
7qNVZNk0kEBYdUaLsJkErx0biJXs5r3GgS/VT7ZGxvtZgY4pIw7JZ65+dztfZKS6EpK5Dv50hS02
KLdzm6CzZl/kpCJbpkl+SafDFpSzud9F4ozgyi6F4auoW/VuAMIwL3GKUHlhNLu0hXAI8+Qwmxmu
EIhCxni1px6aFsfdXGfXtkoHjPR/nzFtPLnRTDp6UZWNeZONnucR/eEjPLwOALl72o0sHc9hRXof
x4TMlLnnU0M7+zbeKVUrZu7yrX+aLyjKSLPTN8PcADqS3+eAau3J9POYm6h7+XiWsdgjwkUOIxNB
jD/KiwSw2X0I8gzqEELj3tYg2EgTDpnW9UDEAxG/EClewgdXEMDKhyi2/62DF9S7sg50/Lqc9emc
HqAMt49MN8E6qaXsEf4d4DSz7jcJ34o8dmZlQFn0YtGprt/8Iw13+/fprMAze8f6/bPTKvR3f3ZN
T5haMl2zZJfSjX+zgtTNqUuAJfFYoad5dKzDKwzyvvLQLDZbhf4s92YZWtR0AqHsBKuZQ6uKzPBe
AjN+LCrJsEsHVnHpb32Rq6mmq3mpypaD/keP5w97bVEPSsUbZze5c3htaxZOnQmM2GmsaD0DwweD
4lkgH0Oe3UCiLJWVxDtGDf+SU8doO6mHbuH00Iknah7ne8PZq4rnjyklncx//UlrZ0atSA8Y8J5G
3RQRVALk7tu2uqqpdAZ4QRBSGgnt1f8RQwLzVSum5sxOgKFubDtrma74GyM2674uMV8HzwO5cgnl
RbmYZQndpxv0s8s+GCILlfchuUjsG3uNKWJ+2YrywiGOkd7Sh4FsRzFdDS9IzSFwybmDS5CWdiGS
KrLfZPEwDtJTEJhPj5sbabvJRgzGG5i/L7tBaORlcfaq7r7wlLFltzlOyKBYf/HuaFeI5g9pJ5Vl
MiQsRM6r8tRjiPOhh7BJCwEhrW7KOTkzxRX31tScgC6Ap+ktIi//vNHEScrGy2r8nIT+6Iqjrv4o
hhxv9E3AGZ016w0qikZ+D81/lAt4Pf0nolgMQH3SwXJjm6h2rrAlDMsWDQpqFLpm+ZNw9h5OTzpr
j0Z3LXydzQ2bxNj1WbObFN1+eqRH7ypX/0Am9yLM/C1ufkfvPGWjCrZh9SfbqPgdWCrLto/1sMaQ
tviGs1hcZGLbRllmQa4sa8rNiKdsaO57dDLZNFyLstow5kRtxNb2EvwqhbWwIt/hZKYHy8/9T8qX
vZUw579Rg28cg1OxbY/QTmL9lYipxDCk4p87fb5q/09g9IUYInM7ADSTdgTdclvKfDTS/vbuuYhv
wXsVqI9Xn8Mqbwz9YUaKzry/0IyqG/e978v6pfY/uRImwfS0duQBKygBiSsdfOJsmVgyTGuhyY+V
GDJPXVm66Eovk8nG8/e2rGpNtbiMXn/0j72ZbS/In4YUQoQDL2nraSSVxNO3FleZUvIEHMnaoeyU
ORYMECOYRhIYCzfS6D9gFx4FE7jfLrJMDnJUtc/DsNdybrWZovdnEUJWEEpDGulfA/CD43yhEnqs
vrswRjeKTPKwUkKS/TvLFK1keqKCF4lHLHDKzqFrJKQkJD2mLsxdG8b4FscbIA2Htr4gey2HkUID
yh2HmCipXucW2iUYXoPogVOqeYBc9CYp45aMub/p/TYPARImS2ZhXHVN0feYX+frSioxpXrwwVR/
SyIpUfQse08GLBWPujTzaH0Gub3Y4kgtl1vO6rpMR2DDqIv74OZYBtwklFpHXJBTIJW4q624MgA+
VnahjZUEMVZXSu8Oz4mlhYkAH/F6N4SNjecmGlsUxJ4P309NZA3Y5ncG3njO2JkkqVQkNO4OibfL
+CSQ8I9uX+I6nNtYClTSdhg+YthZtwcAmL1CH/Ncyx7tUUr/Yti6Gi4R4XdmkqPa815Y+Rb/Ijpe
ujXKaW3NkYHnCNfS6C4IfgM8DIpReE3X+emHcvoqUkzA1LkfQPf50x+hDBUb1gIOdqOSC2qKfkJ6
YgRgoUQ1oEDefRW/zTCDn+vu8EcQHly9yj66MvpDa3V3UVpm4arML9+O6YmCfoWyFyE3K3BVFYya
Snjd6dNcS3GmMUjPQde4ZPJT1cb3ymCESkPmf/zjgOk4filursj9NHrKI+UMyye/axpM5w9FQKvc
P9ymHxzDPfmttpAEhW7TAnPqcJALqJ3iI1YJ0x2APlFxLC4/SKGi+AcHAAjTKRa8mNHpNnna1JVt
bLoH8SvKAmPltO1TKNHiRsbTAVfWA0kQhsv2pFUYM6Eb8xa9XIVxhCFdrKFMQRJf1H4kqUcaVM2E
tuppVy3i1fLvjkKibId5D5mtsUK/014uxzrG4m5ZWbGnRkLyyAuJb+J70bL/Z7gIJep5dmWzr0He
sWNc+KCIVhoGorEPyT2ApFHjl23JhUiQegs8r95uCq7wb+ZgiNoSleymzE8xI6Yt/78kKDpMaAAE
yGOLzelO6CYkSdVL6x74s+rG6gnRknJdXRABh7+BPzwPNDhpVEecUrYZRyG9EU4aKFL+x+HlnCue
QkKrKeB4VH/+JwvcnP96TyTN5EfGQ2Ol4vF+i0IJdr7cOVXMxiDo7bFwG3A/4v4tqcrnuB0o6N0b
h2N/7KFQcZbZlARGszQ/cM1UEP3JlqzYqjAp2m97pLY0LPqWTZTTlW/nCOCnxa8GrkZn5wSf4O5w
eBwqeDTRx18hF41Zap0maNWtr8r+ZqNd5GzENBtUV47ZPgwuoP1T/mA7nL4fYlrlRcbXIF7ADLhd
xXSgb1O0BDNvEpzKdB2E1qq/PLNjdHmhdTKiOJAHnbNjdz8z9uSS7T6zfR6aZxG6j6yoiiDKacMV
qbisDhIewUqhexb+q+NdifOLIBEfpMHXpoCjKqaKqBIng39WNRxGq8EtJujtHi5L2HM5RiLY1Qzs
ONHpytw2+sJHH2SNp11GA2OawqsCiEpmgVc1u5f3BDYQBVrEakyU8HRbdAg4JLDFBbVFezmDLvyf
1o3tLDY7POZMsPaJjc3JJAPQcayJSPDh2HvtUGSpOQXrrNi7p0jOEs3efsOejen5jtC6FdM9lyWN
I7EB5byWTVtr2Z/pX1HwRTHzhxANmxdFyUySyn+AlKRZi8Yo+oF88Ri06fs+IOT4myfgjnMQvRCQ
gPQaTQ/dTz+0OxE3C2qTzA1nztg5tI6tHNIYpuAWHS80f/kxcVIVuM0e0qrcF75D1iR18yCryahF
ianDxgkYe/ef7RDyjTNaOlKiXScgkrCHJK0+brjXDAdzB9R/fVEmlMnRLgZTvWK28TA6BAGVdChr
kBX54SMBxr0awuMxyZfYuR6a2bnU8aS8rVIYvhtGDujIXYKvrNKOZBa+32k/uy+IcVukYsQ3rTFL
hAAbzI1XDLxYgTrq28esJTUFCnbTOnlkdi3a6jbPcXzKDRjxnQjtIlX0H/uDAJ8HcLtyvDf5bNdR
BnHEuF2qsN3y9hz71fnqzq7VYAM9+VYk2loocvF1LuQWGuAiEjxdREnUIOwPzT6Kk7rZUDtwgMXH
PZPFK2IFd5af6d+V8tEeLjT1suBB9iiUhg4ykF2uGBNAhkUGM5VOfC/Tgomswcv52BFUePVM4reY
XoYtKbPwKatx6JUT+NMC+fJOVAeT6KZ4/XoIXYb8G5N8BaRVdnkHSiHAWwHykvfD4UaqdYBuIzy4
IyYAWCFpLnN75BTYo1t+urS15X1YGwmHuonuYQkKneeExDBCe36r30FzhwIn5NAtQNbbxxrECdcX
lEZ9NH6uw798xIqSPtWEWr2EsNehqht+Zfsm7cU15kDGEbvJBgG2Y88mUCuBNpVLkpT5B3WEsUFw
EqVh5n6vq+HCkwPGOfu+JPWrCociLyVsQNDq+l86z24IV9ZP2rjf8h5epiv+TpXxH+aYeFWWL6b7
3nOLaqeXXOqmAkzPWE+ujWQmuAf7Zzjgvp+FoaXQgox2gdfXRXzyfbqWaK75NuUl2/I8bS65bCXt
Nv3v0jwKr9vVCMXzyl/O2MOQo1OqEq8USZ/nWhhQnTvYpSwEq1kmaruFrpy2jQ8thuRGNU6c93+k
ZSQ+nTtfcLmCg5zHdHBysYfsVA1cA0pAw2tf0knzReezzEjVRkCoGmtn7KHNLkLGlBez1iJ7o3AW
rr4CfGAiLJfrVjOh0XsjcAJW/XHxXlpoNNJMmVUOFkFfBUhTapXNsFr4kycZji/CqCnHgT+6mvMi
Rz0DYBawDxtpLtlpdv6AiLJ8jN4b8pYlC1wBHOjD7Ts2S6eYnhE/0Xo10ym5khOYYTDU7jOKVj02
2GaaZzC/YgcREeN0Oy8nFXtREcEXs40jehzhXJ7sHZlT5HmWtjtwZeSSFGACZruXT0uClVcrMnqD
5cy6dt6yM4f1mISSo7fal4yp9jd0zkZyCH/fG4balZOYq5B6EYQZIuc1PNqlZgcQ5kbF2Cr2A108
PP8MPIGKZS5s4z6XtRflisUbxjC2oseYFOgcJ62trahNzmFhavMeLgzy6YV29wWEzJYQOARppdCC
E34fYbKC0xV75m2Yxi1Arq1lTF+UPNUAjabybn5GKmuhGA/ZMCcq6lQklfCPC0cp+1ujWxl1Xnx2
RQWH6GzOHboGOPW1aYAb3y2qRGe838WSsDIaJUhO8kPKMHPSSyZtm6nEtFsFtkV0Mc0qlAnv0K+J
ovjv7IsW7tJHUYzpzPBFl5EFSaaFaAIg5DYDbBK43dKZm3+lMPw7Z0ZTr607aVhudNap0Cl8vKYC
2JohEgWgIwi8JKItt9ZzGaqaUDMR6oxcia4wfLWRpW0/tFxxs7aq5cIdbTmiXJF6k/dvzAvAXWdH
WcY7UJvKcRMNxw1AkQyFheUXbqr2auGwbF45zYe/CC3yj40pS9F6sFJO8ZitlCpEGSNlqj2rC29V
0thn4G6NshFWswwzcVrLo+KTLO8H/RuZUu8joSf0BE3TtY0bIKYnR9sjwg1GvDPQ566FSCH0jepp
+oGwIVxw7KFPnNq6hic/gKBiF9qa70zqsfaZyYDw/r7ZTXixjvxV6m4V4slZZk0VLK6u7w5mLmRU
aveVSUKpKUg4/D6J+winR46HqntNuUV8/Yv4jJ4azDbv4bdpfJ+0TCkslHovbHEsyRE8i6eg3MWK
WMuq7mOxeXRuIEwkEzWlMUupbhEqA/fxSdB7d5RX7GrB1zNfO0/kQZ9kGISy2BmZ/YBFp36OpCDl
ou33jKdlwdLn/WUawOoDQJFZQoWgmLkToEhhARFYqz7MY0aAtrx/K0MNLfgEf6QFhk2IpS0W47m9
OLwNKiEo5rN+7ob4qS91f6Ks7cGTeaYsthLzxQpDtu7Ejlci1HFm3fQQ4eRVNbGmiAsiUsPxetc0
v6FV4Tpx2sE3NGROkKfpwrsq8Z8mRwi7H09QKQ6QMF9ASWnqxGmz+6Vy3slWPtyo1H9XJEjE2cQ7
IrOSna6mslEDGjtESqR7p5m2sbUtMpDgW6R/bWpanvJs0cHiRMLIK5j6Qe2fg7yA8jUYBQUXZJro
vd6NlmWnhGulxwjTstBM5tuwxm1jBpuVNvcVklIOnCUzYXBawYbr0SB8DTYJTVS6Hyx1UxAi/yLT
xwN7010NRNAJKvQlL3VPXRQD4bwRnid5T1OUP8Czuhr0B8C2U1ngc43W6xNZOIn81v22AkHBgqaf
qeZ9USMbHipBto/gFVhmcwh8N0xA5FxLxJOKSdgtmEfkbdHcXWTiap1yM9QR+yh0OB2up2Cm1w9X
XfbxWuZ/jBZ7UocLqWlLDwySjVxw6E/rQTmqlbVSU2vPZ6ozOyLBQGY0sR+plrk028UUxpDSd5C6
GYS4YoPyp1UteBmLYLrcZ93tqc5D9Zf2oojgaL1N6gFP8CKFIIQ3bF9FMYCPX0tH/KnwKr986gvw
DEZ3TA8uwkDnXyhuTBLdEdDoyeQZ282ka2R54DPehwuH8xA5ffLj9T/i1X1LTrsr0swj14H+UhfW
YZTecIyd1Ot3zTDIebgpEx/MyTqXolEwJmGZbWsQwstXzaVQ31adJTIqf3GTO/dH1PfJKzQnWyLV
tkQRobEbA4FKvW1NtjoAnRQFcMathV/gbfzO6IAKGknGQjsDGbTE9d/Skm/m6MNlwek2JKSpltB7
JeDWCtdSFOkwXs1ZYIc4Zvq+m5xhezpPxUCpZXxQM3PMeft/If/Y0r0doPWn1MvUwL5l1jlLlNaa
eTyn+OaOlogho3plOdjebbiAy9iJ19i3gvCp9GxJBvJKbrwcwSB4UlCGKGmx9ymPUXtBHOQFr22p
YyrTpZhyhJ6/RL2a1iYOONi1X6C9J9NFwgwnCgAEy0CP7moQEwtS54LuU/sAEJL3ZeW9qb9gCD3L
q6+tEM4ZS9e9tdI+TM/UW1C+pOg+4FiuYJ+Oa8tB0sU64Kr6/KSov7Ab9/GEBNa/u3DvSUgwjXN1
IPHH9S2XT1BJbFyn2DwEm8wUry1amSLkNIy3v7udx+24KBnqAeN5NlALG59Tx6PwsU5jxlqiRmjl
w1Q65q6EJ2RSbEwKejhnDa+f15vJ/3KQwVmhsCuwW5kxvw/0A+teLPx4dI2JqF0llOOUBR1Xdui/
WofV0sfuPoy+kWpaC1pHPTk4XW5VExI9/n3qL352+9Zldpm2CSRWJiwdJfTLLZ5l0icrRUtt+lc0
nCzAd6giU8N+BSAW/MWxIWg3OU1apElgETBzuIu5/PbWWvDitQT+scuTNdM4++qg8pXl4Bs6PhLi
wXrvaowjsoLDUimbwrc1AOwna+iO10FdM60xqkhd9C3/gaogEvwsZbICNVnY9L4GQRY8NEAyqyC/
LYiW8lk17s2TMmS5s7QcRGY+MJP2vd1d6juelb+/9aYGEjSoHbG0dm8PgLof4BvP2RT9OPgQDTaI
DWLvQ1ZKK5vl19Fov4mt53P7686d8p/kfsBRhMmy/rbnoXbmpd+jBns2UcH0+UT0+kPix1L3QluU
vCSiIJkHVhoyFToElFNYqUZnnB4pDUFMgsCYpBDPc02vI4SHyu4lL+9Id435NRnhwYwINmT+5JkM
V8/Zn2bHu6DvoCiGv1Z4P/XL9mnNQ5G4IMHvCLN9XTX7xQAYwxHbz+Rd2zihvsu1IfXAWXF9eWsl
X7cc8//TcJ0Wq/Om6ugoXoCmRPnBWLt2rmh8WQH3BLh6Phbkxj2xT3SLImsVMII6E1/SORwIr+Qn
UnCt0QtOKOgklc7p3qd86A2sCVPdnJ2UNAH64yzidBarhq/RShppC1k0BKOLUUQSx8lD1svBjucf
OuY9N4MnTsMRPQzefs458meGWWnir0nRXO8qiK9IgEEvd1lEkBJFOF3MaJdv9wHxpIcpzZBS6eT8
j2DlhBhY7D/fzmNisFkBB4lfrNn7ETMJ6NJDQQzxgcJ5Jpc3eKoUeJ4JJiu7uFgRmS80wrIx4iYL
bzQAGXx2D3rb+7HxftSxd250AB9uK72AKwNar7VORqQ+EksVknTXywvBLluwlNT8/1JBlwdhL10N
YTcoyDSUszRDd9qTKcLL4AHBqpLRF1CB+ZQimBUezjyv/IznLxEb3e5+d1YUSN/f/LVSQQYZx/rV
D3TPvpYmXRKbBtIapquhMa7EXfwP20zPlAo42q4YBfmMrhHZJjAgXZfnLW4nHyAfzJV5TETiZsFI
sXywakQCD5ruaPHamskGBH+CI8wL6P5fDRpk+X/A3UEm2qW32DSMIY2d5wSvxTohKze6y55mICC1
czLDZYvZDZ25yKVOglNwD9t0pBNbqwvkuFwg4LZqyd4t+DcQ6DqzLFi9L/AwbpnJEewVJWb2zywD
tnGQ9rAXtbsgq3vDT9sNZcN6SIQ0W8ijZy6eRSzm66ZLrkQr1gHBvmr9JqTWnTinI8MRthhg8cog
ufLIbswdIlO8noFPEFMKmaPK784s17sMdm56bsO5hIZehXn4U3ZvCMzlRwkrorfP+lfNhd/eosGe
fL1ZIZ12aXoXx0HzMREhVywD6U2HDveyhp6sKu14tGnIPWDvcWJWddW1Oeqh8svm9W/f7qNBYuqI
3hgRVfpNH/TymU1TVpMgGn6o60zlmaGC1Sg3J5RDz0TC7wjM93R3s74HTUGWHlcOoUOVo7j3nTCC
NV01GNH4lhfXMTmrCfdVwa68ZuZOIxDRBZMW074+8NL0DBCAAcMd0dapVuskZFF86Ha0JGs1F628
Se3ls0wvFyLbtylYSFbxdWBsY8Bz61miCNgIn8L6k3/3AJNIb0M2EoSfjl0A6SebWtubRDfzNEtn
NtB703gFt852doZyM2b+/3I+NoVuxbz+0SNh/9Hf09HmLeChMd1eHuE3+1th4PfUm90fw/qOih+o
5L/C0QlgL4oIdKnEKd/jvMLIXcF9Jexz3QinL4pcmYVkpHhxLsoQ+MPLJYH+VDw6Q07pfTujWHLo
Bd4jQ0JpIVtodjMJxsSQozsZXkFuvMPBl/NkVU/R66PvS6GizSKKDIJkdIxFVtDK+3NthVPeBZ10
axMLeN9PYOBKAOTr2TGd96EoqgyVdQeDXtmsloTOyt3oaMe+YqZK1NbgsGv/+oFUpQmat9nta6Ue
GCRcGVhgcRmn1/kNP+eVYilNv3E9LEd15qYDHp83ND/CawsSThZmMVrYyD5MR6iiRuig+yR0bCxV
b1w2cb5rLLFKkkKZlBB4k01oQeIK3JG+zhmE0yOVGwsqrgbrijn89Zs4yH7Hp9FEEik5Bug8DB0I
9TdD0eKttl9AUGEQRZ7+jfTWdfR/FMyrVIN00SmYfdOBUjEBBZkGZ3sgSZZDNm/oci0aQ9IX/aKT
8pNhI1dVa04unhLoZGVfzj4poTkHiqtdTzzTD18WzrJkG6/4flraQtsXzzH4mN9DJVPfqZTM4v47
gpPPmIvdV49Q3gHJjpGhb46Vw+0XBfd6bLo60ZmNcxhdnQGVdDssqAZ2J+gXYJppxUHLtLhNcA6X
FXR/Qgo0MjDZDe7S/vIYqy/kdmNnm3L52Y+G3c0jFEp9JR0rRJ3TeBuuPq5egDeAa0U5FFUF1Aa5
4xOB1YADEeTM/BCdWSFnA31JwxtQDQZjZi45drTFYwKCnZrZyqgTwQ7eNh/2W6e1ogQYY31u2GT3
Z+QPWlOF4I5bMLEhfIzLTHSsfelr5o5HSvJ3S79L3ZUYF33RRnLdw7PVenNFM9pZxCk+tJoapX0t
87MTBYgqZ7f3djduudj8LML7vPhIdFLMJc9rWTAc18V8Evrr3/xS/F98xGl//019b5TiabKxE/jp
xyMOEOAVdBJQiwtwWUtRpPGrvLwKop8ZhQEy0VWrTdnqkGSW5WkRv9wM7StqVZ3uKM0o73j2MIHu
jco1Bkk9XbCNVj4R4CK6GtDaof6rD9AMwD4xX8L/yPSAcVAbt6fSWOpJaEMTarOkgCaHN3vViYWK
/EhgO5fmyG8ajT0QntXh/bdxq2+jsc3bw8f8V3Qy8k1SQSGeybrz0MzbQSLY95t82NAgwE5T+77c
Ccunss+f6nmZ1qz6ZEXZCnP5LoxNtdSWxSjDGd2x5eQoLalzNmacgh97KvcBD+Joj1fVcHB02YnU
jyAGUt9e6Nyjvadj8rXTOpqsHtY9D967bYMCDWunHWodJmXweFJ0J98x2CZ6VB3whsiv0lsatwUM
R0ZF7zSNU5C0LrdQ3hd1qX3ji8hH5wKEfaLYpn29KJZ3gUHCJOMweYGMmuFhQrOPdw/QHhsyg0s2
yFw1qBFuWkHswBSlfa5xgYOBtEgmR00h8qslxhN676LmsA3H8Qek8/1aAMH0FYkvaDZMDF4htYed
sewwuaOTRdxrSnqYgsnE/nymT91jVEmGv85gHiiD27eS+JH5lj+TnG6O7hJ9u4rJ3PLzPUP6trEV
+ptNqxjNRQfP8zb1UjrBM36Kri9CyCp4BkQe4B3h4d7/bgFN/hDlTt/lspnG25hrHKkFzAGUCLP3
qNh66oxoalmItQ/7GjMlvOZdmkklH9yE9EMeteS94mJoGiWzY25LTjV55N0v0vyR04ZayZBH5gkU
6Xm5NjbkuEq5KG3z/mj2yGl5+dVc3TmAud2f4xMozXYkCidFjNsIQch1upo3hr1e05coBNRV4hiQ
1V5ZYzLRKrBr7b/D624WbDs2iy3yjXElvSPWWP0lZRCuvQ8k1RFYk7DQSACrSpVUfHGfx7X1a82Y
R8zgQi9P9XxhxCjWYacYlZGgG1UKeKIuSDSeGs8kCx2cBC66/GX6hjWK4+07iEkONtDvLGPXcmVi
8AOUa1pnHpIKfyRFbXvfKvAOIJEZDXQuFDS99aztmQvz2Bh9CtZrxX9LPgFEndAXqi0Ix7YUzXb9
Y4JQv6UnWpuGfqXkojkOZGAw45jBcLPuVXQaCeW+hSLMYYBHLyGs3JNpXewRvA47OKd9mLV4uYWU
Y8dQgPWM21fzWsKQC40bQ8bL4RMSPt+u3y7NYW92TrWieEutT4M35+6Vtp3wNH3KzKg5XnqMW+A+
vxcySjs01jWbSFc8qUSFyccaQz9JQL7RyToUpHfS9bTNUfIUFzP4RbwyYGpY9/Mb2vM2suKLLYTg
qURMI5dchi0UfrrtcwBEGEB216kFp431vDqXmyxSIF7vCp4c8SaCcpzQoxQ0s5Qv9oYBlsG772ix
g//JKthJlqeR3qXv9ov15glBgqHt5pEGBPDDIP6jTk6vkHdr/IZxVcPwEqWzqpt7WrnkLCNrsxQx
pzO1/LxE9s+90plmACe0tWcYa4Tn9pgU53DRoCBL0qdorneI3eNrr7EN3S7vJH9SPkp/GqM7HhjY
emAhLEj1sMXcihdawlAS75MhBtgQhcH44xMTuAv9guCYkcmVm7AciCeczQzrb4ELeGj+xqRXw8d4
5ua6ZxpFzSQJjXydFqlgvfowpLiauBGWtJTOiyPqL/dKd2sUr4THmaCVxovu/EZBRvaafvjZwZfp
S9nuzTc0LZnUuep+7znFMgBtK+4p4xnknT7lE1WXf1zrawr2Na1/dQKTQa3jSW3BxaGiqvClxMeP
DWIbfcRJ9EBNcqck9Jm/2iydWAKvKj10m/yUi6zi3QY/chvRYr6pBNxesiWt5rdLpTjyE1OT7eNu
g4QVKG1aKvw5L/i+jyCNzGvhvbEMQ9I2qFZjmka4dUEF3Vu3lmH6WAO9FBIVxA5Os/FMJp35NgPw
JjEnxMfIOf4MWxR0n5l9Agsycx1lAkDU014qNKknjuzPcNSUj9RE5lJNuDnLKHmpx1M9Mft2RH2q
BvMiYDsxAZ56J+5Q6Se2w/eDPLhafTojjGMwigZF6kasSPjLR4+EHcbbqIaWYTD39iGaxoa0xxeS
Wlq1E97mqeH/iqwF2iHfl0tx3FhtgVRkQo7Ioa4b382ckuysjWdABXF0bXcKg02qLKUhe50FDsCJ
kCp+wzV4H4ATJFomM0HLR4jzC4BjKpSPHYAKa5y1ynEEobLbJaxXDBzBhaKXrK+Oaw/niPH/MezM
EzRotuMYweL5+NGLaUcuegeJFzXT+/yCm51L0ofyVOswbGI6N/0ug5ZEl1+taALhubFZlFYCj4sB
LK5mgcqhrsG232M4FXG+8j8FFou8zywvGr3vRG7EO5qlGd91AloKXqHuILo3VMfq2GiNt5AlBTod
FGEBHSveEMsaOcH01CdSrF6w26OHUKU/qwIR5T50FlyP9AZSg2pebHjbM2cbYyQmY9H40ZBRahxf
CszxQCgTd6a4mOLSvkHM+hfIkMg/kfxNn9CQ1i2FGlmzIl4m36tdtk8QJr0sWJJ2Tqm5ZO8SeU9G
AaekQJXnQyWqc3B1L+WIL+KOyFG9xiRTBlh8wRUF6ggcU34Gi6CNM5/ksiKRyMUrolX0IV46Shuq
6OFpSyhw/kpPEap02mjLZy45lHXFprPbPqjt8uQdt+8z+1WRO+cjJlGMwhTSARX2S9xEfgllKYjM
cQZmrOcuIzVS+gRKj+L1x+yyuG6Jn/NCC7/in3UTO+17ZiSgyW0wUbjWRfpUsriT5NlQAx5sRSlx
hAd+KAdsIwG9/UEaaHM3wEcNP/3cZ1C6uSUIAuk56++2soVzTZr/l9skPEsB6IbTCM0Huk97oOcJ
AJKDyJotfyvqm9CnIQn/LheG9KX5vhFoFA4QqS96+dMDhpAVxHro5e5iTcOvniZV8tcjPLJXMVPf
/BnI41TP1uRkRlxVOd8EMB+yXvVKsbskjU/1vvYoMAnjP+Sjr019niwsrj2n8FykZjLyxvx82csK
mfqMHWFY9a6jD7m5CfJWcBkdbi/Vz4TF7Ebw6tmhysKMkB7ETJBC0X5Pc4lJWlQu0Lf/hN//1VHi
FEqhtvOxfzIOxDjLBtk+ltpMFa6/gWqXheCHdUWpTJLI60+s05X3WP5/gU76PLA1/hIgpLM7RZK9
A//ySqBC/gJ1jQP3sTwWCworxGtysLx089pbAD6Zp30aa8yx5vfagBGg19BGL5Yx4JKZlWhYENHo
w7R/6jatR7h6yNvk23P50U/rueeQWc41/YVWUuBhoxCnrNdOh8JQtad0onowXASPppSB6XSVYraa
HPKUzelXwjbZVO14tGU5E0w/jQTvW91uOVuhke4SZWIDuK/sC2r3jI78Z+SwkWFq7C/1ympUYJ6q
2sq8bEaqX66ngU625Ig+XrtGLBpMpa8PwVpZGdF+UXHYrocgrIRPuE6qgTX5YwA+TmOKTVeVXhM+
cHxxxF4ZZl4sYPHw2SwMTzCzAH7td5fS0bLMkfxc4fqOuUTmrqeG0tRchQMrkkgQaRnBCxCHoUbc
c9675BlV0+6uCNSFQu1WgkoSwh08QfetTUpRtnGaJmiPukgVmSBF/Iknos+dTSmL2wnR3X4ToS1O
FQZwCaePLJJ1Kcum8TvJ+NLS4TTe8CjqksYKIHjZnDaHgw7RPUJulko7+RheIqJBE3KO1IJAXW/E
TLDG2U5zHbIk+ppICDdnuRnPSH3gyTjQi4He/PKXy2QL32z61D+JP1VAvJTIFqbIBBU5r1wnVlzJ
mlhxEPQJ3p7DCaRnRXKiL6+Hovdx24WlAfrUH+MppClmUDrbySAEJKRCLJCsRQLE7s2XBA9tBu+J
CoEtACJkGZiF74azDqVzA6r40gCatjaNJOpryVlV+DrM29iDxXlI9X78Bh7HFU/4Lw7IZ92yx4CL
BbgB7cmUUwh2IaqvtPxfQrhXmutiG6H6DJRrg9x3uBcgcVIeT9S9otjUR7lGVnvdpHD1IKmX5h9f
ntgczSG4pfKXuKqraEuo9thQBYsMIuDMpkvUeDogFg04TE5BmP/2kirN/PUvfbtlU4NGTsuZV9YV
i3gxOCiS2cOzmzAzAO/TKOBYWdrJx2asQFwhRCMjbP01EbHOTOlvAVuU5HSaHeMjNRXF+WEsget8
Z1F5/fkUvbRr7mONJG1QyuSJObrm0N89URBh19z8GBYhHR9wF7UeiGRB70GY3MtjO0AfcvRkujj7
Fed5+q8R3cy49uJ6HAOAc2rHVKTe6T8KImg9h9nWaA7SL/Y2bbYOUUmaEJn2rwm94IuH6P6aMqk9
CbX/tj/iki5FFOoDyH1ETsd0A/aQnGHcDwqBsixkirQpo0eHk636d/cdvojyUZg2jV9LanB34Izn
K1zIQ+XN8KWh2ccKWoUBUxyvpIm87bOmP+LkhWAMJyRFVPaxKbidW6E2Qr4/X3IBG3PQTWfdi+L5
qnWK8Kx9D0YHNUq4Yeem8DucnaD/rcwaAaYxAOZ8rph3fWBHzg/fb3F73Qhel8kd8B8Tl0nIpRTN
G/A31AMPw1Xw5ffc+0x/pCvo8ga+9qxDwwboGglbLQMteNS0RKU/O0C7a+EwkuPzUz/aNGZGAt4v
iI2/nl+iVtek3NJJ7W3nhHYvstS2shkA2F0QFb5tOPnku04y2Jew9I1szl0GB0u+BcEg/kVUDYpF
9RL5QPdzC2ZbSZtrrS6E36pxkYRLFJ46gwh8HYHZpzDhlEsu2CKA5rFRSBBbkyI7o2YAbbjL0dOI
9+RRZ4VecIy+CL8fDAbY7evidlBVO0nqLGXH8qJyPs6e2ct+I1YJLbXd5cX2ZQ9QTv7eMKZuuUc5
pkRF+jHhJqFoXqw1qspj0KLrM1imoVy/L4O6wiWCITM2XG4o9YXQ4SYYKHWeQ8gLkaQudsM9a0Ya
0O9Moy94barBTvTkrlu502cGJ7CAoXKUwGVhzwkXpvnsguNA4mFSXPU6urefzHAKxDHx0SyXQgc7
qQ1MbHKzK3kfUYMwQKCNVcreTnfqgTZESBPDETrXiP4lvdf32xgIOU8qjcLiGovwvkpyH5eH2hak
KdnV2ybz9Al8KbykDpgpCMLXzN25kIJI2biZ6R4kDCHPd+3e943/WimVA2rRCd/l4uV2DPgzrJHO
fl1gfXOgv8kxW7m5MIjndAV5xYQ/Si+tyryCqe58xU/TuCwmZv8vvWTWqLczNAgM2VZfHmiWCpa5
VzELA1iwin9RNPdjNxu0PreldWWY2OKMbdJafKjiZOcF9RgqFFWyFWZtLrpiKdru8DGig9MyIBQd
R1CmJ7CjVWMDOm/57kyzz6ODSZZCHr4SmnzHbr3gknk5zEsIBe473A+upsc0duLHJrq8sxGVgeAl
K6lgPXdVWD8GFlgiock7uqEj46lJl60E5T39z+W3RMhdNUUnbeQ9RzoKmxwL3JBKVbHCicMUWi10
8IQ3jnW8sZVhtQewtgP6WVi2CiuNmoqYdscHKNmuT9IaJCZCI4YuL8oedne7BQ3qoYS9Euai/k1P
NoB97oPQRUaIXk5hylWgNR22+3YKjA63sKS8FD3nn1BBGSS1rIaakMuZ/Smr8zXxOPOQkYcUgrm7
9Hv6c5Or9R2k3t9FMe210UkY+2bMv10k040/EjTe0ZVRPT7i+vLmaJQwch39L2n9v35wOH/2F94T
ZVgbocl0MST/Nyysnpyy7jFXkKIb0KZt7yveqacyyV7QC9UuVM6lPq6hKrZrfY42Smz2/BhvlCDe
/h+nHvIYQcV9EyyZ1Im8c2RpFDuQEwZEjcUVqsQVBVw0NDPcFMP+5wyUyQBCSELeo0yAgzfGTe0R
A25kr6fRe4WKOulKwMhuQrqSsphZI2Hb4uvK/yctaowkC1gYD/AhotiCVs2tjX2pDy8WfzXqfdYH
sNy2lAPd1knU68EWFF2GfkUbiZN+RjSgJzTgtA5v26lT5+bzlD3EbaHLLPJIhtWC9vO+bmlorMeO
PZgaAyt42cp69FxAhgdeSXxPm6Gaqp3XWhRcdsl6e2aXGEohQSpjSEDRkeGj2WjaXb39d+OQLcoh
+z4G02gR+zqRW50hq/JSgyNM7427HqiYS5K/wXso1FLoxB5/aFnxB6BQ8Ys969k9KvNmh3wnJv8V
evtjJHCwRBABZ7jG5WfMxLyz5Jy+jqOQw2vG6+Pp7Z3qRek39WDKL85qvVfeWvk3uSZr65Q++3Ma
Zq/QyD3A7FTY322XvRBy4t6F+mPaoHeg7JF6XeHl+fFbkhWzNjohRRBHK9cIZKZ1UsGJ8P22PifA
EUUbKULKrOIEAR1GlZ7rVsXWFRdD19XBEImTsYhLbkqd6kYgLyyOwl1JcsfUMPHU6XjX/nB2Y5ge
Lo6xkqkvGuCPSMvixCWMNUpNwJ9lkApMR62gRtYWwa9HPu2GoBvbxoKMbza9gn4kko/sFUvSwhNd
s+NrxZhbhDafSTCGAqA8VEV/Y7+H3s4CQmhVvwtJdlBNu7xYhGVMtSBAklQ8x8KvwFsR+/xbpkQQ
at0PpQxZFtr/THQtplG3Vy3s/A953NUez1C+D+WMcWD33sfTS7gBP/ZpIzeZ4+APXT3k4CaUt/PF
FEZGjBbQc/2h+2342W4nnyoDYOI5YTrjI5VTZNOiB3BG9Rcrr84PMMrYmEeTCLiMKGxPaDN5+WPc
pZC7aq+qTpuixWEUdPt0ZxVHI5AB5QeWQ4OOgAczEQIJuFGsVPVZzN9pvvUKmA5Y20hSDerZIH0Q
lKsQw4Q1zltxJFJugOPjoGGFSqDzua0dAmfm3QM41rhEIjywx01emCh4kGh4xn8QKxdlY7BOiD99
LbMFp/IAoXwbhqSN0nHF97bfGLHlj+LQwmsEFUSDoG4Q+yfcJ3dUg1oeIHk5hF6q///LwTnnTo+m
4FpX87xEhZD9EK1dOQHO7jN88U/1ZsJZQRqH9UHYNjfjQSsgX8CrvO0SMZ+fF/CmSm+h4nKkS+Mg
3ZJfs/tKSMUrBhHjK9iZNBtewE2zUl5uNL8edLmq7D51pzokyScQaWNobuPkAIgnl5n3L/AqdoiD
vTsqYeTuvmriITjy1thkEprKXKr5IsEPGZCNqqSOQSX/J3lmz14IR+X0YgLZSYPC5oo5371T+sm8
oMzw/3p84/C9iy8ygIrtcp1+sLbNQBObhlAOSjXif0R0zNbzB0HdTNewF5BZQae/73AuReeymjAs
NNN4554WYuB9cAsVtY5Zv2lcM9UDzBUmpuPvVirGdoxPvaP1eBBIDyzgDP7+7ySY71+PTN6L6WAP
WbAm2aBbmZUDVLuOyZjj9L3QZBM5cllwsxb/6TiueZRXFGAjA2zAkqoHFJumwsXXatT+HDp0bclj
rX67ugxmFwCPV7ubFQzorg6PxrA3jW76FNo89uyPM9tflc7SyAgoBvD4ey+g63Mr42ODfnTKwJyG
peqx+RX1T1XidpjnBL4g76UAXeo2KNbphGCONblKqafUJ5+ThK+zvVTeG1BsCYyU3ZMBLemq0OeD
YhCBp8IK6JBIlHRhwD1U980PJTL9uF8PZ7DqxvJD5Z0mZnTvliWv+zZykxyFb4CtFf6ocpDw6X3x
ZljALPrmMSOva5G1qZKUaUIWnLfmNBYVr55aLa7WGD2tyjYntTbK4q6KmkQkHSj3aclTZk965raj
TJ2wv33wzroOCvBEVzdnxWuUJ7fvcbUw+93fuZXtSc6O49YUhaw62aJVQ30EADY8EDA3bvnHSDJd
xFBZy9ZtaBiErp8TZIjtwcYeOMyrPlzaIihlXzlTMXmWi1DducX3HBtPkJrRd8kT1144lJJUixGD
6/wYSD/N9jh2+OBM/1WccHDi4PtkQVJVBP4M0REm4wCaGRSG8Mcm7Tks+gXdIEOr3sGeRENIqbWt
X+RzxDSozuhnarha1wcJdEVDwJFqsP3wsYq52ncU+dVA7YOOJtReeTweJQdf2kBxT03qwWW/J8eb
G7qWnxaRfFEVzEGvyBLt2N3CHGZfdlBAFMyLgF4spx/EkvxBnyvAralVAbgYGXRfvQEp5S7GMZVy
9Re3LZApj0mRqML4F5icTtpLAqwTtXsxh0bCAM8GTU+a+1h/gU4YuvoI4LYGDB0qcGqzkooo1L+l
3N/bt30Mog6jcEMDD+ujSwmLGBEiQ72qvBOHWWtOqo+D26yEDn2C442atoRjVyMs7FyUB506WaG2
U0cdcJ6i3BbTzCCmBl7Hzz3CyGuE97YXKdwudjHL6p3vqww61NzyA4gIs9GZlxNHmJdOlHlazPGU
zx8WoFHTFjzcNiQNUVLuVxS7fpZTCLW9EpMcxdEUxm4/pOea41lI/cHfeRd0fMOVH3nN98/wMNUU
Zl71G7UlYb++m5QqQqosMgRQEQgoyTe2IXLMk2q8/Nk7M9jYua14UylKQdz1333nwqr7Zk4qHNT/
3Ol2UmsCVDGkN8gpgt1iLzLEG6gLwsYdqseajVpUNKVVOaWP+k7UC7NU60IKxUQFtT7GcczA7+PW
ehp3Pkl5rabtuR9x5r6Gd0mU/blV3X9x5S+1np0U9gAuf9wFxJ4mJdk3hNs+fmVPbepsOQm5MkeJ
PmxQ4mrNnDM2y8jVncNmiTJexYwWvEreu7u80/v3nT26cJvKeWE+3/CJSe7nuK5ULNntQPUigCUS
IIKkKz/UIJoFvAqZZE+kZTKxTNvoOJ/JpGCd3Ad1MhpPLOp/4zCb5yxYnOF2TizQvFPSKSNW6Wxs
+SqZam4d3axhk5vLwSb+wP4mvb6C+WKgRFJCFyEOQ6Ob3+xOTzncbCU9XnRNwSJgpgWPXRyS/ZRf
jTus374G6me+FIbwsh9eqp7VKlhF00dVEZvuemrGjM78fPJAKIWNlmwqLyO6rRmURWrE7esmA5Oh
ST45hbFjsq1SAGx8SsAvEksh706+jOzJrE6DxXvN5D2f9Vb8Uv00J8Y2atyLFrgxxPWsGLm85cPP
E7DML9ZACGfpbr7y7glQQXZg6PewUldAVcyrYxnn1TlFXthYZj1tNsgc2pA/tGOXoUacijlYLaHh
FhnXTwCw/tyVjIPcEXQWf2flio4a934+bvsuJdnJhJnrrLrYcFht4A7syzloUoTjGywTQ+Aoyf+Q
1IyEP432cNg05mI1Ogr1Yl8YY/KMEyE166Gnq90HDpCmWSrU5Y5aMSplRvTPYOC/tn8N5P11wJi+
GBq9lVjDlbqg/25XSrHNuPbPJC0EaLQllzRbuLYAftfhN96yyTxaY86Rli7H6gL5D/O3HNhqH9Ai
agAj99lbuQy+29nqo90SL2yf4CKqpBDoPCFHI63oUBhs7AnLN9g8eM6jDoHfujysq3PPmgff4I9/
5N7ye0SOcosnMJnnOjjBiz3e+gFDIepi4hcvkf+eXWEo4p+1HeSbCGm2iEmw6Rs6GEYm6c1xgHi2
x6KIoBN+z9k8dkxJSmr5MVsTOMYQ2Hj7LM8vkuaxPZSN3VwO1igvafWaWqbM33GCNZUi6VfNz4WB
TfhaAp6toE86DE7JEwEQYkQ7soee+N2znQz0skb9qlajKB3hWCj4Q5LQBd/fXj4vfIm0rT8Pdf7h
T6vK99RTHo1RWtv3X73flHTQXp1nI9Hqq8Yp6h8kW0JSBrqyGoaI1qPvhf6+bHK3VVUy1NZEbOnm
R0uHaHB3AfMWIEbjUU5NZVPtM7gTMIG370zGmJwDv02Rnnge/EDs9D91u5yGq9nLQd6NTU4gkv5a
rEg2hmmHgdWYGO/HLZLilLdYpQTrpQ5Q0OORjqMLt2GUawcHK6oexffcrO7GO2cfrH1poI8jCdEk
5e8TGtv43pDI7erswX4L0g74FRNho27m9WizhkaUarVHKhidDkpOVyfTSx+NlJU+Ixp6WMsRw4kg
jV9jtEy12cpR9K5HZetJkxj2ZbDQ3x/Gdalk9lF7VQFkxIItxDN1e9Ye2Rw38/EiFcDKqh7P4cZP
xfanZQnxCsoGeLswHfkZeRWS8b96osmLRL7VhXqAUHv5Muvj/x1m/gtQGurAQSB7owjpvuhuMpIP
w3VqRjUI8HQVck+8pjyRcot9Le6QZULTtDghxM/5J3RFKV9PcaUusyXVgwMgVZJI3voc2xEVMCsx
jMSrGENMLx/kAG5B1JJDQapTJooLZHOMhVkMfRLDIlEAkp37Jvc7YzjVsUBKOGQW+clojyd8jAik
RsYT04kOKoER4TeYZt2Sl/A8YgsXsBVKA9NF1cuY2+bG1WsmlMlRzCWyF6xWc4EE0b/HVXgsrulz
i5v+9Zrg8MqcaOOKcTV408coZX5rNAy88IvJdgJllelCKWOE7yfBAbZ2+oEjXjx90doNpdlCla4o
1beNKIyTv52quomL6/sh8nkktAjbVCv3jpVorRqiFgikyApNXazlkjq9xN0WBakeAxyTwfBInqVr
5CCjvvSNr0izHbpnZpbTM1NcW2dfr9sJw14jqmVMxwRWXXOAx5PLIR+JykCNn430Zk06tr9ZW7oF
eFPhDF0ie9C0Pzw62nXOJedJlG674b0382vmuqUGMpgiL9tYtyifPegekQueLSM2fRMoxXyWxDaD
16zrWdlTXCEUwdt89RKa8zxVQ2ewxAtkkkx83REMVsw1CKPFHHi8hlqoY4CSuGmnyYU/V3fGwCX1
1M3svuEijb4ZrwVAU0G46AMLNYnI+2JrOzU4+aQVNibktwlcAewwCgFEgaPYMFb/hDE1pfT8VGEb
gIY2wt+YTACiFTHLrejEqBZ7Kb3MEu/nytsO5qAWmh9zTWoys80KiY2/W7Aixv3KGjnEhSxrliAF
KzgKvyWHjAbbhyQgAhUyPurZR4XQPt5t9aR3PHGyew3KaKlFaUmmygF5vTqa3soJZ27rf6hxVqBF
F9dv1vFZx0T6LrhhmwaHieFFlAOxzb83IucyMWimJO7mCtiaaVaUrZ99P2e5mrGHU6tnWV2VnFPJ
BHo7EthNrzudCHupANXgMD4ExY4DsdAFo1Y+hlABBXucoB1wSNINK3QGrZfbrSI4KXSmvYkDnvM5
WpkzPI+OnGpzFjXWZ08IQ/h/X6KEJ1FYfdtuBhHjpsigT9z6a+GRxGyUFPCAN0mzb+NVquEw8Lf7
t305YMZHFVJaoQ4zrk2dlP91+8qlZX0H2Mdsw4pdueonNPCoycVCqJi8Mxjbhp6ccqzvWtYB/4i1
CK4/soTn03j/8+cxrV+cn8K2eiGoWnq65g5twKw7UYDcmVYv3IIttd2XtNr/OzToO8Hot2DA0kZb
lwQccneCQnKGGWiR8wh651a9h6vcRygH4mzWiL9ZJ0kbrJI19pHeseBqOC5FFKdVlLoErzEBJyBk
Rs1MOt5SBvX1YpCnY1g8ea5+UrHSmegzkIyEep9ryM2gRCBYI61UELN61LXgtrOyqoRANTuLlJFo
nZsbywBQ/WC+LtDwfkAUQxFjDnCr6cKZkL23CrESrXDje6ZPTYkV2RTNxjE9PSWSK/Gh9085mct+
0w0NVs0Axq+21zCednakCGPyxVt+K/oz9wA61OJiDY/dZ7YTQERylhJJl3KWCojU/JvmWqO5A45Q
8DwxQ+71YOnph7PvjnBuYlSJxZCvqzfUpe4XNJ664uOZ8mjIHGAdNGM1+exyJ7i4dWE/SrkBZvOD
mOvzOmpgdC2bkYz9bd0E4viiRJ0IlYDI0RpSEGCNhPmsqg5MZabKv8X6JwnASkqEBgLiw0AsJO6G
k+/ax5k3Tw/SmM8IknP2rKLTZCJR393IObyzFqHw7GwYmLCXbRxuTeALyhzP4agl/hOht9rQqtfB
N2Rglbt+9lzW37gnALMSVhxksHF+WxQDC7lOy+4JOWUioK2az8bZc+8gZYJsfjSN/k3+T4W7XK8l
CyO9Y03aPyRbnrBbNF28bi+LiCaBR4JdAbuhPrNE6H/IKjiFpyQiq8h2bJMtjqkKQp8+/a/dnE+U
gM5blpmID/plAY7ZugqIxhLhqk8Sx1DwwAJLt4QrEipXXoMtnqEhX/Ap7GzLI2wuuMsimS3aPDMb
SwlOGoewoiV+MAX8zeNBCJ2JrVTnfWJFTNt4Sn3B7A4RxPtAW6JoSIDKxzh1VtdOOAwJa3KvMBa6
c8QYIDkRRkvL2Q4mBNtdjz70DkdfVsaFzT6ddfN92KJHlB2LMDjYAuaJArX9C66+4K6KIlLrflsE
at11li1CAwF0KLkJB7MT1DPcmcRE62ujbeQjA04KWh57odenNAJKZ6rB3fSXYMgRjxvnMc+345PL
auyvJXlmD8izxKiI6oFLVc6CSQW0KrQbT1OOXyQVzFfLz09lAY32oQqVrHpSjHRNzpcen1HJnjMt
/R9Ne++bTnAtNKFldNPxvJAZLH87SdsbwDJv7lF8iy2tM0UTRW57G1RGmJpRrjWp1k0NazoffMa1
qrOxHcOkzT6mXi66eanFz/urPterKcYhGaErdXnT56D0K08/6wWFKd/c5ss2Y0Uz75GlKDOZ8Hpb
lATk4vHX3hTJ7kcIt49QMnAMPrDU33KJEluVdyu4iGn/e22clBwWEK8+cDO/Yq+9TLBTp3G9jL5I
YSqMpIybdmg6uxdVdRwYFDE+j2+fWvWYKsoaifk4G1sfv9cortfO2UfyvFiowGjIjrg8Pcb/6RyC
LVez9AsWR/ec8Y65Cia8VCINqfCpz5r9W4yxDk4r8dDosswdgLIV5AfNZe+4ni7qT8tVsGrx1WGS
pspFh3xItuEo1VrgSiRxIkOrWvawSI43kOUY5jr6bPJhUVL8cW58zcuivKAOVWNduCV1d8SClT1q
FI0xEE0wWUVyDjCHwWr8xB4FhS3JudKA+S+EYooB1W6dyIdPqhkfax0gcmZWNi4yLm1aEKepyp7L
2De2ZB8+FTwKn/UiZvIF/Hct6WdI+/LD5BMYhl03fu8D1dROS19PtwVow3zaeoif758QcIAvdxMI
sT6muwgdR3WZ/swdtTMqwGnG8Nqsmy9a2R2Gy8MPi3YjKZywrsLP3YGZXmFLTkL0BVUolL7HpO3o
hKnmWGehFbilKL82wWf4fnVGRE2A9DWW8NcetDarRNVpT6eTnxOjWxQojf/Rz/q9Kt140UE4SQ74
1KP/s07Nuh999RaKGK4GRMbvUL+/pkVKEjH8Axn2L2ppdrL20tpIOl4UuPx15LIH8qw55yVds/TR
V0+wT0m0ScpkNAMVFwnpyLBT6SWi034vjOWJEyv7qpUaLy/MUDT9cfqnUtlX14HP/p3hu/kvmaD5
iVybziJlKzwfzQ1i4m2Pg3av5UunvWHqzNRnb4RU6QWevH2kYVpWrPWvsU00y42zGibAmQmwW/EZ
UU/zaEcFBluZfyXs1YjqksqrJskTMOfmULCnsqi35bqxMg31v9lkiGYHI0vkyIosFWYhO1VgOrjL
9AlwMr/0QV9spHSXa1Lr3JcNV4cGjC/sfsczSGBR6rhpnLvkVIInfmD5Kva9JJKnhVmWVZ805qLM
lY18Wdbp+OOqG08VYKMaymFwMNopGGQLIhruMn6NoFDHPHMmn/gdCZ27IKKx0G0jO9l3jSGgRq2E
0wgSxTyxuRGA98knJD0h7flfL5WPkj8nDeKMP6XMEqWJkGQwY9groYwkdq2s1GgkZg9d0lgVOLxH
eNVVezsUSFtVOu3aGidexSune4V0pjvK7oqLvtACGEISBa30qG3pAni07gQWWKym3d1lToLlXwgO
adYx7an7whXx+6741DcB4M6WhHmvw06IAetEIysZdb6Q+PcsG1hvweRyo4CuQho/lMyekB1lx/nI
5wcvMPg7CiZgqL9plbIrnwByF7loz+466sDcUP6SXCFdZc4wKjfFBnadUwsAATsy6ncyNM62/3PJ
Q4siqjFa54ArsIiQD0eLfMV2OE4lj/cQZ+MHg/g9UeCWkHWfcfgkfDcUqNb4Ua3r0poQhgTzaoUI
emqwVkA2ccC4i4fArLMDVog9c4cr9wBFC0otFNtJvi1UUhpQwIezueMnQaWogo/xv0vtuKuli4gj
hWMjRMMXBPkNiHqzfFBpfstPve48vWWHGeaLkoLTWL+22XKNte9mZ/fzP1tHZ3AIUl/ME3bLsIK+
6G2D+ONSkQMIKArj0nk2VnJ9SwZFne2x8ZMmHp93xAbpe3sVYkuNeiKKemvRJm7d8l8jJPXR93M+
lvVNcOWqH9bgtFAl/U8yWz63hi3h70dzhCSmOOE5GA9yxJPrxRxU6kPuqgSai2Cm9nJsS1+mg/Y2
YKGqYphV3lztjp4924AzvEnan8qWtqcNWTIb0rk5YWObHxKC4yIQxxmQk42g2md0Dl5V9Wh170EH
2B7Y7OtP+uHJhVmPFpJAHzQoR6T82PnnvaFulZeL+6UbYQJGkQh+0cUpLs2P4B9a647Cge/xhbxO
ed6T5Q4O01fxDJmJN30d4T1wRZbvcU1gipUPDZ12nix1Tdr9r5FqaJS71YTNw7C6J1p4iAoxE+C2
W8BwuHBvQBgzzbDrbkDo6CQeZKivP/woNJGXj5nsTVplkx0F3GfTuNlcx1tgSAALi5KTBaSsF3X6
n0eokYpyCYj1geebOcjitwp2vw2JajcP82D5KsHjSEZZrvgF5kNNYAeK77QIb8lxr/FdRVSSrmpw
Ru/7JDli8ckmaAUj7xdszYKMBgnSU6KM8heFW97uhDPNYqMXaCxeJin+/Rb3VTDAJ1OXJZUmO2E/
nkK9epCchF/LnVyZOM2LA+KJJwuNBMaxhnh8qk+AGqMWh8WS/3lyqMWdyddwIiPzNWyHQU/4fQjg
SjvYVjSZeIepDXhvyuKbHzK+Tpk7Mvr7tNQkdV0hlWXHE+EqRJChuXzI66hRYVlvJgzKh6g37hjH
o2ChtU6HPjij0Pobvty5d2gPR7w5ulJPTj287u8z+PsGvMwJelDB7TDNIwUQd46frTx5r+4ejRmV
o5Nh8kHLJ5ysq9ehmNin9M998y9VECCey7HJlA3cbqVbQlHQXFmPcaZ0/U1n+YdOS8vDe80I/9L6
5kVKAlP3G2XKdIvKy5aecZjbuDX8/m8u8BXmf0EXhZRgBKQRi8pOPPLQIY1ydAukDC18RHGr4Zur
MV2N4hpNU27rQ/OvAUk7zG+7szijtYi5FK/03E/ZiLNzzTD8+WuDdeXby2lOaPxrVd3wPAHmC9+T
LFwOPTM82oREv0RXjltwHLxGwao/Z00D38WJ21/Ub83nq/mw2gYmiJJSwmTUBCkmuqIbFHKR/KVA
D88wJPYxJ0pjAOqcDfRQaxQZFBFifbIIKlLg6DcGiytU9NyOwg8N/GI1zpDPrFGI/QyCrdq2J+gt
lh0TorD6X8PV/GZuWVlcjedgRHNuiMf2tNKN2+9GbdJ0mAFliVrph/rAjw/8kwIOqR6pkbVQApjD
RKJtLRyVFYqovSCjFbs/bu01ZAA1skGdrOuk+3AYxLrx5OoDGdKEXF/5D/2BqO/G/OSqIUMXq5dl
12kvfseHdBgZsiU4Vna9Nh8gVlXzXT8hIN00Xnv7TL7Vcyz26x6eAYtl5RYVMAgp3yghc0K+zUOZ
sk3yV1MxlaUvc4XDW6MdqNLL6JzpHkq0Kez7f7HTFab5EH/koeqsfSIrbvViMUQwpEt2akKBO4JC
U9KWfio/WX4/DHDyY8eQjwO/6b8poha3eGHlsuCf1XIvi0gRQXDbvQrKgi1OsYUtKL+V7QdeGqm8
imI5qGQLXvXN5HYQNRRFvclZoaKIasD05oitwJK6gJvugAHXjsyyaxeEJTs2CpLWmij18FcwkoXw
uId+3pOMXxa7kNBchnPcVD8imMLekBpZraYIY/NDgE6Pq5/sVfB8KYqara6CdrOhFtQNtYdyMyJm
sGTvZol1Q5ymNBTGMhuBUDzlT4NaJtpDhSBrcceJA68+u1WPMVDRgctyJ0R1OdhSgiu+EjZ+Yhnj
7wtBQqmuagJ97i7b7PGN4wHvIXA0X9rleY4UOk/OL3Ie3r2H1u+SC2Pe4etyOvUwoNtuBHWOtnkQ
++B/dtXwTdFt5ENdk+M5lZS96eIkxtj/R6VRoxAhP7VKSweP4VlwJziZYt0dwny4NLReOJOa7L8M
DlUjqXnURuy4WZTkRlcQGGC/raDmT91uc/j00EMyEWzb4dFD/RemhJDw5G8DKs9ehaHsymXOnSLr
/svpynzqSyFM9AuEGO6ZEPg8L0azqxK5KGWEhHUNE41DXJo6z3ZUrm3Q+QURxKe0/5Lotj5Htseh
0OTQz1a7cenTljGOlSUv/17bsQt6RtDqHWPTnfkiLTgE5H8YDH1FR8GCmTXaIqtHAFkygqB2xOQn
3lFMwA6PMFhAjJLmaI8u/6hYBI5fL73HLgB+IkR6rePP5PM3wpnGETxuO1xZNDP4BEYdLeofRHoD
LvGnDK6cdQCVSBayBAh8B/wMrGqw9y79OR5GRiiQrkGWDK44krs60tGntumPnFpmXN5//5jUtb8d
2G/XIo0egLovSEFw7pJTMYrIrq0vzwMrq4oxVv1E35N18I0cXjqMjCOyhorFfF3aV9iTK09qnfh4
ewg9zk8+Gals85kbECxtviT7uA3IG3+21ZDVeyCNMQcR2QDbJXV5bLe7DhpmSSQXwTTK3oNmpqw6
QVtO62ur0ln2j2fzM97cHrJat4TukmGFrHo0iuKYUVLIjjlpRjwsaYFfn0Z5sv/bpGdzy9Mo6i9V
il4Ca+gVfWzsNp2B6r2osouGRGARJFazj5NymSsXpOCGT9ZzKNr2191dDGLPjAlabgulHWR91tJE
ZwthmTtxFsRCQGesqz7jAS6mpxWTB2VRbth6lL5dFM1kpFhOdyArdKWKVjFW7wpvUbhxTZkB9ZNo
Wl94zThf+VKaJHhdM4L50eYk5/F7xZMCKZ83Yy+mhYg0PCSdAWZ/S0Y9teTB8ELCmGg9udMHvpMy
5OTW/IfKoKILh/sA1j72H9T8yKqozgd5od0THPyDpulbwyXNLJ+SZ6/8BoQ1kkMRgF8n3OLUwlGf
gA0fOQMkIcTDk6ldLB6ESYrvlAGOz6Z9LtqyiqBtK6Uokkcy3pgpeO6ta35eaQkB+9p0/1E6xkko
iB3hsPAkYI0N7mkCYHgfBpzB8Ls0JSJRk2CTUxHVflJu3fsiOWbDVnVQlsuePnn5giddBFss1VGR
XCleDlYNdAJvxq0jiRC9UVqkWAK50BnC+nehCKUUbQMveuZKVwjH9Kn7bdP21tpOovrXNCeQci79
rs74VNkuer4uk4lOiE3lKmWEnPZMnxNMZFVjomSMsvpMotk22vyxW4NyR4uFqtDmZcAetqpZb6L1
ao2G4UBlD4uw2duCEBGoE1LBRFuUkOacetep31BLrZhQJgmvpQAIdeHkTGg/m+DDYK/maUorLSYX
YaEf4m0SdP+tTIdoHmBoNJ76w1c9E3zVby8fi3Os8K+4dExkHyTgbOCmflFYmXb/EmWi2B0oVa8q
auhYeFho8c4ne21d3EKfH8TRpDz9YUFDsF30uNVjoNh1ydpIzVyL4/pM3wHTOQMn9jq42UKSceVD
4grOGmhrLX9uEpCJUCAwCLwMJ590LcoBMmk1K1AaFc/PfPXlQEyHtP3jBe6uVdBSe1EjpK8ChYag
Vu0S7U0iiwnGInEkEli0gsizCbeYrLdNGqgqPOHPMdMnI/SSXeOXkgkuoyuUC81JSUlnlrfw6BFk
Y84kdZrZX2GVOCl9KQKdYD7142FCkIKvhAisvMYs6LBBCUIzDgnJpwNaf8atRn8Gmu5To/kRjxcH
n1tuCCd2Pygv/CHhRINutb3qpFv2JaAsqhsQ3Uvri/0OeYLw9RuUBXjLT+UvDulvoU2O7RtrHJM6
QmQDXNk073g4MqXuM93LojPPghwvShkxZx2PKI0Upbt6J22U+3GAO2qk0mzuUfEbs1qMzw5synFV
Ywrapt82hz8QgZURtY7jgAYW90TxQDCXyNaadviKTG7RaUE2H/rYVYgBo9QxyUr1hlkmqxerBwBv
i3Nu0rVYXTmlj64QFLaS9IhVCcgcI3w1cpc0bhnwunzNJ+aATMmRlhAZX2CMUSPiib8RuFg3QcKU
5OOQx603cTLvYO3t4eMRU35MjrBJ9cbAm5HifJwFr8KYIzZDp5PpmRIuPgsqlvLM9RX3WBhaA2uD
arLm8uVf39DSfMytOHVgrNcU/deH/4/cVYK9Ubhxhg74uf0pdFfjTMA4JuHM9oPLx6rX/tJmtETR
0cMIlZ872XohZnHQvsCCrEHJIz/vUfD+hSeWCOAnFV3NgPzU6daoNpyyHbCpokGSo6AWKh3sevrm
8eMsP4AeKYJkl7o+GYSvYICCkCy08TfTqRa/FIzw9Eisr+2/L0BxmPhKs2h+2rRDXlkf7lK1fiXi
XP2fSOulpQSB7Vd+l5lSl63BFeK1j9XLRjS+TCKy0rFYcRPpADiYbckdNC3GUiv9tmxLzFNuCgoQ
c8KXNejIK5ZPlSj9OjP2UqAQ7A/XVxGcvXZ/uC9sS2TA5TC631u9yYSGbt0x8KlQ+3oyMLe/k8ke
byrIVRYbwlTS6MT8MI/N0MBanT7xSwwDTIAVc4jpoI9DvJyzmCHa8DCabIkEO7c/jxf6lajXc3WV
l6r69UlAR7XwYA7Rg4tc6/jsvEFQImwXBrfcQoeocNG+3GxhppgClp1/D3IxCa4vWBEwTYH43kl/
+MVL422mW0PbK/m/E5s96IRJwrthZmcy67Ky8VAQDY4w229lw6yLXJal/aRylLtawFSWf79yRkia
oMHWPdX3MoKIQ/tvmc9E6szcrlGBp80P7HbImKx6RcHbbBdvFJxZPulJR/PJ4nZxS7F31ge9AC4h
32X+sEjV9ayTkGy9C9SVhRvSxWBzyvVUPdUQLkE2mC7lUqLKMTQbNeszEk1ggX5SmicSmenQh0zx
XfRazuK0gUeSKxHVuja2rI9rpRNWiWkiBHN5RaEtxNiQUuY8tXZN4nD57zX2ZcukjQa0Cko0VoMN
lhwoY1irY7gn6c4dFp5VPNTDPXECzLDLU/n+JW9hZ7UljLMnToUFG5kDJwhrYmHbQP4mPsNE86wX
EpweQ/CeEprKI9Xvfo26pCnmsdC01BBXduk2W4qeVcz1nK48HUAFlJ6cshpHYAd6ehXbR9ZZs8cM
zsVBh6tHzn9HcEiVs6R65jAYEgfDXPFmm0U5B1b0NloS1EGPX1BM4U6fabinbfz0CX/hyStWJTaz
oFyfmCBEyDvXIDIDVWafNSC8hMHoyZ09qu8slCD5oHo93GuiorP49cD1vkByHvnLoimegTebvIe+
Rii0RulxJ4bThYRJ81mxaCJl0+ly9ZahKuG1lMvr2ShTQLE93SffOM9DhuvMrFkXAa5NpkEKLdh6
QtshR9TB5MZqbfngUliT9XmsHDz9AvERzarGkmD4Jp4LeJC/WV50il9rLvaB9K0UDl07+dcEOu2K
eaz+N89OemUEMbnSVWXMYjGQTXE4Tu8aFoX2CaJMlIZBDca572u2648q4n9ZUCFVtMqBhh6WmH7J
2uDdB7uKmYIqlVKyNjqhWGDFQZDAwgHRyXCtSkEML1ZkHVDs+MtL8CE8meJ0qvibjeLY5LBzxTfg
1MO4dyYkVy6mgdDO/Lg30xAozbk/UH0UDhjIRKmXXHI/24dy+EhlPTDmDr0NoznzIPsNPcNVQobP
2Sr9rSNj3HycPncSGq+PwDFbkp1HDYb5ei1+NIH/3+NKXgvvfgeU2fUCZrZVMe0h4UpJdEWBbsEM
1f+A6Ts4Mg3x2DsXkVfpCZivJU0/GJ17iNMssQrtzy2qqBhJ1iJKono5xm9NzbP0ElqgdwJYN8oZ
n32IW3aFtpEafInWNMMMKqEwjAubJsGy8Z+6ijjh5RLF9q8BxxSIzmGTNLz8UY+enSc+dcHfd0dO
qOwgs7jbE/st7fuP5fuhnvwEMS5vlODZv7MVMDXoFBv+2FTv/XhpuaLbuUEI/lQv+xkaiNjn6kgN
aTrFF6K9hRO00KN7O5JYHnugsAbG3ekD+lCfUn2LUpPytywzOkPY7qA36tnZNF1Smkz4VKWWwOCC
VRv1Yq02OfF/bvd2I3w5V4JzNZjkzajKBSxhgqDJzOWYRGLMEsK8PK5GQz/48lGp78kfbElrcO+z
CDgH1GshnUpzh527m+RC5YV+ZSQ2hhlARyEiBbmVaii0XYQoYzflWLn7i8m3w3/rM70UjmbSijvg
MwFtEzV6AkMKR8f5UGa5uJkRAZXIy2v3N+NcZ2aB4udChtqpSJXwMdD9I2JUyIenASYvOP+O/2bQ
A6K4agrzsMrSbQ42T0+22qkPImnhjzQhmNH/Sh04yORWZdEbZQzjIJDXyCJjB6QtcVis1+JF57Lk
/CVOO5mUrYKF46+OpiQM6TMSIBK7U39V+mHSsC4pEmEHAPZ9xgQ/n3/ybAT+jI0EPYC/RqvdXQe7
ic8py2bnXgIyehUs0vQIRFf4b9AAOMGHuTSQvj2/em/WqTZor0sd7XL4Jm7uHF3Tao5+Sy6ZS2RB
XYArAt/Le4WDnRBAp1vOsGDmZIOqRWO11iWzocE7eMK0NqTBsgN8gmByN8qnT6k+TYdsUwrtUbxz
UHw3r+j4ggns4K+wdPwV9Pxe/8/zy+VLFvu/J2YNMDa1LHIihNWPbAMcxEKIvAmKNuVApMxEEZVC
0wh/21vx/6eGw2Uqfm+CLDrBS+a7vw7Z7ai6Kdgoy4s9J4iccukzVgCUIlpyi+eJ+HMBsS9U4KT7
SA1Wjj7zrOlUFgB6a7jU6XQjnWT34nL6Bwl5GhMQaRv9TBX5v3xNGynJnYXVYjA3OsmvFOUe9ZMp
HwswATNDV8ysm/Ukkzc7pGbxsBqVeEsrFnH4QVABBJ0jBpLR94yxzJI8jqdZNJ8mVe3o9+6yNyaS
r+yj8tgn/1oVpsZBZ820zxYPhfxjsUPg9iLWCnxPOhqL4EMLFcRMFQhzNkBZrEvZ261jMlmjRO6R
WqmNwZTgFlDS5gPytK0qnWCON6UaR+iyav8dv+jCLaAAjthO9F+3CrJgIL7oGXPYsH4ASayOrQ25
JyGbCRz0pYoPVUVclUVcbFrlSf5Luww2RN8WUGn03sCrcKVERApHzV8ZchxKuEaUAtT8oU20ngZH
dXtYrfZOSAWOii0qTJmi0dowlhZJzSBR/DtoysTvXyNb3+giQcxuDuMK6G0h4gl+xKNE4QEmW2Cj
Xhj063LQcnltvrlaIgzhegKmrn2R1JlcgUXI3BOz4czhJ/osz0u3z2te0fObvMIzMGc9WdhVCqBE
8igszgu4MDDp2Gyg7A+fml2N/S8uhVC3FPsD6gbxz30xL7NymIV8RsutFvanYPaYSzazYwKpknzA
U7BBj7wf7AUFqhQklOwucmL3Mg/TeEPmAI1YKp0kePVUAMcEIurZZ/R7vnOX7bP7UudXTn88Z1qI
wUWNd9x2sHt0xLwa7wKECMV2aYF67hLh6sTbp97tI1EO6Iv8R1KdmHMYg5zG/rizoU6U30NsWfWc
ew+PV0Hplc6TwBfVXZNg7c4oloqavM2iZ1euTFB3+6QzbzyuZc3VlGGnPIa9E0fZ6NACX3STdWJF
3A4mRaQt21MyKiLVwQg1VkkQH+DjiIoKkLcqOtaI9ljhYyVPGx3C2uOAUixA+u0JppFzO7x42ymX
XMhb7fOgEnfNG9xEQNCam1twtp1teP8o3/XHZyTNpd50tx/I3Yu6GHv3cz75SCSbGK0S2k222Y1M
wJ4Sz8lrdhG8qVaGx5BKSqaIkf6+fSGIErqq/DGaxptjQ1LdjdsIibToU2hojmYqdgfH0WNM8pt4
WyI4ZUBuXq8eiom+IYCUIuC2qPMaAfVHbOwazaxfhLHAA3lUl+hBRDooxxI6wMZFDnhX1BYaYyrf
oVXd67gnPqKlAoFx/Mp5tJ4sKeguHR3pRHnRq4NgO4KD0UMhk5EaygEuDtWLufPrl6V8ko7iyqao
+l2O8bQHEA9ws5ZWrM80RDFxydNc1QfTPyjAruji3O67x2ua/9+JrXr0Zb2Cz1482cOBQDEd15oQ
YatQ0cQXBirjM+9e+4QfKpnYXE7ZzazLe2kxzFqabVJ90l/rZZpaulabeFFrxG4kvh6OPbjRY/pc
354W5gyqRQWesVzy78MiLBb5E33eSIOcyTI5KI63LdLs1KUA4MmV9esglS4ROMkLUQgK5uE8JaP+
QuVbhFoTr6M7Gt9quE0nYS6bCQMJYvmXyTg4Q6tHeQRSGvY0RSyU8xd3FECDD7P+2L6xLzmCtevq
PB6vsHpDPGD/BWx1uDJr/Tgzp28wfA9gmtKQ++AJM63GVeSwGh4WqkJJxNUX31TEgZzB6u8q6Z+P
n2/qOteBSthY4gdijWPB4MUX2Xb97s9VQc75mdT3ew8cL4rT5u7ErtyW2RAw435R30wY1nbuGdWo
cu/LvVsUKzEwFxU558xfEnmKNLWa2+X3Eoj8WX0GUxKH0osqAIIlit3CTjtBSzsz51tyjQnDwBvd
kBwWh7gaukE2GpBneL+hTI9qSIodV3SDJ10vwxElFuO+OW2lsosBPVZNooUuyyU7WIsCYlvmNtME
1RTfh6IYU6fVDIfkq9lGRTVyEhcYgxANRrrohrbbsmFNtwepB1LJRuMEwZ2SHXqhyNxzBFpRBJIk
lHKx6GPt5hVm+VyyaxKS8y8vG3OxtwhhBWbf7ZfecjGBqELAYqEaYIbEZCzbJk0hbqXRiCh2nFE0
TC4++5kJS4UFBRnHt/Oj+rI/yrNILC8TP9o+aKBxaVvgENRZa/MOltaOIg6awiw+buD2HMbSNCXM
RMv9sS+/KPeirtj4gtKdqjW7Dd2fGz2cNED38Pyvvk8HkIQ+A49aDG2J843WtQGmPTI+8ijF0OwA
XtxYGpEBBBKGwF+I0yRoWcTJG0YCxZhLgE+/CMf4fZQHOZhOpZPnS/cgiryydrqwUlqUGZMF0aHb
jvCZ9v7yI4YJPi/wqZwsv8LYAg2y2rFy8fhvYGgpGTt+eztypLJCBS9lIcKU/uZ6kp6Df4eBONuG
6qemo4weVS+ajvdbAPtbAtg2AWxPIMCcjTQBkuTqQ+CbKQdU8Cp9BZAtIsSZ334o8h8PipdK2Chv
O7avQG+EmlrsMgZ28nnLn93aO1kV1tk5UGxDWSs9QVP/K6NETjqX2gIVrPnVPselRpX7n4xYarRN
xmCuYmPITKnxfLTUZg97lyN30sSUo+1Lbj2UTJEV1/e6xDnWPvZEXp9a2xNgjMfX1JXnxt3Fjnam
lcwMQi9uPUfLTiE4CGAxAoElwJyZJnrFZOa5deW41Pb52eM9ONJc4ayAGUcN+Xb72lzmzkaiXiPr
P70dptYYaDHL0AbJwK048f7HSIxWl+Kdw53NEq3wKyMnoL5p3HBQAQMhCkqhU65lmlXppXpIdt9G
KuvhUE0y/gMPIS8uwva1/rDIElOOnvs9h0GZOsVIRRyr6uqE0qKH/3jKGnWywWRMoYg6w+9bL6F7
Vz/HD+YQ/VTRthYBjjIWYD2jS9mNQi6NuXoFNsAswfh9yndCCHz7Z6Ztg/1qdYPcwNh5CgYkOz7w
uBC4/zoV9PtINxVXdT7axwh+qunURz0WxXEglMJOV9tOrnBUgM9wf6XqWBgdncEMKWHK69XyJsEh
U4qN76Hln4f3VI2d5mKAvOUrTsucGI/vFaECf5/ynGYcI755lfL61vgFuNKO9bQFqXVgG0J/+UDv
hRb7gsJ3jP9NbUb8RBtxHJgQpmsFgZ6zqgblQ3JfIGq005wEanh0Bh/XxH3xKgHX/T3+7+HV+qmW
D1aZwYqIHCjRteZeHQlpT8b9KfoH/k9AGh9K7NTbmlX4qlY7ClEQSIJa1D6YrfUgN9S5g9qzys7m
GK4itoTHjyCEWIgtxU1B3pfkjVXCO7w9iWB1/i3DQEaiWl7+YvQdTeTPgl5Z55QNHZyVEVqDfbry
rbvjQ3iFkIkiibznMJh4UWHkIPZcYGDkoya/ulXtOhSka5OQnsQqjPX4hpo8gOcW4wU8HsB4tCWq
n9I3jRNSZI2kjk+aHRqN7og/pTF+XQNw0aMmreHSkeYPZ56UPDs/rUsNObqv4Phxlxv71HvblInw
hSjiwP4Z5Wfe3+T74j5WrLj2ERpaJ4g7tLGxcsIGnzMES8bsjWE78KxAjvBHvlZpempISBVSBmO9
yuXRfw3u8P0L8kx3y5UjBSyHrHxd6by6PmA5ZFAUcnnEwamgRzpt3m2QWSGLtR5KF6mmJD6u+Cgz
qp5an98wOVUqfT1XjpVOXVvLkXxnNfLMMyZVebtrvQL+0JAipTxAmDfsBqtAnNttXcW1wHv52FLz
xUlN85dqA1ArNQNY/vssc5e46Q2s3xenb8EyTn5q5mH9VNPW/0I+w3dSiggfgMAK6bebSNtGat0i
fA5PXvTfS5tNOj0Fb9LgoJXaocRpMnX2Ck9ovmmZmOodRbZUhrwXFU1rL80YNK15PlVPX9zqEb2o
mJDb2Y8ZC1Ylybib9GZS/B1MeZGjF8G5Zz06xGJpLQNm2l4KoNXsZP1BqSNAqYCnMWhJdj7jnRB9
/GUKldsS3oIIsGyx63IJ9c4YASSa3r595OrrnTyUrUXanzVSDX8Yd+eMqdY9aGawJ0/ouIOxDdJR
sllAgC87ispqBldjAMaO6rM0tlGfsu8Ml095EO3y6h/5XauT7b6AzO1ia07yO06g+l+HNykBpO+t
oyk9tFvQjjn4rrut6Dn9fxtHIJvIh23bL9jJen2auBu9CifdtD/hcFauy/VtpSInZll2rs1oMEaP
+bmkogFdAh2jzHAih7vNMw/tdWPwI0H2z5mrwl08hDEBzKebjnsVgzWyvQM/b/zh5HhCyjsRuxOC
yTJX+ExGHYlFJwMOBPVAt1Hldu4gKSbi9BUnYeemUj360rUjRYaifHi45fV7D38lW1nauEshZ81S
YMqXQx5oz+/znmqeXbhMOPqfCvBWDbcKlSs6+yHsX7BAe8aXiLr6j/2Ax9HDI6/8T8dnJXUGx5fG
8AiRza4L9Mak5o4ZQkfB0Y5bldoV37Iy42Mmwo1nbeiEgWD80h20jyflf2OO1/hqccfBWwqzlQOF
c61C4wbPHMrudZAaMnQBhrFcP9l7OAaDN7W/96C5QJhfG6tfWBVtqmrGGdKnxS9DZxIEWX7/VCyF
Qb2n9D1YO2IU5+wgJ6scemiOTOcjCnyKasUvkNUlNWWOck5Keu3yhrZIMJcUBXHT19UxQr0v9ILX
ASCTcNvyqxD0i3Lnbx/mQLK3LShsolin6bBRMCpILmsSG7cGjZCDKquvlmuHlCUZUh6EA47jXenb
RfITxqXjswY5uGOhQybi0tCi3kiJwpfVU5JdX18BNLMtWQqlbMOBKNCDRiKDyDd5wh8l7AmsKOH+
YbThVAWa1gzI0b3Bk1HQnqeWl1igjektEOL8zuw6ECkpGdlZDsgpZSWGhi2aEXu4C9H/29wBZXwb
t5CHVAu88MdkAtbGPgFfopOrPhIlvOS2tzYQwJrMSqmLFJyxIEBv9Pe3AADKQb9qHNGuzkg2xvfm
8nW/o8WHdPPfcGDqEYbB/IHEZ5hc7sOg0yEISVERaDwYx9vBtjc5QqM2cE90EyRUyv+c/sEABZip
+sw0enKx9eRhgZIN5W1BhBj+jnbd2nNbruHYv6IaImksHSNiCvx0NKriq0Sc9DXa/+Ro7tRqqyPn
mFlBbUmR47ZnyDX5jh+sq6CJ3L1me+yMKm1RVJq9gz43LJTpl1MFZVUZgs02cTqR0aHUBV0bxjJj
o4dIRfgWz1eNMtqmfaattpPrnmCiZtGgYN0XL/47lh/UoRV0wvwwyj+uxpebWRzPvyDVgLgPf4Fz
A1QqNlHOQ0NbPEgoIvRXDSY6fQBaCbsdmMG3uG8YQgqOmUsMRn8hpG30rArp6ngbaeBRoDlGl0Zs
fZsdocbAqhrquBTzbrqtJxPFAPL29SGPlXCkCbN2BuOI1udph2HhOqNU8y0ZBN05400f2M51X+pv
nlNyL8+V5Yl4n1VeYg636oUfoK2q+Nk40w+xtIZW6c4W4JuHAadgr9PL6HEygy1YDu0MKbM9S1If
RahJ8N3al84/xdpbuce4LiB8fUxQs+2pFAWId+in/Z5oLOP7uebDEYCDBnI3eiKCLTwWAhuFX1LP
VlaSR/tYSYZvjDAthzh6tBHoR4QbrS4XNtDZLr2zWZTgIhC7zmi0JWb3IbKwR+d5HblaU1k2sCqe
u17QKSEh8pkyQpJ1Cj/x//s9mrrNeHXRJv1Fxc5gGn8rb0VjqpkdnE8eVKcZyFDDqHMRhKxFKdQw
UkUYg00GHSDW05bjeCsZEEyOdq6wWC9nZdyQa5b8DwjL6OJ4rN27kQtUNFQOPX6XUOQn5i+UemUV
lHOT5DyTfuNtMnSAr/NYTdrynititzTUuj3vi7C7wMhVx7xLSkV7m/3gChYvVYbJoq7tSHHpQi45
+4fc+oxFZOVerTJQCIXa8DvUbmHFGWItWwegDxYOiE1a1NF0KypR8bdgLP6Q86sJMW048Oq1k0RO
LR4l8mWphcIKCQcUduILa1SYZqEkxEkKUdA/V23qpnmWUuGJlS2e7/aHKid1XeiVCouxddjHLJz/
Tl82ORz5lalpbggE6jNi4ZqCiXF78+PokqfjKV478bgb6o+cHOX+Yv3/bmfOSfJYmRmf5Vhye5Z4
Vbv4lYap2Ncs4h6902pnTx/xdukfZRoaIqGauRZ5ihMSZ8Yy4e51gOmODuqAbsi0+PVK6DPMzwmX
Xw36F2kA7y8XS+xywRVbO/eZyIiY050/pEQvAk4YagBFTtc7J2npcbQesXZWks8vJEVaJHxFz3jf
HKM4lhCoV8191zvqW7TXWmqaABBOmZd8TdI7vJZFNz23aV+orprNj0libE4MZFqyz2vrr8GZkQ36
zM+IwGMJ/5R7kBJRBkVqChuxbIkrRGYd2Q9TfgkdEbXQJiPQbjUZrlMAYfW6JKdjDaspuOd4Hms1
msTKT9nn2mn0MdO3siG3UPVuLnhrvHOd1RUN9nfuN/NYrPg+yheisL3G99E4T098DlStlVYd/Zex
BgcWRYNVROgz8XHe5YsqsAtMCtaOchj1rIClGMk9SC0dvjFb//iHContRrewaib5lKErmpupWmw5
OMi2dlres8sqWBCgA8ub10kJSmW0ZaZX1qpFh2Uo+u59HlyEALhjAg/ibvNWPzmP49NmOUN4is8/
aFe/NeZdApeELfopeZXjfb0Wy0VJK+8/AA3uERLITCAF2zz7GGcLLSX+TURKKBnXPNwYx/hqR8hH
X5YZPmlJBCgX0CbSOHOfAd31NRJSbeQ8ES8hq+yfpIjBGe56XojFfT7WFRTrjSyLekM0y/hJSSL1
x/qQBEy/2VPpZP4TynlOh82w10Lo1AI6zFxAOn+GRsAT1VSSFuuS6bSvMWuly82XjGW3etZhlNu5
rrJK6N4P8dVgQAYO53VRAo7338UvXfmtuuJgsnLFZtC0FiY18VoQ5wddCtWG6pAuoxh74lOV2EIw
F4t/yx02WtRpdbhuSU9cTJeNPyq7vSllIj3M+/vV2ZRHTV0uU2u2g/s0xJtrhVXWUt2lSbW0r7U5
m9E/XYe6Nh+1De2IwZo8lBHbHQRj+h/KCsbgbiChVVsBHeNWFcrr/fp7GTRgSM/cSlkrgZFPDL2W
bSekBBpOHW0Hna2yenhXEwQhyX4KbBC2T8yMAQYYpy3j7i/qBxxlZGh+Y5nlHs3zi97H0kS5m9Op
4Dy+tkvIcmS+46GN+C+xG1B0UKq/epEXMGaUMSY3ZDStPWGzYKZAXROw8Ki7wTEjbUp8YGHpbibF
7XKY82zVDH6pIvGRpbChGtJPC1RqyK0fJ1FhBNdgrJs1BkjgDwufAfcsZfahV69h2oe0Ob4A+gMb
VZaacmZp3lLK7P9askNtyJHbqMmT6N5Fx8X986FTcEnoOjC3DK9Hyn8gRv/2RgtoZJf5iMKSI+Py
6NGc3dBps+gl1d8yfJmbqL1uTzpdNc9AYRDCJ/mNZt6+CTsJfttUjrGlfo8aEpYXIfptAGuapI9W
Ix18F71+q7o6R6IVgFpD30Dt08X/Fmi+1yThS/jJmnn9Im0bkO+pELSw9gdSBnJiiy8eyKaglf/P
p1uzTnHzgebvJGGLF1j/J7ZMvmK544sE287i9LyICfRu+Zmhu0X/2Q5UIVEaieu0+wj6at6tTpKr
CaRI2Tc2hXsIFYZyNtr2Xqvf0KptDx5w0N576pmwSXOj+kKgdBylCbY1n9Lk08y+exzjlwIO6pxC
z5th9bRpiplVdImDH1W0YX7QHkzd6n3TK+J/gg/ec8BUwtFIb7NjTeLeNArY2b5/Q1JgKYUB6fSQ
IXrXWcvfwkJnLxrra4D2GmgNZzly+dUFvizSs9RZxwLTqH52G5JcBN4wrncuEeSUtHEHsnm1L7f9
or6Lwbcir9JwIOKN8a45zZtEUCIfsd9+8LUf5ky4eDbjClNepjTgw46G/d0kuBqjwIZYe9BDaZDl
c7JNrCeFpRjEc8k93Pm9QzNfGAgkbvzgM/4Pn3OztUgk9FuXh+RF7Ymfs0FZSZjq/WTQ/k9Tio52
UUQ3J+B2yPs2JlWKajwb3i+yBLEATsFmn5bMVGtUgtng/0sErW39ddgJofIQe1bhnejyCu+evoyj
R5/GppQ/5WWb/11xmtAKcZICWMRaGJ5ncJGETc4WvX6sX4cWYYGn/1zkXGaJmWCzFgkARh3Ax/Uk
gGKY05msK3Z2CRKMP4mezIU+6gcgh+AdJnoAtJVZCADQzQNAd7WPK0nIpGXEmO+aZtZEQ/q3Bo9j
nPQ11LCPR5QOaGp6IPbWU+kErwSEIsKgtQ2mMjGztgtcnf3AE9peYmvn7u5DgASN9dQPFz78nosg
NhN/TNufQjB80gueVGEL02DUkh/sMXxz5KXtPPpbFYmDMHZaK3gM2zt4pwdA1D+81M2UOrVsaXn9
wD9xbrm5Cw+g9hAaThbSNzcB/zOXf+lqd8e5AIwQxhHo/4CTnE/yYyTXuL/bhGf4J8wZ40JIJsI7
4zmWY31VMuoEQIFIa/2NoBaW1Kv3hvr8m4N5JLIrSiXdpQ7WJYI/AbVjHbgaIqS56vJ/YKMBwl02
dGdDm+3WUOnMWFlOahDy/aP+S/VgTMlaOCuMiUNGBJg79ofMUPWy8YqnTHYC9IK5toMJ+bnfOmCy
aVZRymC4jqbuubVtQd6A5NNkqYjnnTgVs9oH+oqzKSlj+L64O00yAU3sZe/yQoWp14JplWSoI2R7
vJioThD3hpHclQCHHcqSLNRf14c5EOuQj+xP9WPmuyncmDb6liz3ARu5MMR80UYcK4mHqiidaVaw
1+Vq9ib6uRyV/4BFRs3HSQbIFuAs7PoEHsU1stAaBiaXvKXYtTvzDN6j5wYPQ5EWqKgs/i6TJrYz
BI4GJSzKQxjSxWPor5n3WT+hWnsMMGuBUiiJI89aVKZKDgHhsie9MAKAfET2TappIcac4Hil0plX
UbbkS/o5dLH4qQJpGoT9e+L6Z0XnOWsXrcy1/rWQgdah9CSfrZDTDpRekzq/g8WFgtAQJJ+PS5Ha
2b0MC3WMJgbaA0zzR5dp0JplQr+/x2pdGX08o/D5Nfbzgmp2WHyWFPsUP4jbqpah89ecPV1UFmWZ
eOVR3jd+1Mmn39bDRbSLUADLQMm+V99JQ74hHdxc0B9xXZlseKeKtbrWM/L6iC33qemjsfC0MKNc
MzKV31+Wrz39+2mGWXnuzh+2n6ruG+QpynGGmlr47P14wHOhi+yyNDrcgTEi3FuUsJd4SkU2jfuw
WphPts7gt2bfxtMGLiHMPKH0ewq12c97850g6ujQhrn+wdGP26bg06V8RbA5q+DZBvCyg3kOe3BP
52hlx4xxbApe4lNc6xVmZr4/RUxuOtjaCFNyLEyhpFaVtT8XnO4i+QcBKaARj5nfMuhNkGBPsCZ9
tcQAGl4LDm8IWcovVq/CMfp+6kZdVAKeZLbIv+L7ZLYuLGPvAmjRsoR74jV6vUqIvg3mCuNJALP/
RWsNahqtc/Q7W964loJslr+Q8LawliKonuXbRVa4NqwwcvQAOG+GlKcynnHy7dDg21TuUE/ye1fb
lmzAZD8dr9DiZ/5rqkSIDCfyOvobG3t3np8mFXgVZs56lVhUpWnjkR8j5XP96wauqYvNveJECpRo
nUt0bxGCEcMm0/HgEX81FmGMhB53HxQP8huvjSzQucObXDAhjDIM0uEpxcdZSlkxlysjgN//0jCl
jxZWcuENxLQhNNdj9+txQghecgjAGdH3AmALXvghja6r046hrqs69kmUt/m2WYDplNZCpQPRWtEV
X4ZZ86PY+kdy2UnLVEw8LPkuZw3HPfsIEfPmr/RKup4jrgnbCvvJs1vGBO8VK1nS+q+J3efhFyP2
B5mTJ3b3TlBD6ShfI7XBNPgLe6kulr+NCTix5NTUR53qkEOdj6SkBmHxackoP5d208C6B+sgbHf/
lLPcSOqoYSPXGWPpRjQGl3k8nZ2jKkzGI9GtR8lNfpyxNtnDREQrH+WVbMxQgmuSBuNHPC0c3d5u
+WCAB1zqAukVaNAWT7kCPorGyKdUhdOVDIrYp39b5mwP+XcvvN+peZ2I9+NdwHWQq4i6+QwmS8vk
gQ+Vg6Oo1AnOTiy69eP6Xxv1hRX+FZjvxnrZrtNHyzKu+YjomTsTkw+0cG6l0L7WDEN31fCmMxPD
t/C/rInxuN1CeDsCfSLcOjy5stHsPHt5t+uVA16kbvZ5c0iuOFo7iEpwaV0wuFFoEcJLeVxzqnUn
tde7bTEgckt9RAg+hQfrsBOROdK7fFzlYBfDj+Ux5FpBqZpyLIRnCFOeI953VX57XVoa4u2KyGcQ
nyYlIsAFwmvQFw+33W4dpfglzIhrSpJlHvuFd5okHaJI6FEwsk3aPkIVs0B5cn6XS2f4SDPGT8WE
YJbN6IE57OZ3kcwNlLwZv8zfADLOh4Qw1/9BotDQOiOU5/Kp+lJwALgTXT5Ue446SpfG2+zoqXBz
Ux8uPfhHI43j59yFbSniwKA2q3Lb7T+g65lyA45YbQ38t7C442wfQTTCen6WWMEF3dPDL/unbmUy
SnYWVgpyWq3dhvqHiCuRer5iyGtE3Mdaw8k9QvfkgP6hx8gXfjSBPCIxKp0fkrL4Oh8XqVpbMuY2
awpDq9BQ+VXremiyl2MQ20dhS23b1LB2aIlP51QtqGzUJxpxRqv/dtVWXfTygBj3BUEv+byk38ss
MNneHUHRhrrRTh+3rn3ZGa542adGpZla725gpwMkDqIvZzr6IjAZrnis+OL0jqY9RgRKBltx+ryM
dH3fL6m/yZso99+spigYF3PeALcv1zh3YseeP4nehPedF59dyrqNQdxeezLPo7l+RtT0VJuvm8Y1
AU62ZzzaxaEvjdKxKI8z825xBdpGqvkTy+7Zj1oxK8D6c2vL7HeE+ZjIeuNv/Wcq0diRTzUTtzq8
bvqqevMRsLVOJpn+h/jN30R7reKQliisxIYy00gQTbSJjh9usJyy92dwVMx9r2EyKzrbXC/x4epd
wjX8WUc0uu31T/jdoqrFB8Rq6kAbflUE5LsFRoLgQampNUb03tpSg7mu9gNBlu7R9cs8q2dKwHqX
tTyuA8K2CDITJ0Vdcv8VjVcVJPUvhqAVMOger94cxh5HnwKKO/g4nXW7HooFvUaOFzaX3XQz8SNS
ce7i1gPydXbJTgcbhahIkGgZQtMSAHkd8aZbJIn6h6cvlaN/kt+bFsy2/o2hcsOqx++e9+7YYzKf
CgUCbU6914GnVWRBTUKJyTIIHBEHTokE8FRbjeqqxnGVrEXt6A0ivwiErm8+7gJL3fKUsu+GP0p7
M3uaFCYAlNV8duQNTj9TIgUWMR3zdq7I+xDbpuBTnMGGbFmiiXJ3yanshU8zZaiO/jNX7bAFPK1V
O3cesGBUe00HOQ83uss/mgJ7q9NhDdE7rD0WSQKrfu/1/bWv7FmNL6YzAW11/OsWzh50oYkeOjXr
aIjKWWBbNy2l2J9qRAZe5ao+Iyi+/COsuLG39HTa4C6pxUVQpXLMXKEPQOkPSW/Fi+J871VGtZk2
nVxjIVPN4OvFXLjFFpO4eercwWnDeJRMHCOXE2b0E+iJFQ+eQzh8lPVeuNsuYIA6X5CGZNXNucQw
fH0rncA9BtuJa/anNpJIMngAj2pMES/zrbJiMGrmDAQBXu5lDqEBd8Czy/bzROzztC8qosB9/STR
p1sZ8RT+gieNIuTQANuXV3RmWOaQW6IECjvbK9O70DP4n44PZGtdxHJkrm1putLk9tNZMzDjtWi8
kSxpef7RjJID/Xrx1OahIoiD2RalgqUpxgqAP64KRhfzTpEKx1SineclZ2P6shmCu5X4yDwc4WyX
Di4aWmBL18xKoyPReIbpRSTZz3tAAS6VPBOBiXhs+t4R+JDZsEBZ/UBB2Lds+X4MdeExq/pv+Fif
rsh4PVvkWTwbelvyLjTLAf3DQsewL7msrM9pWse8zVrGQocE/fdXPfTCDNJWClf8gbDF6lvnEJrS
1yHl++bgI0CK0tx7mgGX1msyGOwLr/qbfBwloo19HscH4RfqG64ax928DXmb24mZQOC3lUtP5kNC
4IAgnBHNC/OV4YAK9zm78FWvqQxIDpnJGc6o+9a1oJxoexLCO2toYwFXeHqu88x01fHULXYNLeUR
uRVGRMmxhpLjiAynFCzRejykoGlD+7avJlqaU+FNhdtgeUVQYMspVddxdhYMEmj03L8cm4LFErvu
StuikHybRFQPMHM2xXXPmKRaDsk7vqcVJGXp+OFsZk3AGqtKh0JGyScHZAz/my2k6s2LO2soO7H0
qza9VTvyQ3vJFzICbgtr1svD7LXzBWZ4wGSS/oxbzWtc6PV1gbi5y1XHFykg76iPzP3g+d1y6K4g
tJo1LXbNQn1dcO3M1r6mq20mdEPaADzDoCSjNN+4JyigNXZqsvpQWWu5vKQVvpkBIu00xazqN1wo
TDBk04Mi5H6MPgdle3D/0UzBDIkVbhZTrzgva+eKTgGjNjucYBnGv1tgZpguC/TJS4LEvln1i+2n
9tszCrMNLYeLnp8+aIGYT6aQStDz55zJvoQXZrIWxsOxsxJTsXmVtJGRKiCW/UOM5SNsa6yaWkFL
R74sMoHk2rVlJP2gR1mQkA2EWkaZ+mQb61glUZsBZy/NStTEBevDedHCAcfJortb3lLl8FY4XwWl
PxTGq+tU8LqKogn61Y6Ide3nmfdE2k/nJ4CyBinmFkYoWLjeyPc2E6Y2ZOoEpjP6xpeK6iup3UoW
wJRT32fbUOMMmq40MOEZnoyOiENwz1UWUBK36KWmFKEuqN9DZ0O33lES5aEAKk54i7ljzw/WgWuY
5/E9lU4piWTw54w5PWaEKfOrf6rEwhj8az/Pc7aBaM+czC+J3/g3qu6D9kElEBsaVFfFXg7rZTa+
qAUb5i7XxfZP2TTP7KffmN7SjpwVqIG2hMTRzrL8Crh6W0pX91cL6D+0FT1fPCxzzsxGbH/i5K2P
HbdB/wXm0xP0oQSmG0PayCk0EqAR/2uUGEYbW1JvI4SMed9OL7OAwNMCM+Qm8vlvaQhWXp4fmD/7
7SX8I8/KBzQxXrR2y/BsdIjR2r271GOeg05JIUhEzsIUD8y9xSqQuA800fNURgVfuvohOpxNjgA8
n3JCctuDx/PpJZ0B8CCb/9dDQ42lInkox1+rFvVSX7inwrs0c9Bmw88SktML01CcDFAzVOdELseY
owsHEJiC8VUcUjg4BF0AInBrEVAoqlnqE3z0JK8Akj49I+p3Ub7lWSfxrJ2vAupx6MDQlPaJM1P9
wCoyNHKGNqeE4a37CqxFF34ll1QdIt3rfL7zAq1AAtTMuINsrmiyTMP/EuUhLO1rArCDqjSGJ17q
twngNjPI/KQ80/MGMoQQ44DKTUwAUVRvS436DwX8I7iGkOGllDnnLwDqOPt+5KDD7bPZRMLADzUt
/Po+Xiw/+nlzJs76ogPV/a35lyRZIyAuLOc4cX+xo0rsRt09x8BO3xU/z73hhGjFfndpiqgCP3iO
fQb6OnBsOD+TJVmUkIFCp8KeRzTPlApUVB+bkXzDxTZyhv4Q/cvzf8w+1zH7z9Ds7BjtmJMES+m7
Xt87AkaqKqCQTnDmWfQBNWOcG/fzGy0FYNPymaw/5lwD8TYwikkfb8bxNnk+5JgaBtibS8RMGbvx
itH4Co/+wkbJG7CyjAy729XdROSs3aXkkLGtm5sKcnqx+fhOQoZarTKmjSkROwuEc0IF6X6q4Iec
3bmvGe0UgIT5ndqKbT5a4Zc/hQwniIU4jtnCKNChxO3arrRIgcWsD1tyiHTz3iL6NvOHqPU0jH8g
8rXe9wEtJiPrGTBg4OOzksbpv+nW+RISKRBUkRpPWH8g/Q+1Pl8m2lXqxSXLEMjazakomIfLOq8e
/sBH/c9uBWV5s6WdycXuidnyu2099lLTYWCiwEDriCoXkEI69uMMQoBPqdWparMF3X7n6Jiz/rqp
vL7vxg70f1YV/axm2ATXPPv3Qd+ZHbzjkx8nGB56F/ZaGsx0p/Pl8PuOxryAJhxnwWwx2L346ARo
Abf4X8TyILTojTbiIlsRplswxFRjY9s5pptWZGU0PFZJ2ZgCZGFNBuVfz7Sh/iIhjvRV2KOWxxXx
umfTx9Su2WadaczsHWizSKetfwkrNft/4TClXpbbBPZFCB/jdonjEH2wDHxD15S9qtaiLOYBxs6D
FsgxgGAD5m7sWCoIGzfLYl+/+NFX9SkNNZ9PBx79xBMTC99Le1jqI+CLTLC0kHjWbTY0PlQcM3ot
JVOL9Cub/HdghY3ZoRBj+x6wwsyoJ+Fz0ks0YXb0eCb3/YHsbtZRxNbLDzOc8LPPix9tjc6VMhhT
UiuJ2GahPX/0xzoUlRqi6PEAYbl8jPXBktvLSyz8VeE4EO6N5K8hVg28L3tJlSsz+8R8nEfQut0C
KgieAbc4ax5dWaPQdB02MKvwn8bxjh26oOFlW+v3DExOsvkTPfnOrYTHtd7EE9xLHOuCrV7tioof
HGsh82j0tHLch/YnEDohRP5V8xM3Vz8dVGT9c0dta7Hnj02hTLEPEQUulCqtk6nhZevD4JsqgF7S
PiMT/c1VF71O3zkJC198yfDKArzcbAwPO6Gz9g4BCsWvHKqdlagMQzBhj+mHajBDIQSMy/4C6+p7
TCCxJgOgmoa5s2xLHIUYXkXjMWDRduAi/VFmLnnEryTZ4oHl+1aYpmg7vFy9Zs7CmlgBXHtRtV5q
Cu74+sYPhfYvzCV9Vlv5QwReq8+zuu2jA4JF2TgTPsTh5rbwM/UFClMpYwsoSIgWvQ84GHO8N/WB
WhfvrSfI9p/STwwgLj6qgph8hKH52iSX9PqVNrYWzl5HZzTd3eq82K35FYsoTAYVnEZyXteGPZfQ
0NAEVgQcKWREkw6GoFDrszVLrPd2N1HMvRcNqxvt1kSyQO02kcArgYXdGRElRuN+hQ3UL2XoY2Sp
2Bee8Zjv1iw0OOyusaqLqqvCmPbzVLHhyNyaCY8ZhzegZBSD67zFin5W/Xg2sv9QH2czHAazk7gg
5usIYaJIHHo8isNLJzncowg5y/gXo1cA17iIEbQci8R18kHu7gNPZ/gHjY+3sBe7dJOs7nc3CUwl
kv785qO9vh1AtF3cNbb7TUgZ1GppJVYXZby5yPxdAQKc6dFc8tHgpLnfXTcbIpnu2TaJEnoOrIkS
lOiNfiF0kqChg0pPU5j96EioQIcfVZm+MVpe2/4y2jQ7bzlcxoHJ5r2gzT4FhFbTw0d6URh++3Cs
sWvSq7n5PG6xrr+prAxLhEchzeewXXwtwtrVuYbsxE7EWFiZSxGqioXX8t762hfi3dRYNRL1lIYf
gqbUtPWXvRMPuKDnd73nbNJCbmLJL3+MizV+aE6c38+P9aNsF6Og4MRXNeTPle1rJPWg3UX9O9hF
AQlKagchlHaPy1Eov+eBXoVIoxkbFa42dDxqX3GsateGrbIviBdxz4YK/5ea1HfIto+Qyg4Q20+r
5Rd2ZVVjsaI71J4amkqmouZa33BsZQJiXp2nGZXYoBBvJi87BRCynso2GzXFYB4r6JryN4hPOpAN
TUpk7zVC2SaZrq4bG13zIwIKiK9p0HGQ6X4I5im0IsC1OBbA2tWcdMRMn3HN+579ftSa6Lbts6t3
FoWyAlmh841XymfJFT67tuhA4GSdZk6q54/qR19JB4Dz/+DLqMJYc350lZ5Ti5vPJI49/1wK1LRI
9XdL5zswyMgzSOpZstiL2ZMvr4yVaXt6xM1kdy0162l2hS81MAU8GwJxfkRBEUsqKrDJ+e9ERN5v
0IiFXT3gBvBE/UTWr0mpF21kxc/Cv0rjOb+9og7n7w2le4WFSvsrceenrIAsyRREBOXBSRaiAaGM
dI8DIedPz+LW6xw961LNSgeiSKNM7oVOBkfM8/CgiYXwPh50YKw1HM1Tn7F8FBlGeG8CEGAkg38R
Nph/obU/1zSuZZdAtNAGm4y12r6Ei/YjdpYvewiOM+Znxbw6HYLmKv9zUgPaRV1dXiZk5CvpgnU7
hMIXjMyhE5mQ9/6q0DxVJTNSY0C7afEXngDGm63s1qtwOmVVfJXhUmiHGbfqDDMvvLmhwQXNaZKg
lkXNaVlCyqKcWCNNdN+Q0ReI3AEa8UanWWNRiJdVhP8i2sTvHBWp1X9ompbMd2wcO1eeiy3+2Irn
sPezsG0YTMTxXQu2iIpxARx47lrcSCq6+K+1He5ASWk98FCRGmVxWiQFJyDPRqpsqNlvx3xgN5+b
sov27VysO7k4Yti3STmyff4XiJsQL6mM6Z5ALFIkIR0TcGm118W0zwIoEWeTdoIVM/QJz8nzcsS8
+feZCJVhxvzDqn9KCujzV/NOL+tvL/PbXmEFrhQ8ApfErZi+zygUmrX9dRD32s1z/EroTOq3ScUL
7U2lVPIEJQamYVZxdMEWLHk2tFTPYRsDlEoNpKZ8vMirfnqmcnHApxgWq1zz09gx8auWQG8ixRAX
f2GfAND/nGragogOJRFg+pzBnmz9U/uekuRBOVTa3IJcsHnDnGNU+QIUvgnc1kymAIAvj3ChDFkF
hzkbwtI4u16WzPZKOjgaJZAselSH08foO7XELjd0gKOKiadvZxnOjvR1EohQGxJI/pfLzq6yrMpw
xpuO/7NH+0/kMcYqa0VJUNwHCzIdqFv/8QX79u3wzG8O5y17a0YeMPAeXsqL0kdTgw0Fjwfcc1yy
98fNUfDlQdPganKWlg6L/P/F4Zcuy16JP2QaIZz90fFFHqLKi3gne2l6zdh3rWRnCkdXaBMhklSX
r3ZaaRLFCCJVDbCDJ73ZiDF0bHUwq5ssaaaUXLFkBeuso6LJBzaFYql7JEGkqR0ZBh4MRnFz5NqU
I0VlyhRVKH7331R9n4WILDyZr69Pt7BqT8EzTr0B6FgKg+b4P+wOzLgjOetRO9bvk+9OoPCq/KVK
vOWhxiNz9fo5I9I3+oDbng/g+oBv9eumj0IbXmDXeRlfDdcNlBxhgFKshiHbmUOUIIcd8Ac3q7ti
ijciLgnfef29JWm3SUAymSQJZc6AXN22vADnWXnw/CuVDXUNjDwa3ILzoUIF3LnuybD2A6z8Q8ms
2UygMCx9LQSm9xLXUvaZBNhES6DtqRQqlQaffexfD016Ve1/53NpdJi6pN0WADY2B1Mo/bYLIehL
VzYfDfBWn792YHEU4OMw64j9G7i5pChF4EcUMD0TzfoFW6QJySJAWsYTQumTGz2rZfOvMIfhp71E
ZdEafG9mLTs6wT5TVonWX2OFGBTAvHOAJvxCC07epL/Cylkw12qchCgJLpLb4pKoi8aGyVRApmTy
T0QGJhhvE2TNSWpctVd3oN0SnxmgSzfe60Kl9MyFylCuVhop7MMTDipwa6sAseqS/6qPf87gs3yZ
ly1RjRn9IwQqncHbRODI8ggaqsP9PNTyYzKaxdti/0Tv3M1h+Y1lQYNsY8CYlItAGdteX/uoBpaU
+zIIvm7AH3W1Wkp2b/IBSNqCK8AtW+YYofCAq3JhVkj9CVtPzdAzYWxTCPsnynnrKQ6bLe71giDI
9aHhzxnIYoqSUoruGMh+hb7UDan1wm8W5n2ETw1YmYMRtOBIV4luEin59SOZZLVyZoSCFPHImJdI
M429ts+YDdO6JQ6m0Fe4UF117nFdSiTk63vtyxqRNGAwAkh4vr2iBOw0/9m5yJ2CSRYevVmdodLA
vl4jVLRXMyTJTscEn3xBIKUXz7zvNsdcVTUghbxaNsamQ9UFcSbhnKxYILG7gpZzpYo0cFmGKIz2
f90BUznz7ilU+MGMLghQJ6eJ57JGXDf1dIzK1puouxzDZJvWOFOTRtOj6IfLZdYrCKgJoh/J7uPd
S3F8zt77FuW5WgUlV92L57kMdLZHmarrKs4h1rslukhJUm7K5UektJcQG2ikUDdSvjxVaNIHwa3p
t+431RkIibewMwZ6mI1EtlURCpYG01o5gXrbo5BoJ965TvpngroRgK5BqYrv04m6c897x97DUyOS
CM3Oye4YO+HNcCPmL44ShhbgOdakpwAXYEy3oSmWtIhMWSaZLcufsLRUMDKR5tgbsQ5IEzo9D+Wp
jc/33NsPwzYvl0tUkYnvchLaTdK0B1rNO/RtzfVm7xpn+M3Za+Xfi0D8LYwwEkJNBQIyuBwyfpM9
cKnHAm6apdAks9tw8iVUPcDlzJbRz5SAT2JV4/oxvO+nddCEoElJuNHiuwpEHKNV8+uSsuIytyN9
kvDJ2J2kjrMRyUNNxVPrifzO/eqo40RFUUhaot7AibcFH5StO8Qh7Y1Fsz6E0KxygDLIr4NRk6p/
L4wjllhcJ+/Z0288DRfbD+WvR80UVfQuzAEgO3BXUdSnLz342xQMXWkQUopWFgDunCRyUrJeqmNZ
32uvvhv57UqBq21rCyimvBtm+X+gUjnRFO4eenSiCkrxxFpXgoJVqO2HMyDxCWREaqJym6UVLs5Q
DeKjFmKoJhYAweqyVQZS/b2ncpKdfosV77VWavC9Tvwk0QxV+UxhGCbiliwWK1pa/z2ztyflE3IH
r5RXSnF0CU+EXkvdcp9LJv4qhaIemR+5JTBrlub6aCpyYtcZeYXWgdIUp2OgZ5eiyPuLLkwnSROm
mU/Dhz9FpmnYYQ5h8ZKBnFbU/hdXpdaNdv7gqEDG87eMS9aK1bqzF6dcTYxKTOV3PmTcdyc6iaz0
yYCmql8NainJ2CCylNC2Y9eBqEsfM+c2CI9rUMv04X8q141y20fpyGlBUXYiE9StYT4Nylx81v59
NeDCuifiwWbNs7GrIEGySkSlTVfazBM22Dpxq41Fta7Qou14ihGFvSQ1vRja45IDx4VxjWZL7PMl
elFkT8nZ6tEUH+gWL8WAfU7KgrE6ZDzezAaxTFB3Ce3gb/sq5GJ/2VAdCuQMyIUtQr/Mc+mQDXvX
4ubdqTnCnPs0A/lxUEFrbEf0KauFmDzLwK3CtN56w8pBp5S4cz3USBrZbCu1Zuo+/zYKGKhmaIZr
89Nkp3Gm0/wxKV7YxwWVz1GPtcZUE3hmswdXz61iLTo0nw63XmGweLdoa9ZnSln2PBscjcb1cTSC
B30XB0lw/p7/RPiMjvtapaxyDp5TAjPDwHkQL39Md6SMmqPj0xhybv1pnR3ebR1b8Y2u7U/wFdcK
shmj4n3ACNDNvOY1/CCotGOlAs71LwF28Q3CB/uO5TUUPS4X/PK7hT5Lm2A24za1YLa4OWHzvigV
MB5P5FlhijWKbSrjkNEVhpW04FEf6VEBQSVjc8rZeVsL1QMtsZtENhvS8eqrSvR2TYM4LpGwY4ml
wdI+xAcM/rsm6Q1knpaCPgXX5vXHWq8RK/uaxvXRt6UEzm5fuhBCdO6o8G9ldWe5VmvI5d4LOnBG
nvmxS0FtV2LLKvdMfdxraEof0E6goqLFYs/4nBK5TJomSRkbZ/1VvfXWGrgNb/Y2Zj2Gr8ylj8Uf
mHJlnlydkbPSEt8V33Hc6fZ91BkJFH0+6qa1ejv9j/dDbWGptR+PheHGFH1eG6l+snBiEdRjjR1G
mtemMzCdG/c4s6dV3Vh6rEjFdge1o5sOqyIcql8ULkB9D8wH8mRADp9uWmfvOjZVaoifMt7oXcyb
vpVpn8RxoF8QwNA2cs9S9PdYnKcyFD32CcqKxWKevRv35WDz4+y4+x4wyLeApgpIBLsKQR69TwKi
04cCecr3vTw2YlUA/yqpeB6C0re2td8yIdUEi7jSaLT0UIBVRJaT2ZUqrjD6R9RCArbqhJuc8dXU
Npia+ZddOyFUSI9+IQl2StrcIOZB+YrCQYRbBhRYEwahRrRtamCgEyJ++lcKPweMtuAEwBI2Yt0C
60CzA2bZJfiayK6UpncEBSOw3noNylX9Eh9OAH3GYYXdwc6fhqrme39Ju8i5dn/lUtU7hLAZ67wk
XSB1RTqToGgkJZektDuasIMRSU5YMcWUxC8HaoPjpmWPrlQeIT0yYZaaIYYysjR1ToXwklkxJnbA
vtdPW+dTvKhpk2Y05KcceopqnpwvdIQwT4aMQakGnqPU21jhlM9K5+roM1CK/2bxkRf0no6rwumA
g60kKH703TDQBi2DBNDyZix3FRox2slVwHrsvbJCJTTaaey0RyQ5tuM/m3yFKFKF3pEJCpjB0hcS
3sc+E0MMl5F2I9OgANyXSHgzTxy68d/NWfs3bKLJc1O/3YpimZQUJKF4GAwzTfSmJ33R7MgfUPvz
Hvwh1PcpTHqcApr8AmvSHZPl/WionDSu1l8Sp/kzTgm7+TkZv74XemSvwGA4CUfl5slHC8rG+Euq
hU5WrpuRySt/M/He3yeGpe+Hg8hx4LYDlSfPtXWF5kmUegksiEGq8Bn3Av1VoR4sp2lTFAB6ojpl
LBSdEmGc/q8xjPJc3NKP9Pxy2Y7vif5hO5tBcCb2cGiGlb+5jX5/V9y/yOdCadRTJN0nud9VjOTt
Rfh8Y9wUCKp48+J2MoKuKt36l5zpox1lJeOv8HnDn027YQs6KgXy3pku/2ndrVUGM9dBWyVliNzk
hzzS4xFOxZ5J3RkZ52DOJaGp6psi2QLIOFXMa9BH6LjmRLTgNuovL4GRVjgjhs15GDDe8j1xXM5a
ZfQuOMtAq3Bev6kdrcXdtO/Rs36YVVND9XJ5WhisXIo8n5zmm9p6MXVB1tJM8UCzu7RXdmPVWC+y
ijWdUb4zXfZPUVmALCpcOdIBZLGVYsLN8Gh/iK/u9JABYpRPioOEE6xZN7PKgUjSRY3ZpfrAjRg0
O7mOSDxGQ7zOAAuLah6Y9sKujTaNeyOqYj+BDOrPx/cyH1ISwmKaqNUuusiguqxFnoEK1lBJXPoh
uGfgiwTJQr8WZAfMmTDdcEBdPkx2kFdF1PfKnN5dzO27dB8+7fVV6mTPccVkUZF665zwPfHPznxn
Gh9eoyXCUuOxS6hFa147O9NWxO4XR1XcD94CRUDEtKT99DSqVEg/2B3Xb5H8aeBjMMP9VNxi1bdo
SAE98MJ+3PJCXkwVC7cVZxz9tcZ0Z/WKtdqlYeuHS9LCM+M77EJJMrpF15ZdstbUN/ncbLSK9akj
mU43kMVbfjmNBGedvec5ocBHAOLNLr1d7209lwAjh6jGokG1TzsdcqB9NlRnpA4ss30BCwD/6Bse
kzfP3wfAJ9JNkAMHf+wvLWfp5pPPlrXUSqXOnKxca4d6ouGowieJRVN32RQRUeC55dLpu4N+mj2g
MNRcUG0Hj2K/mC9+NXN/ZOuWcxwIof9BbapzcV0WZ4J9JGYLdQezVCwnATqaKdbygSmwe0qDpDCn
MIT0sxsyAPYwBwT/EpLzCGFQGGBGKgrriirUXIfuDiB+Zal3qt7MO5cHwQxyNPnDE1Eed69J9sMB
Prrw4YOdhG+eMsXWYAR8j0ZGcwAH0VUBKkuurhwCmslebAHjxqTZ3KtiRUnPQjh4sYNYw7Lkb7BA
GJT9XicbymLp/sX2QTrk4GlQfFW5x0/VM0oCWx0MfJ3Eu2hdMj+Bp02w3p/JtHlCmXKlFMtSEg1l
x1O/2KAJB+4pjMTABKVe730iTEPxgaceececxoYBbaCPvC09PzDzSur42u5ogi7jF3eUU/5ChEye
7hOaZSp/WJ6fBtlqLH5ulYYVcXao/VPmyJc6i3F4joIOpmauYSEt6UZKaNk9ebWGuH+jM663ij0k
8tZhpKC49AAkbWYbiOLiz/a4lxbb5hgrcrPBogyv7AeJo6gaAfBhGpYSBqLltCDp7UqN0e2zYJ6Z
yCWYpgWWHhx/k387bACWcXBUrJcmvcCRaI0kkrGZNqaEslvqiEZjiTx+qkDQoc0dCzEHZ/J8GkSb
tHkJ9u9kydeUtm1gdM2QQSv2S2zcWEFi/RHk243HCnIReaLmeGvMfBYMxjTtiDv7SOd9UmWIa3dF
oRk7GG+r/xf1YcFXjI+u5SepO/EW39C+8wKkgfwWh0EnubysF3yfMHGa2Wh018ON7l5gkiQGlGLo
2zHmKvk7f3jcPbzVd0/WoypJJtymYmg7IK0lTwa+irJq530Kx0U6ldZWxVWoBgvUu4WV6uE34FJj
MiJhpRoyHJUkEgYMH76h9fS2stw7pRSNZ5DNeCWjAv1oBv2lslZAit5MTIeHPMVrbnycu0DqsJ/5
r9Qrq7KiRzpGgsMxpXGlcYg0UpZLqTVyJqD4K2hqkdKm7jiXNflR0Y2Qy+RBeTtbgMtz4nJqXflG
fqPzHLaVeTHqo3fZeT92pOEtXx3R2fQzGy2TDVnjFhpNtZlSnPs7i6BaL+biZ5quGiuePCXDjupK
Q7R85FGbb4hoU7KhJ0RLR+dzEuGskWfR2YNrkJBkXkC7E8d0/QSSz+Mt53bAhqtGv5mvsddSZusQ
z+bQKdOz2y+6eSxHeAwQy7eNtzdRBaFGPIc9AlNnvD2Z7QWfUtupFeHeswlV87tu8zPVVV6hw1gQ
KKbx2UJbo5YUnyr+0gaPHJM0xhk2T1iPNV1M9Yoj4p017qTxumuWLV6qtaQo2RBQ0vIhDyykyFET
9mRUG/+faGo76u6IcEeNULK8TsLrDd+oVSZ6Nt+yKcg9LQWTJshMmNM6I7BsqhLw9BIb9doR/p9I
DrhBDe/PBjK3GpyDzIyVTrTbMtaobKEz1f6PG7ubk+4bXDBiZdz4VTs+CvU8WnEEWWPtwBI6mjNZ
Wtm0EglWi3+TZJjNZNu0cJ2MSPxvt6XU3XrZhoc+D1Lk8wYm56k7B7byjREiIMJXwR51xFT0K2gA
bmQbyV4sgY2vaGjajBz2kJiPLTk2Gs/rF0qrFHrYf9YMn3UnK8NjJkKQiFwSwf6zdpAQ+Wqiiadq
NtXjlSZYfUvfUoWTvRexFV6Nl1TTNNCHwqPFpuqrAgx2+0/40QjVRr5AMWyNlL+WsNxiZ393s/1a
UwYG1o+goHOAvMkAK7i3h2+V4jwll9lZyak5Tm3G51QWIZu7FurSBAoHkFYIAr/CBx/RQvktup9G
eJ87cFMm8oi8DZvVDM7RKjJ3pRkPEfKEZCdreYoe3Ja4h/mwdXEHaw8apleA8lGN4uWOoRl6j2Di
M52P7yYghWOBGTwRxJ2ctgZvJId3bOo5FO6JRffPnAXfbpljhukJkw/ti9wGEY+qv6fu5eXCdefG
042kTLRBQaGccuIibhaK6+4EqyR7br9w/FyhFkcV76fVUtwVjr7jkejfeun183x9PImUhIMgmOLL
F+ubY0Ae8jWkRdNese1/qWQ4Ku0IDvgav5ykGuPRqNadawCJmY/OfpZEaMoQjd3PPC0iYAtqBcU0
jv57aIzU47gj4BaCRR8ZMZPNeHVMTPT5NuJo6+PIiQgKEHDt5LRfOKlPw6i7D2k5b4ZOyohKuGHo
xkyD7weSBKp9ukGSgAHJBw/fYKaKmD76IjbvdFxLwAuoMytY/cuiTtcLZiA6gmHVtWW/+YItN4J6
wK+LZMnutBLo7jx0T5d6AoKitaIz4viDbrEahCLOVyeTqSAxhDQcQbCwrHa/1E8dS2aeBbRWPzeI
ar8cnU+114Czb5HerzNYC4gn+DceJXeQk7F1h6v/05s4o+d7DXTxYW3U+gJfBWWIdB5tZ8DTjEaV
XOB7CK1V16sGix7VXVUrH6jHs3emZ8/7OjUjrQsWGtY77ZvxmRngAD8SMjYahz1uHNan89X9ij+d
CqlCscCK4h47XDcD9RXmhuQyIRZ3y5hTtB0JZIqQWZ+Irn2yl0l86rJthcvTpJN4LbVhyNyHZA2F
vFO1PqfXPerjL2JqZEcmmlWVrZl5oEN36weERIY3Zo0ZLzMgcFmS+e44CL3PqdS1wSPoJiN3/Cxd
Xtj38AWe+WjOsCGh9RyKX25m+Z//gOvVFlWPtJor9PjrVYoXLTOAsf7dRdpuQ4IFh5lXS6tSp4IZ
koeLA1BrmQLMW+EK8E5LpH28S0bO0n6IWErlpaqN2oBM/qlBAiUgbZUuawn0hgD3lZyXhDbgPH7b
3Fv6LsFMfhxHqkWmgHL133oIIWycyml2Q8S/gdeK1bnGAVz+yp6+KKc3ZaHhyyLtx/dY0CIbe+j+
YLvC0QpT/ooGPvVG+hvkrR9+aGZZPzigqzb1EPervcyvh+tdcr6xu99TRpb08BfheB4FE27w4eJg
MsQnTp+Oae0jpDubTwesFHDFmfiHZorjbL5m1j0x1jjsmFAVlDfFo4n1wzWZYqRJqRFVOV7Ae+Rc
xjJ8LBrC75kzfqcg1f8kX8evhmYHknUMyDAs/YrD9EPokUaCmcRDx+uQ0LMiyTAQlyQoG0PUmxjW
wEtn5pROL5EoIVjtXVNBAN94cdmUgY+thADol6ThTTRnVTNOkHmt1WJB0wMWmvzdusDYY1gPTExv
mnTWDsZKDlU1F8Johy0sg1ZHyoG0c9nzr6DkevHPj45I3c2RMODCFKFI90g+4yDAXeMcdi1w5OMO
n7cEWiJS99R+8nC7eFhjzZPS8j6tL8XVOB2pa0VC7REV1IHnjCZ+Izx0lEYMdHxKx7EAlxkZ9QxQ
tcBD4/OH89yim0dU1RCFAPVabjFMVFPO4gxHfkCI+arrICtJ9zqGJYWweWyYAeo3B3YB7PmzdwlG
4e4exf8OLt0eJ3rcPY5N39piPXegSEYNlil/s8FKpwQeoMBELBOKCnvVubIZTRJhz87pZ6JQUChT
ldHbZMlWng8eYfuHdlHKOGaCKEyrTPm3+BsEIARVz3FMGow9UnUzBUWyzUEteOa3pFcLtFrhPfTR
bgD5SzlfC7v+qSorvWKsY4GWUibSdfdt6wmh7CE8QKuGTQqPE2gUNUEKrfw8xHrL4ymBtSU5e30T
L91MDQ7WYfIb8MyI1sJuLc8LJGyTUAr9JRJmyvadailRcYhyYSjnW+/pRcM3gJo+/AA3Sq++nCUN
B9KRZQs60xETs5fG9rbvqN0751gvvvzVCTvq6ZwMIIdXhS+NRNdObdwkrPT30xShvbp2TOBZOoiw
b4zuuuGYoRJuBjvnDY+t8dIynLWx9P1esEfags76O4+FDZuwcC72fe6xLpoRGG2lGRczm3nc+ANm
/FrpLkW9UY2xO57SDP5AkH54X8ijwRUJ0N7+jNOSTckXNtKg0TVWFMwVPLzLI0ouLyR7/Pp3qYUt
QnLZbCdX0u4JpgpKmi5/wezglvZD2oGWh3GTef31vgUGxH5y16/zktsFJ1Hup63VGYVV+iIp1kI3
sIlDsZj1fDwhJ8VbH8azK0WUUZrj2lt/p4HLJQZhh4kSQoTrFiHM5zj9zdo7qgCRli0tI3P+IAyF
Omz8ts0DRSg68YK5owqwLYZxG0g1CfMyaq9Nxc0TGQiOjI/EwCHjJbHCYrnPNvinKTdOUiZyOWae
jxdJbSkwGvh5P/nNsodv4qYqOE5+RH8AD3bTClIvxhBpd8K8g/Vc/E2T++D8sEpLfcGeTUgVoiXC
V+dF+TuLWbyV0xPY9NpyJaGMVS5owrdDTCwbSzcVy35tPmL9L27XqLtAewd+/1eBRj2PejhZWy/B
FCp+Z/XeqfgukD//PxyasazRhPr6+NwXj0EnWbCrOWLi+dJ4Y5ufRey5SWcZqK7Av3mpNnaGpdbb
mcU6sft/XVaxJVzE3UrulFrasw4LEOX4FyqjufcPDKoeQU5dMRZQyo8m0QxABiLeQ93zjAw/zH6/
NUZc4o64++uIDh7F5DOAha7b3FhsM7SH+CSabD1k6qEM9y3JKLiKwxuRuGfMlRgpnXt+VMXQ/2WN
7OqwfaMaCh8e/SA0uuKrMWllSatO+/pABINntpPynZABjeRo0BUurkitVp+gF4PhPDsN9Pybiy3K
FeD3Wc/1voaWEDYxOTJaQ2UPzQD0kv/V2Y/tu1OO4tpncsPrtOu8RjYRD+drW9xqjCXrkdTUbaFu
+n/ns0knCwjJVvX3sANskqGLw1EiQZmUI2K0zqV7+8l8TwpoeRlHqcVVXNRnqkNZmmLbblSwglEg
fwXlTXJzYqZwyjoPpGuClQjYFrmVS0u2SiUNGfgcgo3xRqKn1g+T9b3NO+1hSJof1HE2SN+dm0KJ
YwKKhoKoquiN6Jz96e85GDlDscBrSex1s5iHjcbfbaPtBter4iNObLZQaId9agUxDKqApm3ffPOQ
4MpAKGqyrjnct3Diuip1xc+Bjyy9x/utpAjSuEoqlLgi9FG7qGlF4uI+wDISJf3zkM3e8PfyHPjv
8HSC2H9P2Hi8xM/NP0LlyIKcDWQWqa8NqT+3jBLtM6h65OGzXDblqLWZtEU4Suxm98fPK6NPZdlR
nT58Uxl7SP3PKKmSq+NdWM+Dk7t4bz/x6bQS4K3JOuzN10t++B8QWLsBwhjaPkpiZJO1lzG2fqzw
uwoJkJ7DFbcioJMLaJcUR3cWqp/OlgCCHYssmImjQog/HR/RAoYtchveKZ+NgpevMCuclG+DuV6o
B4psd2gsmIWhiGdr4ofsaZDWxqJej2OW80BP3zkkTb79Ce8aBD5T8hx7LcaV/6AYly8PJ2zb2eGE
yCOb1jASxXUd9ZK+JuyqwEfj4nwPLk1Z0d9mzHGhfaVB4ttUTsXduSsz2ZNIBTFCZFr9v2uQ7hhP
w0xNtW7bsANqWj/HXvceghrz0TcCGGa5K6Kmkd/wqq57y1xrukD5h8uR2q3tn2zL73+hknn/aRYW
a6jbFfHvdr8tgRFgeNqYSJgYnZSrcQdlMqAJxGNcQ8/YKwgQgP83kYMyD9Yk+2mD2wQbO7R0R++I
L8LpVORmnAxRjIrywTcv1qPq4PAJ9xwg2un+ODaQzlpSwSFgLOP47JeA8YA1JUj2e2j/2P1/ECPT
1iAetc7L2c1eQNoO+YkvPKWzrXdY/maCWwemj1vs+2yDjp8dFQmehRkYV8L+kyP1UCIF6EFJIhIS
j3uVdJvYOdjprzr9+9kr2A8sC5Su7HsHjwYhohNH8+zliyHTaLuvKOZ1TyWQWqUxAp5USZ4+PvO6
VfGdBxULgCJpkW0MNs831LFphfB5HpVSLi5h9bsig/os9q3WCL0WENOlJhi4YAguh+yAhwgdE5Xw
JEZ8FOcus7cl2v0ejtcp3Pqv8h/UURtllZ5OaUnJqtBQ8SJHAb/m+/VR2RCAFUl5+EDCGK+w4LPy
gDEincgPEGEoPTVSIeyRZ8sKIif1NUJ0fQzAlIRzhvNsKYtnGI3x28fmxT2x0DEv1resJWQETfIw
2JR5jnIVcWrE63q6k9CWf4ipVmxAwRQD5IgaR0QcXnh3UILlTFc7KsY+hL7ahJFWXoV6rPVL+EFB
GuQnIt2X0MTKC3QqRGA0diuxKgaaoFGtwmNerL4DuBGVnHqGzqDSnvbI04IDWWrOIE68OH6zLWQJ
JMyHxGXPjj6GjIERnvR9V2WXuNhL2P643EA5XbfVO0uTRb/i44anSNTCr+sqqbPR1RsSt0owX28r
iy3zB0VDSu6MLFgBptic4AsyWmT+9hJew4U4Ao9cjSTdEin7569nRVHi+mSs2LctqEDphVJ3qktr
iRCf4LNLiHfPemALIDJ91krhRrJeU9wSDr14QGj0tDbhzZuSZr4qiA/rsyM8TGOMFSUYzpWjEYGQ
GZbaQ7QpLLK/IRVn+5zqjtKJS5TEhL6Jq4QtN0E87jXTaXO+H3SZurqgCN0NGurHYlHgpJuxVfcc
FrvZRxSQAKw8+N/sNU6Mn/PCVUmWc4kcyP3dgPApXN4pNK7XZy1AV/np/o5c2zaZAAXMDqdGvN8+
CQv+Tl8L0reACotSAhArXub5h6NPTfZdFICuzpjzArHQcc+ll53hKPWsZJDO8M4PBb1SV66trpdn
oe+PzWSvYolP7yVkuX4NhNMJhmOJebQ1IWuyFFBe091VArqtjD4S9ixhmeR72FiXVZKmx1Ht5hdW
oc+jigVG5cmXWe2/OF64X4VLcNJ0iOeT7htoHVp3WVoKId5QOdN7N5Yt3r6U4DiFBxD+nXu88ndH
wQRYMAq5e8iWMDNQsvmFriROIwdl9GNWULn+ZadiZw6M/Ng1cyVJfZkpTXbgsZ7YQfDw2Zh+7NHb
X9+hkJr1gZDf8C1ehYdHQyb3yB1omQqpMXnJ+CO8cG67An+pYdNyqOeIpOhi3F2BzXVA5BYtIZTK
OJGE449900WqFft4wdCHeUx+uFYKAb4EgG3iKNydGsxx0+pSk7TH0I64LtIAeFwZ4KgSh9/nKsDj
3kM/mCBnJmH+iV2GdXumh2hra7EUUhn9yKhnrQkruW8igvpK0WMWCfRK0xaqdRhHyOzK2LKNV/5r
hlLw8TETGCuBgzoOltU94vXSewVHbAoax5qrpGlzlN4a5F2jyJSpuxrbuUXvFE8FwsCAoxRNzNxR
x4A0AFF5tiG5kZigf6XStVvozEWbjl8BHIelM1MtI66gAcsNdfnc2k2FaafulOxVIXENccZltRVQ
FLFf3AzusmnOvRmXFjuv9WbYVJ7OXt0MvZe0ctBNy8mO41euaGY9VjEcsJqNE1etYmunW3ve56YD
ItFRaB+9eD0pP+eTsXpXELxHvptgZ+faxtrKVndolHwsN/hF95AxAASoQGo4PtLwyk/ZYeBze6m+
muWNsEumPN37obPLfiLlDF/0iq3nO+kDbGSyiuosgus439pbib6vRFYA8YA/GXKbhr9T/P01WK7M
VhCNEynzhdvtxaiQ7Fd56/TDYXcRBsA+8NaR1EBzH8L0CabBX6EBbElFU4iAIUWQpCfiuFxMQcjn
rQTkyQG3IlPLnjXBg3XfGcAIux1YYJXRpnJu2sH7YhzrzhVZTGUfvgf8+TENxgZGEXyvVrHy+MqC
26RqVmqLk0CsZSjHjhZciSBTrcJhEPM0+xrmnLAjvMxZgaTCagwHCm0L9Ool2AqkuYZA6t2fke1C
MjoElFAdOWHkQE8JPxt8I6oznHb5C5kJWvBzY2L+JgSFXuh7TJA7KqxpLBOgb1e1pyhyunB+yrOB
oLO7tDdDLx2CPuA+R7L/F3Sk5VW27hZM+Uvmlk/6x2Sc3dCMN5/NbKoWooWcduxJFrbMynG3AVvh
pqL29+OpPrhNJeDebMgnXv5SYt9xBGc/OKDbVd2EKyEUngTrZiiQxwNwxnR33qTvRAjHrJ/CIktQ
O3nnIHtD45matwIXekQ4O6KhCpIBn8Icx1VN2QcmI4kzbQa89Q8yO4/muyNFhts/J21rf0rQg72G
ljaP7G2enIb2bowDfn9GvlKgQJG3RneTDGzBWhlh4flAxChydLQ8vdmDP1vSyuSxAopmDyUmOFNr
qzORoL5sMyDpLezGBvLMtFeoH43Q3dpCEznqS9AtdnhnjqKzTn+tpkQeobAZ63Vnsu+XISUfai6/
n8lyQfhEoQ9ZhMcOEyxb34JILGJB/rx/3csCHs4Jq8GP3eaPUBlnx9rzKBU41A2dRZi08AOaT0M2
s7N7c13gnkJ9kRc0MeDUxln9lbCMeHX7KU5sopHkPXUfi9jVgiAaUbDu1GWGlPXjrjqc8S/fhNxa
CztO4opHbdPrEnpLOYBByUysARy5JE/DqhhbgwBVDQHD5fgzZ0iYRFv5ZhfFlg2FqXdq3YnFclTI
yyJvt20C57P3tJ2FSGanypRSI3dJnRo33f1UG4A8Ai1WiI71DbT8GYJ9c9F/zJzcw0wMLcCEmpMF
meL5RKz8fcpYUNQU73MLJ+lVpDNl3f1d68g9A9s3O2EMnsydR70SePkBnCghWsN9Y1mUeLsfnswo
MpElH6Bqbf34ips1IACTxIbKYNB8CKa3X/WjMGKbR5IxqkQdS+78HxZYFmHM+8z2jdMmYP2QCB0T
tP/85XQC2QWDDCGkTZTTfNWux3xOutwXjAbfytQmHWJXwbuDojpBXUVpVZzSjry9R61aQ3PWIJ6a
y/hFPJOGz/IsO1YBKUiBTkyf0X7lJIsKyO5os+h1OIXz8Bv5j0pSRRCZaeS562urg9eq7VxcZrIw
XCyY6kjEzqh8XThSDon6sI4VP7II4OjyRSVEXR7jQKPOPfUSk41bhm+nvBcNddXNBjPSgFB9MwrG
xsDGcoTfsHnGM6BEJo8688X/TX1Pc4ILDGUdWdi1/sKW7gXZEj2NuJOfafLxLeDAuKh8wjHeDASm
xjyGfetOTgtnVebqf6urNsJhCAMcr9B3FK+aXXgdebuRA3v9rWHVRebZKw60EMXAYlTUUISP6V48
LSNCQDssC2euF7xAVwFVDMtlA+SNtSNJyscD/wDD/Dxo3FQfaaSQtCwtCQ6OXkiyhqSCdU7dKfKX
qSIxXadIB7Xom4F86zwCbm9An3T3VQQbDtylk7RxpKifq5FTAW2fuT2DDlNByf6zDF/h/nPTgPvw
/wy0CN4ZMqzm0WMIZXY+Bkt11QZcgxspu5XVgpGWiy3F7c//n3/ozdmx7M/xEpDMTTaoGgCOYPtV
Mp1XiLrwi/rFUYWtROLPsYcbfov+9/cGt+xwf1F/PFQ6SMjbSUgnDzOluGEyd+qCc0nTsgO58cF/
N5/AKQRFziUo1KuFbrYsLsjKK3SUAg2OFRFyMx1qcuIzU0kl5su8PEZt7uNckDINbjfU8sT0cVD2
p5RlY4i84MblL+CfdUkBGutDoOtJdX1NTz3Wecnats9QuS32CABW+ezR4MvDjeEJEKMSF1Ul2DJO
0l/AOQVPKo60KUTM6594BMhOpZxmbi0HS0usCUBbRLp9kWPLm0avKiQstinELmbno+tk1oAbJVJS
S2mbV4tgYsNSfbx29Gn619cKAv0OROkFxve+vLLq0AuKJHEIyEoUdI/1UE+057YRj6exMO8UfyP2
bHNzxmR05+mPD9FOE6cM53/EojULrXQwdGBQCwEEocI6DvLTYp79EMHYmmrgFWA0NyrCUu0RkKqy
B7fuE7C+JEiln45Vav3xzLyDEylNyRRSIUWsycA8Jb0E+gdRfEfx2NENSQB/iTtHL4q9pmZHb496
D2aSjav/XTwoaGE4hVo3xjtHE8RkZ3guxIPWrNfTH0GtssH/Q4DEF07UdZ24gM1CL5Zpj2cEkGhH
D4DYb9c9FBOfda8f4a3xJTD3c6bbPxfSZydOkUjbTxQZbBUbliaWZKKYpGPj1hOLMFjeg9QkAa7h
5sjlaOxOGoA77PBKIv8BbzkEXrz/6TO0On7dCWcuhIlYuIoszqdbZ7yJ/FgM88+VM3b1qUVD/DFX
cPElIC3HwxbMhyH1HMtoHFQfKBDhS/wmIy9k8hY9AC8VxoZfzbims2Djz78R0MzQ4G5vDMxkrxsA
IbDj9gH15tLst9BH5qHdcLq4kDXQVAsg1y2SmAZvt9QCwOZekCkYqQ45o8WmkeEeT2mbo6TD5sSf
Ii1zGKJrTEZCwXpd/icHNrkMfMCK7ZucxjhOYIRO67B7uUpqbIQ+3DwGhRuCb4xNowAm3euBHtq1
0xN+ZifUS0jf/+tfW6oro86u0XdF4qF6YUBBgdsUoUcmJyJgo2FLoqHWoAnkkDycoA9i6NEdBdbp
chftJ7nkV7w4hpwavk/ZmrO2IDFrMY5fY45cfiTGmkQomL5gvST8bGD75+KlEqKQOgz8PnWPu6W1
uBtdc1B5t8iR265u7iXJ/Av5ryfWDKXcPXkvRstU5HKtUCPaXw/wbNtx/iF4znsuKOF5O6IEcWD9
bH0ifUB/H0JGAOWsiu0ptlw7y786yaFScggFwXW0nxr2J13UVFerfUHaCdnZ6991qcoMVzqOjpn8
ZHpNcfS4VBnsOkOFSAD/9+ump2XNDINlY84iR19KvxabvvSvNWMxTbBRXz9EzJAsYCTRe/PAX8Lh
ceIPGToVKyg72fRguRlGe8H9zGcgqrV4rI1psZOeSzceaaW6dHptFFqtZr/pJdSEw3HnWDKKDWkc
qP+YBLQUgnS7HzxsXV2aHF/946Lf8TFJxQI2ggtKGdkaYawj9kj42nHhLcqaqrguo6VK3bbtFfZ5
5Kq/kX8nGKsELDdn+uIcFssPUCQn0ogXneE9zDiMewKXOai5RGIP3h1sa0oosGUKyD/ljl/Oz+oM
Pn+U2pbdI0A5QYNa8iMdYBeqBJcnMl7qWiVlJQwwQv+UY0QI7h4yMzyzD9JHAzO61kKmDdtQ2dD3
QJrYjOCWrCLQkOmQgY/4Q3GM0M+ObrrfkyEgHJi8zPCnRRi2YDGyQxUvFdnjhbd4EK+XkV2nKOXW
hC/v1BMSXRG3JmUp6Hb8MhbswLO+h8ZK8C31T+ab5ZVcuB8bV69j0OhwPZJQhHXp/NtBvdgV1bKk
veOUecpr4cxRwS62DU7YxgDOHo7fIK0f9hdQnwdxOaDdCbtetWFusWgQoihy3lDVf9RLugu2yOvY
T6DYnCpswOyWrQP1C39+5Bgv3NPyjy6p5aqWLOXGSdEvOUxD+B0wuApV/tDwyqKI35Tv6PwKC44n
PiDeIhmu0Jn0IvjYK6iIXtfZkCl+PZDHmf53F9juZLBqGeCq0hwy0bKk8OvkeIMvZMACO2Qvlbcz
3qtSRZeKUXgGpXO5JDQmXYC5nJlJsnxF9jZpHRofulNVXIndbjJKmFmdFlxZX66dPfcdvndrCXd8
/t1og7KIwt2raVjcp3NoHO5cssyLqyXYCkZLvNJWHi4abx9XMJtqlpezzHHRReCDFsZBXJKz5rn+
n0hbE17Qp3b+BkRY2F9g5S5o9A4KbFhMYtKI4QpgeXJw6ngcoBFm3W/JPPFH4uweNq9Ua3b8kV9j
NQOsv6RE2UvalHHlMJ6C42tr+2WDf1/Xt3gpkcyrP++RuP7zb7a44IwH/QIarWtA7O/sXcaUljft
4mFXfO84QvC9dBSxNtTKaq6aNMXx9zgNknd26oJCZ4RleHassK11+oG0MJ2hktzRPBhHz+Pt+ngB
MfXghumwaLsbfdhTu0r/pyCRrhTdyCDGZ1Q8xFwZt65VP1qB80GJ1Z4UienkoVkzrfpaSgzaXRD7
vQDzxLMMFsONpsr2CbbeQdsswRoJiHRTKcSpPI2pdyznllzOZ1pzpwYV+ohatJIZXJLYK86sOWHN
WTfvefE83SAnTTxaHOfZXmwqj/2XOy4jWQoPnOz4IRCILeRoHxBbUMxTEvrJls0mRD+aRpwKrunU
yjmZFeWCyNpcillGewDObfmrTH745f8nhGozFTaqGOlNI0x05ZaFpjZoNvrih2vT02/0RX2wnGuu
x/4ytkTHRJPy80L6BUCQgrK18e3Ak4dSvJk2qgxmXVvFXtVymvgyGWRNCBwB9kOe/RO41cQc0VaY
Njq6+jFqqtOuwidQIOvkaos1Rd5PKtRP4ecmz2D2Eo8jxIEaFmSLwGFo0VJUUeVIAy7Tz+vNwTjY
WpGbZDoafCPH6xpDqIjyKvbbpgTOtZ066kfolJQ2BHbRoiGJPxF7jZMLGvl/rinslwQcbPA4hDI2
vk0T+HTxT+M4nEI4e84aIMhwfcFCiOBoVsNNbaI6LG9FV/b6+vtX3jBJYd/sq99K+/6z2FGonPDp
kO2rjhYVxV8yB4NN1WtR65xZ3v8k8PkXH/zAtUMIQ5PAifP9MqLLk3Aeyze9zeiUEZRvdBG8Y4FX
BFv0emBRf/2TtTdp1NwMBfYy1cw8mshcm5ak5vVfzC1OMlENVudLyh/cF6+Rf+Nf4tjjl6IfXx+K
uBjrXmXHdaU97JEJknnm73a5eOyODGysMCrPez331X9la+ob3BoykXsFdF60SxfmtKevpixg5KHP
ECTk+96Klt/K1Dgs2yoOifGJl7EF8X1enrU4B90+oiu3eTJiZssD0mXNz/z/z8pmS6wfy2EtVfgj
hjmnTKwuMWhT+jF6Jo0UKv3sk6CbJzQ/pUBqsQoC/PzBn+Dlk7IxMoymC4WAsWVrw5Y+e+JoxHD4
i2UZNqTRp6hliqjzieElq6MxU1o1nFW5odYLze39WC7kk7/bqNuArUo2Pq7qQ5uVq9wkNAuNGi90
gFHYLgFMoCWDpe7+fnPJ/6SX64TBVAEZ7N54ymP54MMqg1M9xxTgDTBKpztxv856Yp3sAzu7aS1I
OoWgrAsuJncal5l/jJt0H0sozpT5+++Z8CufNVgjVVFzH5+XMcBsSZE3CmAJBw1mkC+e8pyIyn/v
WmW53w+Yw4bKwCGkZREcTUVS8NwboRgfmB8OiMXLMIaMxYxQdFFb9XMbs0t1AJ7M514YjtfxK2jG
qMnkZitrg5PtWmbw+17M5F6kP8d/hFMz7gYZ7fbh/O4saV/4TG7eVktvoel3VfJqXFl2Tb1BlVKB
yRRIx3ZWpAzyeDgDzyU+VYqkKe+ylNYFAdS1HYgeb7CFK2WkyVnZa+6inwmMr0uGNn+x7sMoL3jR
z886ZRJdccV/lUs2wXYKZ+jJUkDxcTe0pJ0belfGHywKswvvSpPBnxLELh/AllM/EjmSgdwTgyl4
ijn/vNHtb5+KjKaaIRcQwQd3dGkNoVbXOpbklI+P7zWrC8gsCfRXH+u3uCA85qe7l4I09V1dufLs
hZdly435yDyBrIvht4pJrSVn4SoWzJVCJpJvXbpaQlcP88oxOmWvUQ4MrIgtOWBYGtrkZObRkuEY
+yFpoC2DcN1cnD3owAoWfVntwm8hqDrIKOP3ADi2Q9+LQlCEGdeZFXWOpA3YUP7QTlUuw/8qcvL4
teTDTzqWkh90YuuLUHUPkNtBzPDSwqgN/D/ThIn5eRtMDQ0wH15/ve8J5sbO4E0+K+PKP8M571Ob
PvipnMFu7RYtq6rLD7uEcG6Snn7g4hvVoYtbe1c3nBm9rV+uBndwfVVh5K3/v/isl9HZf2J3Awa2
1oDtF2QNUg3OYcqEROvL4W13OVBhh0mn/Kxj3R1mdboKVwFDnoZa731GfIu0Nq6K5R/6DSpXt1bv
jXyk9EC2hpKLq7iFGtomVA/mWbUU1dVuoRbULk/wJGhuyV2V/eXedVxmNqwsEarG3dM6ZLLUJCMs
kyYfPNgQ+iS7pERcGYGS2YIG8yD/jW+QPp59XCQSp0EfgTmEAEXBAfan4mKlEYnBjIkIKLoSgQIQ
qVQk9W823NWGEVI6KQbyzKFUWwMB3ypVV9lHDvAI7jqoVuUSk8GvS2gQ19tJeduBFyBOb3wVr+ej
vEPTVCSMNRdThjwoMTrnQqNINMfEt5dwezvCWr/sVwAPdUS1LPSd2zo2G6snm3ZnATXydK79YMKH
PU0Z8jHAhbbDMawmr6FTtsbmINkrvbxDx4T6MytHSIBKZrCgBT1j50e88GJnGProU4SETjrsW4a4
z6tn5Hw5B72778cwhCu2IgHwJBKDWPnFrOc/HVuNQP2sSh53+M4h/kJQHspcw4BTDkbOKnGnJ/qu
z8u527AGShZ+q3yxgb2G89HoC67kVzd2G2htYIr5LUDq4l/vaudDCbrFyDlGA6o19fk8YlIHdRHh
l/Q/b+So0zs6me/CFhONdnE02pVYfpjdcy7ju95iIKoFUqeRXzMOwn08DgyUbK+UdiBEYrcVNpqN
Mf1XPh5U3Q9376l1zkud0TowA2EmqoBShRoN173SC7otS4ROhY1FzcXH3oXPmj58HXzMw/dVyqE9
DTcNvWKH3+bGsMHoxWA0CjhCMd41yENyuPzbIE6Jzm7dh9PnJPxHbaflPtqYU6youx9D4T6M5HG1
AEudTcBhBhN472UBUzH6v/daYzAeJV1ggg5npZp0FVF0z8FYkNGHGdshTZoRxyBu5rXGpra6M8rM
C+fQtEMGzj2liEMwld4Nl+pfn+M4YbPwLtdEfVxFpGf9R/qVMWiLbBbuIF7jfsZZlyWuY1T9VoM1
PBX3m/yEDpJjJDVKJ/vUQRaMLQhZkl+Ifpuiw654VlvBXu6X7m/uQVhDOAB3Wwe49uf2z/F1iRUE
ZKFHvlhGaO3SMotpbyQuBp4Y320bohN1RAcDNZWJJ3771t51nanxZgTcfgrIcZpoFwtGXFDP0MTg
zTLo+x3vWx9c5UEQ2/+KkgFnENIBvvrCDknAUtydPwYEmk8zdxI7KU460JDDsaFkRdg9cFNl/kSX
4HmfLiO+Z2JiR5zkhOryZ9r4JJ6onfSlmM3m/l91z4dhFoCjIzz+yyfZ9Qr5npFP58ky+6HglUXJ
HTpLFncjKu+adCpzopTHqjyOjXh8N2GkIn0MkLF1FFiIdOBr5OB2qpl7wL6wqaAenjRr4X7Xg9Ah
TDWJUplCKdweRNt1fyr3QCJzUjP1XMn4MrH9p4W6ufUkN75SIr6L/15ZmbU0QpUr1fQxAjjR3ezJ
XY/cSWGbj7YiIVzEc7V9hxJvv+Sc8yDwSnpRC5STbYlhGZ+l7YxbW4Ke/C4StpFSEfhTO2xr51gm
ZgcQKItKXWHoT96vVDxlvAJ3HqjTis+erXqjHLbmmiKkTOXhkttfV90LCt4PGnZoEUYIZsa2e2Nr
64n4MPcwGoSVfWAMjCvGPI5CrFmMTb+PQlZ+Dk/eS20oFFml15kouWAuSSAf0bzX/Vg0IziR4ZYu
TIQN/EWyuCe8OO3qYoFXZWllSBEBZ2y1VqgzuTNl1FM7o03nYADgmnn0IO/9nO1UImk0AgyUrutg
1y7VIpgjh/tBLN7r/M/IP2wPpvBPLNk2xKQNb7+EH8B1NJzhPh4HT47cCMExIMnxIkXq1j6/J06i
Lp/qJDVYr1Tm1KH/G3sxJBT/xlbRSsVUSn4yoss+lMDkjUJ18rsdBEzv9DjU7CTgyYS6Sz6IYbto
5lagdFNNeijKpRXOqR99nOC6sHNYXEcU5FLOUM3P+xWLf+yAGzRfJPTRfecHVekXnjuZwdvCNszT
YvzgN3uXuMwXc7Ylst8y3m9n1nG3qbvPsx0F1WI/2wQE+RHglHQ+4z+OgrwSmF1qLMXdx+PMuj5e
zOVw0U4MZCgE/xXrixOIjJuCOUYffwYn/swVjU7XzwVUNofQ1DsvKuG6Pe/u1XuWass/gnoyCe8g
tTkwf20IcNUH0iHR5BqwXrZxKg6/9WwMQQC/BY0Ee+0quaU5X5IPoybNfKdYWqgHDeduAOBUUIe2
ufk8YUB+c/KjQucpmv5jN29g7ndxujaj4AzHqrd1N7AGSyc8XObtSiUFnHfxM09BnCZpVn4rMqo/
HoWlkbrp8ckPBBa8pWVCLQdrVUwA0CiGzxAm9GwJdTl6Hx2xdH7l2MlZYA9xHx38rlHyt2Xc6eui
1ztv/W46z1bxD+bnvsViD3kyBIzpsjDizEHKfFY07MxM6JlGz2pj1gVqIJxnrULsvjn6+gQ7w1lD
7/soto2tiNyJU+YUO+l28Al+v2kzXarsS2x6AgXFwC/0mu56SEWsF+4xuUVeQu7N7uVAignIzX+i
s42E0geduF6wv55WRuiTzkQDBOZLdk2C00btB3pNFWQB7RWJgPow7IcZhXnGYNd1GHxxqp6hpDfN
d0K9dRQP7EPjblG0dAFi0gmr8dcgFrfLMFeiQeIfVV5RdT3xWXBf5tuNztgy7Gmk2pWYEDryR8x8
NMOIInJeQGgoDpgnWZEMts2i4WrxwztHuOvD+OZjgItHliCLvOxDG18drTj2VipB14FMpugvsMLi
fmO1FCJLRfC2gcaVUbsdiHpoA61ooB7ea/yLqht2F653arVHka2lZ7tPiVaTJU9CidN2Fs5DZEva
U3beAGg5bhZnFaJZVa2vf8ghs/K0gY/X1m6mS006fdjPXBcZAJooIi5Ny2pGttS1zJlrM9zjYFRq
x4CUCiKn6JwYSvrwEawWyVZdKFjz0jj/O+Q45dkr46lcJZTnQvRo2dyyXVyjAAZk2hDOAeBD1O2k
tTiZkxrfCYOfXzrTmf8S8UZS6fBIkkUMMQbUb2CpppJ2L4XQbetQT+P81I2wh5GhGvq3kfPlVM+5
7ODHtELmAEYntMYAOPGTrbh4EU50tQ3aVQqNaTKMxtoL2ajoRNthNipUA7z4EBwQLs0dMv0b+Uwh
hNy4HNeoNbl9jWd2PGeVxyi2mIoqguuo8ZxYxxM+HEDe8be6StFaD0euhpfNWjwrYv1BY8aq2fjG
Nuia1FHrTUTxJx4v4nWx96Bo1VWz6fWf/gPxKPSbkTKvi7eniDBV/xuw6wO0dMEXncSWk6Zmauf7
ttqbuNsU56GNFhtsgzHLSvpS/AsVFDuwAd1VO2NWRQsZz3z6e0wSXunnGtBIKaSNWek0rqaHk38Z
C/PhyGpDxMz8Hje7uCjE7TeAR/7TZwVpK6cEhFGHGXVmP2/6J4fmyK8jVKTPnd3MgmhU0w/prx2l
fYN95buISNhmyCuV0Av3SDVfGPUp/+9eCf+7R8uQx7YAeWWwWXSg5veqTslt6cnj2V0PAgpDo8N7
rVRlB6jTcxO19bIEg/r0x69zavOFclgY9/i7/d5cH8kea/wP3VEJDn9nKJeFKPq+WX2RRWUjrHRL
wL14+bKHLMOvsIFdAIY21Z6ZVpqjLCNJBtKq9ouLJeTPF+n0io9Ib/uOXEPyIbU5YvI8ch8N68Bm
+HYsX8axHoQ6rJVPE+eqseMFe5LxCxhqq5CvVGc6f0TapzaPYcwBOhmsDtwmThpdNJOyqbT9+UXw
ag66o3J9hPZoYp3V0sUcX9ZzrjJEj9qmySBJSOjWRLS6/SlPIekwmQsD7JIVSOc1uViIDta6C4vc
gXrz+Z7AcCuzylZv69lQRAgQsJU8eytIVfBWgdoBNrFZm9xChWpk8s8pSQyLZIXtBHrFy77/iHyu
LCVt+R+wvF2XQFUBj+gJfMOqwTkH6ghkJuMOdoHA9sndFK6M2kZL5ETrH3pxxzinCxIlyHJfXW5q
7yjvFJhH0FXvB6DfjiQDq2PZZOJYLkYFsoZmuIzTeCyDxI7NNmbEKcPY2nPSQ2PAY9H6eoDY39Ou
Rr1XmEMUEQT3hk8LmixBKyrNIKZKrQSENSeTDr4Nsbt1kjTWrCKdZYih08UCBzsXzPkkUGQ0apeR
FppxwE6svwnldOiyw5jJxcWekLVJ+hd5rNvwWXIjc4HAxHK08Zw3IrmeK++F4uKsnbNwpAE/uCN/
eKWNjImZ0bzCZFRzM63Va7VqE3Lzl5AY6MDmr5EitCl0ABOPG/UUll4vfje7DuoQVrLicJIOFC3J
tOHb9jOUPf7ZMvCFIqJw1swCe24tuGOvQANONzr2NiK5naz2S3RHWhU4qZiAiUsBkbKPbwka0sMO
vfpo7vBCS/ogbidvBhqJYAfAeVsVGmjfelDyyZqW3qA/iRyyxdEaGZK2bZL4FgOxoPqxtk0s0lUc
gZ5A1/i+zeoZ92PhqCz+vdv11BpSdf62ds6ekNDIJxh//Cx2/5sIV9ggw0ReFBI3PecTJ5nd3BMW
Uw35MXqO4aCesB5SYrQllsfw/kEjFs1DSOT4R9fBGCBzJMpSeD4vOvJJy9vsy3YA+eTF6QKHPHx/
0fDUc8Y2vLxq2rejq7JOJQbd04iiiNeB71fH/cnVLfQ6hzDsADcHQsmBRBEwl4BP2GmzjEZrMiZN
byFdx6ahLYcpW1LdEaEgznafXc3hf5G6E5EkaP/m/3pg8+Lcbw8NgObwBzvVC6lVJ8yc3mqMz0yc
mVwSB/MoNeyXq0wY9zjWH5VpC1iy2t8IuH3Ypd1ivGuUocPXdEfo9dTPzNSgrrGtWkfcd+SE9vbj
mHxuq1ocrIOHAB62cMUm9ZenAL67KGJNvpCnaKElUG3RNzvB/ToSf64YJMygNvNDvZ57q3tYZrdR
wz249njMHcCWlJPqqqpaObqeh5BhfFhoXRD8s5t3f+6Ig3I6Oyw8VPfott4JSMPNGDGbXqKGbZxh
KCBFZpe5jsBMv40QsYlcx/5qAViY39Dmecr4TIfVu3PfffVb9lQv8caCxrUMRsLnThtlEmQOTEuP
9OeISI58EbeItfPzweS55gwLALV4mFVBkPknfBDR1Ya9sS8y0IkFHwu2n9BlsQWlgqnmvCSFASLw
rkWYdXV0OloCzCWkxmLABsYUUzOM6PMwPx5MlAT9f9jdPyvZpVh64VbYLmNMn/RwwF0wdwsALUAv
p50xCqQanflwtGB7ZQTDSGTn1CgeMbPZTlqI1wV5Mtnt3KMCdbVnwl0dCccIM4CnnJTd1gS15uX3
bxcobBvXYLnOCDQQt3EA9G9Wu1Adc6+Urm5sqfhfb2051JSvm1den4QAV9JQJRH4yZ2/pkP/d9tY
UaNzC7xND64g1vbwX5PJLCbOSq2EEbDEtnU/aF6SarmsNs7JUXDW8CUTI8wbv5Vx7L57I2EJkCfJ
cObyTo2i4CT+zfE6ZX1FHkGMLZM5DLgYxvra1iV9Jmh04WaolP6xypHMI29ilcSPDqxojvz0pOc8
5DhrNN9ixIZ50Zy0+r2HGo4gs/2P8F3OsYLQbe1ya0d8P81XTBQ6FdBum+dKGJxHzdea2jKgVM1g
0YZQD+4IKLS04Kb6HioK2j5vZcGGUkMXb2M/DeDAC1B+jwysfmq/slaNR0NDMTfzvAcfOuQFCXPj
hVHdvfSzQdcN1JObrP5XORNGgDoH9mDndQnhi6KmHMnvoJaOwUgfTdKnY5kp95ruSeq4ROeBYOFL
C4Xm1lSgWItKDBYcGRrpxyVFAjcyhHs7HAcZL9nlGHikV8OwFpm71PcRF14hSCkjdkxySGt/sy5m
cZJYPn8W5IAGAjJLP3IWJtP5LoIx9KU+2ffzwZwndDGtGF2w6uvq4P9wCeTMkxE3PsSCQ6LxVMmv
+uZdkawf5BRUGWxlXYK6fsOXskkfnLob1A6zOuPUBKFF5YftnEBJeIc2nIf+yJxldEBMSNEmGJ2k
M84DcJFTI1P1i18tmyCPUyvW7aLFXPvKV1A5+c0DDQ+bjDYBO0M49gqR0taqSuGPm8cNYoLgwR/G
7iGs/RvEImEjhJNXvWZgOM/2x2XUlyk4yA41DoDzZrM2HZgAIJ6aprheoGAxNX+i4EehWz84Onrw
A86ZeO3PCBkyY9fl/qt+l46o7j4LPBxr7Yv8NE5GynhQwXcCTFdz5DfEEgZM891mA1V9qTUE3hTQ
9NAfZWpfhIyDcx5a9v1gUvOSO37zoOJkxZtJiLQduR+A7l9xgGgMeTC0Y6ZXIS/S3ahPS7TV5iBN
7rKRxzs/5iliGQWjQ+bdTKtsFxJewP3LKi12CgCzP+ggIz9lXX+kYWAduKJCP47cOwLg1Hdb0cjY
VBb8Vg7cJARIXiug1GJK1S6qd+rmtcuB1S4o3hBdZLshLggrGfSuRAwf6K5Mi0JxyBD0s3Dgpvij
3O32zZGdn0vK8CBUkCkohnzBE2je9HeBRdgN3wrumWMNShP+y7Tc6yUJxuUu+0Tpa8n6jSVJYhic
/ThV0/0UjN8jJqt0+leWvDJpP8PnRoWcjf528Mxw/sw8cu0NUL72u/HZmkCqj0zjLaOqiEIPyIpG
jMVO7IRrwpaztZKER70VDcLqu/mfToK5src/0sd+QE8wJo3Ce0YeFHs2Ld6KwyuOvJYRNBk5az5p
Fqje2GJaTcf58VZ4p/+kQNPJSWNz4EP2C8Sye/LouPoQgII9Y5IaolRURFOy9ivl+efKa8qaoD7f
6/U3c0J79GrBvH0q8b/sls5hZWUUH4USxnYmSEQDviZYtzsDXNVfbNjEycVCLHEXI13lDhNB7+6H
q92UcsblV1+kLpQcaliiPmLVuPgKszQ2I6FtVE2hoXjAOaE7u4aIyI6ytQakqN7nLfyaP6z+FPvn
4iEgWQYCyKYduhDKcCQT+wgj2LEz/XZs1KcdBv2V4T+Sy7XCDtHOMY/PRR77/oZCuyfHebeF9Djr
+jh3IxozK5b0NKaH2UPSkvkRtC+qof0qtu0RaH6h7lCu3LNand3YroxOrMIfpBPW2f79V5GIMnoo
Wr+YX6HPhGs+yDyMA0C4qelqxqOsDmqzltUPlmfdA4sdRpBhVvvWbVrJaK+bmEdULqzNLyirSqbT
0uKZzl3etlSFyvnCQRBzngs209eQ/JluF5OwZST6cLQrOZwJt3yn/FagJrNS/Q+/srPrJLeJsUjn
kT6gIueXJ3EO7dtcXez2MnJYVI+0fwUEqcSIjrV6TugpnFshO/sJKSWj3PCLoZ8CKb5KjBibxLrh
T0+xfAL/Ph9lc1keDw33XwXbUniCfMz25VGVliKKq0dDMQb9maZvW03j0E/d1RlyA6MbAz6PURow
KJzVzbjUaIIpTYcTn7J2aTG2HE2op80i8bPZKTRDSLhrwQyBSfHW1DQia0C0p5Wfw/cCSKvi7/re
9qdiYKPObgpeIO7FUZCluVcrJ8H5qONc4fpSZrkqhzQYFfM4TNyWZSFuR9MxmZSdZe5Jdrx0SGO6
+asRd2b8mXW19sWFAw0TQUapVM2fkHWBrvxMb6V+xEFuVEjhVGdrPqHcSv+HXNNf4CuhrBLBa+/S
SZwZy2YbbsjdcZvKFuJM/mAvObuc3vd04PlnHU9phu/gW7geVH6Scg/SmUhjcFI6KMwyiS/EC4LC
SRmJ2CRiEjx11/r2Q+AJmtBB1OaBkli1KoRn4Gi0TnC5LzqGGABGyBGK2j1IE+5W2Jb+VaqwynqA
vdoCdA84pPiKr3fFsA5s+7q2T6DSCDY2FQDC54EjuZE4jNOJXDRRTR6RyZoH6mEA7LxjD5s5e77F
975JHOOvbdA5mEQiptk4/Ezc6H4qv1MAeYKQEv2w1uRnphqArUi507z8UWQ48D0yGNb4VOMTpjav
r84v8PHjtO7OnKeImH9mPa2g/Pc3XIxrYKaeNDObi96089tVYy3LlQ6Zp/K5q4lbjRHrVLXJ6sXt
hE3xY/vKpdtf8Ob1i8rtROJSYIwfLCBXIbahU3dl6R36WuinEM3jO3omNNoW78oHzm3XTUsgnp/0
nWBQ24ZWzeW/38bdWmYyaHU3Zj1WA/03T1Q6pMd6dRf+NVsSq66tn+W7IF2SiXuDE2PoSTf5JHPL
/+NQt+9EA4QCE+Mt52yzl3HwjOdM/hxDAGIP1osZr1c53hj6s/CCfFsW9OLW8einWb8z9SGppCUo
i525WYhRh3ZNsehnJS/Fd0p9754OBBu8jR3K8S6jX/Pm3DyJlSNKSgS+HnmS1DMKtzXW9HCXgCIt
yCm7DZ6sauLfwCFz6NOc1tZg0483y4IvQcewvE67gZR6oDnSe3ErbLzvSau+kqCXIrDgIVlgu4aD
zMqAOJBRFgdmTyrhcM6VogEJOqVX3Upki5uAps+QCzeLM5UPPWjn6IQcpoTP0luDVs4RhU1pcdL+
hgoq5gHEfSuCS8KnMRHxHdzho2s3SoIWlyNA6sB1kZjqxT85T3IfYC5AW2UfFDhzRpEYIE6xgwYN
OCLDZYr3ctZSl6WUeTbo0eZoVthHjAeak9UKwsnJ4+4A2eUg6f+p94aMMFtq8rKgpyU+xaGiItxd
/EepVjrZaliIj7gUZZCaXad+MF2MyAoWCQQVIE948kQ9kZxCi6OByYHtCpnC9SM8GzwKf7B0QI6v
WQgTTPUw1447w8DQjDpQmA6zqzKUyUe+OrHGlpeTG6vp9fJsAkOuiqa+XuNQ3XdV4k3DhDTbhxG5
EG0p661mbCytrJReq2iqbojHixhGW61OdyNPT/KU4vEIYPk0onzOyj8Rq2ycZvqDlRuEgqZI/Enn
EJqEu9FQSo9eDsI7ap+bKx/0jrddgstSMWFdlj7UccBuGGAb/dpNL/K3VBfb4e+J/Gw4lzI8BaZq
JOF+Hl2Jsx6u035z4DfJH/A0zdMlKJACh1A1q3RJ0KRvVmABrM3mDECwD44SJhtfcGechMgxxCE5
F4d26ZHPjPoY3UoxUU4ViKSeWddVa8ADlYCUl02cMqa4XpENKG3PAB7zeWmmYrk5fPlQ3lmDbeYO
vV6P6V7+swJmWIMJDoNUaNmjJQ1W0DDmTy/4QeWzx/KTSRuEghDl9VgvLDpen4IsTvM769FC7Gz5
21e/3BbUIievhYQkFs22WHF7yvFone4EArkr2qp8hXaTyWCxpgqWCkZnxuh+s1gMK/Y2745wnBib
0GmD0op+RPPP9cy3w2+KqSmM2ZogXADYJd5hBSjxmFWmT3NXA82m06XJxJjCxZlgRe9IvjTllaIp
tTCSDSTh9gtmkKpiFj6mI4iBZSyKK+Q0RjrQJUqU8cXqttR38EzgZIqCAXDk7FrQjHqNCSldNTSf
P8aZ1ttG5SILcKyUSwZAwqOK25RiyC+5AeetgoTXUIOkBDSjFUAxqeEIkdBv/kwLha1DcLBzeD9J
T7b+ehzpPMRIDHy7thd3VkmNqQ375DK3esZyWKcTLh+RABNhrb6iFN7LTcny6yg1uMaRvjKiVjti
GpSBfXjwc1MsO8eafHKIegeffugzd4v0lGdQ425ilMzcBkx/9/m6xIoLpVH0/UKXyrVQGpVmHvRw
xz4SDZ17N0sYPUSE/FKfK+LqGE4LXV0T7U/30dX4gMN1ReFg9quhEDTkz32g1fan/NkdgyWzB7YK
SJMVJfcjqbUyeWVcdbeIyMCaZV4bdgUc4k0mjn5QeWZWTgKtepZTNF2h1e+2ZdGCZfd+PBtauPg+
w+1Bx9qN9lzcbTm1var/USR7G7IroEMMU8JtPHDX8mZGQxYETnhI3l+OYYHQ+5dVzd5NtUIDQRk9
PS14D543YLyH0m+p41bvC2pDz0yBJLps6A4SXRO4wI6biI3gxyHRWWUPlk4lCN7l8nV8Z1yPDOgj
iQhZ9ZSlDZoT6/s82Ki5P0seY8vsFziiwR0L1iO7wxXoPRfmbcreVhqsEQfdpsf7W2zT/o8NDrWL
FVFsvVZi1Krwr9Br7a/z+hN61cJUbodWT7B+jOCV7v6vR2ysZDySX0xG3SjynkWKlYx8eUBOc3XD
shpjlz02TEKv4KEmWbw6T25+9kG75ebdK/Rt3JSjd5AAaaqg2ecNQn8pXtTGXyKrZGktEdryG8zC
Rn+gNTYWAPli1Ed8rJPoNruMJatJx/XmFJ0fbQKhv4h86Znkq0XdZRa2JsP7IYtmEh+5qxScC3AI
QWFYWP0+wvGdhTw56AFF5gnxIONILL94vvVc5R4wUYx/TsLa3WtZbOZheZkYnmH5I18BgOKt45cL
nfbh0vrsvIvEFRaYMx/t5oCcZTzgopkc/gZU+ozwbElp47QBrkBb7jbUXVJxfRQDFo8kxZimEA7n
gIZywWt1YxGXS8e1uH7bPg1Tiu5LJ26h5Vv4ZCLghQcmpkS/upStH5VPbkGrkwfcsWf9igDfPbhN
9q8a5LE3Gi7+Yan6e9ZRlDPFyfttiCYEiHAm3fRACrIB0Ek9fypvtjwsAeSCO97+oDESoCTUyRD2
m0ZHyqKvnaEq8j+XrrBliO5do0vHwfQSYY4/5quafyJlgU0FwtiJaAIFgzR9g83yypyGIE0dujWy
0f94cyChTfkSUdE5vG0LeIRm3OPvB4qiPHgBGBetZnEduSQ3drYW4ouf+tCp0cwyxmRSnE3wZ0KK
/um1QkPXUgskEzoeLfK/N5q88Ix/qM7ZOcg4sUW6YbJmaG99EBQoc8kujkoJDItmmuw9eIQhNKtg
iD2zelTNQQrvCywxEiSZxcI3a86BRL8A31mh1Awicv+s1B+ahCWw0i/0N6JumwWb1amPuclCigCh
wElmzajfvXgzUf9dXyLAVTd2taSj9uznHrakqf0Xv8Lmn+Becs/u81lO+2CCO67CUnOJFhiWvXOv
g0x25BSrc6YSXxI9+7oHKZoJgrXj4V6LFbEWYLZERqpNpgT4FoDbtlJty6QnxW9GPyPFVylY4gKe
tyb6qsGfQkkg+a587lwHhztwxpz83MVDLrJXdcylSTSCOzUTRjEN6JcS9SPX65D5AzC+3hONzQwo
VxpdN6m7noNZVBZdad4qbkk4XsqOBraInTCXLp899SM6yTdu9yjhPO9RjbHAWXG2cXpDe+uddeIc
UDk8ebnqPhvcfRCAAqqfDjjyvg0LmUq6vdKAHo0LMGkWA6fpCrCTQ3QjJaEO5D1NVjVWoL/bY8hO
Iu7pKq/vQR50wfyuImCLXbwwBWSKqjraBdwdbLNwfbAxVdDmsY1gEck1Ldec+cxwY+xmvccBvd7N
IIN5mOPj/d8IvrQ1gEjtrpcEjIWNsojnZfMXz0kQZUKPNAmOR/sM6b/avYtxY03X7ASYhsl4fyTx
8KQQfLEBylUuCKAeZsuTltSwgb/ILBOHMdpfslN8dENIL8Z5cjrFAaSfvEPh5OajIoZMFtqrgsnU
5CmVCoyHxiZAeFWPQmbV0doTEE6hS/JAvckChIJjHUrrntfqKVG8oapdpOB10hRBAvbIL5ONxtzc
nzevtExonSB6YAQRLGVIO7+mhFLcrvidC68edPfhL+nvpqLtNF5qcAm2CyfbCgbAHKBFQja9H9qW
ici963Ll0/NJFHYlAktfWlQLLKuJmQuaFWONFmhn0bOCs1ftwTl91kEfWii4FZ/BY7c8mwmND4dE
Yq1eOQ+/w9eRaHk1DGxmvcdEoLNQYIVTr1Q+2T+H33PcA5rmkr5rARx/logY3gcwq37ii6mXZGdX
O1YgWPr6jVbKws2ObQPip8ohCkjR1LpF+hYRa7p9ybFvZQTO28sh2HTJOaDknw+8qT2xXG4eKHgd
07nVf7oWo6dZGRvfe6fDaSusg+B156w1rUcLYrgUpd7SaYrVEna6fRAX5RlK9l1QMrDqTPOGg1UP
odtNCGE03tUTO0O9MXjPrE8tP6yHwEsf2ai4IoA011/0R+UvNTJplVcnR6JrlG2cttgCpheyJ/39
L3waqvnGFkg0HSKtMvKhM3hJtt5k9mE5MZjIQ9dwre8D0LJi/A0nsfLYKjG6CWH8TwzlMRvL8Ct4
X02xk+OnHGlhWSn1lwl+3SmaoEx1nIIanzsvRqhVwI5iaGh2yZfs0bgSFc/yGf6A3Sfvhrpm93L+
LXL5CUcJz0pze4SYKNTon8r+Oi/tSBkW9KywnlcMbtMKrRMkgrzm2Oc8F5MhSuG/3m8/aGbZ+XMa
hrPVvJtlreAHnTo5fJN+7aMZ3zMqzzwXy7QKy7WQoqAY8K5eAdDKYgKMrM/m05DHPTX5AxJvYFGL
8epmtvP2MwmlNRqtvUSB6/94lb5Bczce9sbMoIpRG6gUmou4i4fGw0qD/cdO3vM4kqLVppEHQfRX
3ELhJZNNZJw02SpNOjII/cB7Srsgc55EaeFlaWE0K9h6Gtu4goY7lUtlr9X/YFNc1FzF9OavgZzs
b9CqA5RzkJswc/AHlRS6rzb5SmjSOjkZ3T7egaBYim1YfMQaM+WtBqKd+Amjk22Z726FxzEWVkSD
oU+j7tp07JGH+gD3VfJJrLYz31Rzz/1P6tsZhl/h2bfaIUxa4G1F1xa6KM9vZDcxvwSZx+SXUk75
W2Qk9L+CBL/AzGsx+sQeCUEGOsHJRSUKQUl9AHdkfRp+3yisFsppoVPQGsoMo6/7LZA+r4zynWqI
0uZOFVuEMpkXTQ+/1NnCFogyRDL4rmzJbAWAcatjMC6FZLxTwyIDAt/Mdgj3Q/tUbPyZvMj4wDEH
g6xJbxW+LtvfUEornn4L/b/VVrNY+7RqGhhCQoNw3+lw3h8WIHV82bO0dVGluEqYZgaEChQCpnAY
jVcfCxBXvH66Fvq+k8M2ePcXHrVpMhgT57GLAInzuexO0+G1wlP9E/VhQaZbr5gmyP/0vj/Jy1w2
oxjisI0TjFKDW5XtXb31vmGWERxfZmdVFxDyX/P7yNuBOB2RrHIxQVLZDwCFBBs1dK4HPzxE3DHr
Yq2DsSLxulQS85zCK3vXAOu0rKaPODjt67/BHfZJQmWkr1CQJP+TYpnHO3Gt9FuSvSYT16aksLKQ
opiI9NCAmI2zPLRaoF8OTePqJdsvZuo7LwxjnMjBd5T1Lz0TzCKk6bJ0SEmeIBS8CdGaXuOYriIO
xXamUXMSpMCvyz0iyh7bYIuTETXEhGUjEfpiSE4ku6LYt+1ega1D3REzs/M2TrLDd5HSzmptmHYm
/0eEzjRKCorxjzaS0GMx/3PKU3VdhR958yA7Huhet+hPT5mUKR5n3B7m01NT7COv8jgD174yoHxv
BcvLkpHnmn75xPnIAqoeQKi/is+W6lLx8t6FrteXnbbYJ7VdapHcUw7QTQFNbEFl87xSl0rHGzHI
nYjYq2h+UJ8eavqqs3taIjZTqzXkZcjODcuRZXTmV0OLCg8vJoDVJr+p3QYtCjHvv4h+8VH+muBo
RrgxgKkaQw8qu6MiK6uN0qiMIsKf0kWo5FmCfXOs8fWiZ4LkPky4mq2Ht4cXN3DoaK5Qo/yEF544
vrruePuOXuc8tbdoc2Mx/Chdaf/AtIbr1uySjUM1qTby0llyJyNyoV+VeG4Hkt+lZjhpw2vMpoST
h+sliwkXNTOyvLeklzRwIL9avwYTY15GHRKdTUx7TevUCT7qYYaYUx/qzLKKRulCggNnr9tb5sa2
wY/qKr/AM/AMRgitqnhu4FGEWfpoPY5/5fcJAtUsY+Uv9yMJuLwRpmqxuFpN3wMYOexF46OhPc1Z
4zVF8bChI5FQtiVG3QsS7z1UW6prr1cHazL2rJalGqtxF7WVp3aJv249tCCEQCOz5sUiw3+1++GK
vXFVKhPPnqWphZmrNwy732KkH5Spys9gTJjXPebfjV7suYNB8IAjwSQrosdqOqxfS7Zm7hT/CLxP
smopy0sqkAGpy71deK2LuEI0THaepk2oCAWd6uuPZI305eXoRUQ4w5KoMqAeUq5XIm63yEbmi9Lw
HeaMwKMDUpkMmnSwUFSDZ76toGl+LFGQIVJDeO8jZjf997WMsvpdAKdIq6KaqJGtwX82vl22NdIp
KZJ2zetOMzFWzw332pLEu17dTwrBq2kPzIN2vlw+ms/bD/J/C0OteuuqjTwyesl1ewvAeevAogVF
dUT2BoSPavk8Xrace/QLxMMnLkvfG4ThCLYe4c+PuGdB0K82K4S4aPzsX4fAGu9UwAY+bgoSFX72
e0YjSz9+u9gFPdZ438AFZDxZyXYCyUQAdLI1GEJVHELb5MFSlT+Bsq2frMrQjTrUYMk5CrMENhbV
M/BihQF+RtiM1kjF3aj/4JyQW4ap1iYFMqtxu7+feoHJxRqMrUr6kwm3LxWwHDoc6T9BYIB35g/n
EHTGxhOEgh1kMMehFzhbX7QtdOaTBXLKu6KEhe8sSzBrxWp4vep+2KdrWGHZVj7n6kenhVAIDk6H
Vi1BPt4An9Er2eIlh/iYGfpZNesQsZMapEHh8lvh6RyxXHGrYc5IhBy90XrqKKWdP2L1EMmGGreD
vOwV6IiPpK1rn68rdMJRdwtpngkGj0PDVypaIEo2mLSKd6B755VUpOaHxVa/y6BxSfkXLaosm7jc
gO2eafu/51p0cO4plugLZl1t1ZbEJi29ChqyrF3pTFqWLFtaUlBYmpnuMMRzT/C6cQ/n7WY7PO5a
GpNYt7ybHMCUF62Cbw4e0LlrgQ5Qr5L39sCuxROUw21Bnk2b94oKi1aOtg7GjAwb87U220eNeWBz
eE1xrPfHQIvBLyXiB0FvwxuBCETDS1kknF7J0LoDmDmkBfFuL8GyfMLqIJZ3gGEN03w50o9nLhhk
V98WXiUhIwxQUpjwarVuoo4785N6fvi0dtydFuTRPb9tpec4pTlLkPD51Apz+UOadrYT+eusfjVM
X5wlfgjJasmnulcCm2OaCve3ccRc5hWrFoOrFtMEnwc6iqHnbhJswBSVlPAY9mXAH8TZV81DlYH4
vA20vSMOeZunQULay1IOJStl2UEXSazZNUtNfStwZgIaWicSEgxedPOkbRwQiwN5TF+e4CcQhku9
PjO+AxRw/5Gs99s2XKZk9knUTNHQ+6gw/plc64SkUM2EHTGD+kud2RbMEo12f2e7AOd0+3WGyeL8
3+X5dPF1nTriHhHmXBj+bSj0fnEeO6ddhc5cBCrHx+M3/tgoC2yyxmnkkt6JEuXb0UVRXQSwMBEM
al4hxwz2LAO0z3VkDc4sCDXJQQ0lTpcJKHB4+VVIMQDZahvNXlPNHjD4qKzgyZTjJy4NnIhvl6do
qBdx6LHQWpqsxtWN4GOe5G/ljk+UkROJcoc1Ns2UXJhZd7zyeqaCPfcg+ssbYU/ODEOOKma1/GvD
2gtXJX2oIqJ/KIMKslazZRVHP7EWrOyzw+An2vwVFwmYK9Atbn/2vy0w9py+3hkiLS52Xu+Ol/1y
ogAbzeBmM+Kdgdld5/H2LbVbnILn7YIm9Xdmqjl0N1jcsAMiaDLaSITt9+HY0jb7lBy7qDgAgLvq
FHSF0lJglyiaio4S0Y6sHcDVlBB8pZFglXYB2ABdSfYjRd2u3B8s8rj4hbHOhEOW/YNPTp+pKQBd
lcKAqwND0Nm9CbY7tvgD3TZRpE9sfLLwNtr264Fa4h1S+JUOM8cFKZUotgHjfloGe1/U6zHI5ozY
Fe22yMkGeZHbrEwSq40tVtIWgHeUAJ74OgTD1TDSNXoXctjVU2OZbcLcVAFZKwq4wW+z9v/kR6gn
a2FuLNUJ0FxWqLWWiYi2uqZlWVw6MAS0aNjMydpderyF3NbdptYMIYymrKCcNSoMIRpVtwmwTVW8
vru0Frv1vWFF5EXFZV303HwHSxAFy5ShLQPb9qC0yKzWWo1eyIshuDihp1ku24m0/h9jlc19Heq8
BbW1YJEa+nLNQrB0VU9wqhFz+Fmy8535ha45esz57SwwlBczXgHiTUpxs74Ybs8qVlDPXntqTHgZ
E5YgiBAzMWwR6i6wXhM/04wc63SNHFBPQE1/THltJ8zJRi1TVnbh3C5IsoywcA9SbKmSWDCOvQhu
RLeUkiKMfkqDkbByp5HTTwgiY0sWnYjgS9MqkayZ1eSw2oDQ6XA4W2XA/9yVhfOBwSgSwitdBUMc
0OEm8s8HABQ/DF38t4KYmgzH0cgaEy/FbxTDRcyUszuAQDgdG3M7zwnLHYSGQ298D69KvOcvSV/h
Sq2LeMCtbYyEGYgTaPY8o/1CsR038RWMbWgf+a9plLqztS5wjSneaNnAdaLPejw9c0AO5tsgaXQF
fZdi74fZkPxWfQvxaCo/oWD4wyRzlCvzGZQxyIFxOJ2F/Nb/1goBPDneFbXaG8NHI3x6Svo6Ub9B
4wN1IXWIK2WXDeCJiaBA6uVc+EqhUorLZP/6fNV9XEYCw6HPXPPrAHfNFz7g9khlgyZj6ra7O43a
5ruOXVmIZIpjbK1RJBXKBu4Psm6nJK7WHd8aaYCucspbbYmQPIh7ZzYbyqkfJwSM5SaT288XXd4A
+BT96Z3GJOMx/4Qw+a445tgqPKaen5WGQZQXzdJhvf9ldvNO37z/z2S5oFJL3o/+8E7697fxrwTw
uXVye8w3u6xZMjTEKMipRcFcUAmCYGpevcmwReS3V28JP0FfiXNqk0WfDshnp9bV5wwFX/DIi3sv
cNMGjbyjPMPuTlwSBNCMpIpnlXyf/sXQhGd3Aj5T7L6c5j4QqZbrksYtkTOVIcZ1xFwuidwpfQIL
iEoDkeybK8hALPvpTratRt4GR1M0Dn3awyalQg2L+CleGB4KD2paPvgDF+w+uQoshCrdYIWmyjqp
GYGgoi48lYBKDQL5BVeRVFXYGwJ+Q1ofYyN3xieW8Zcd/C/4Px6y4rf4c12yPnW1ceVL2cQxUldB
1PZKU3NSIH6YMbxgMISCeNwb9GJPNYhVTwVUairEqoKcHdCwR1k+WHMRmAzz5tt01+wEAb3swpnl
ki6SpHHR2cL9dXoPWtGC8wufLEmYrY8S0vy7p4pm7P8zg/KtN6VdX4pG9DRjPwFvgWi4X4Eftr7i
IychQ1MxXBLeqLvuO2+2lU5KBV+tV3BmXZHj3xKty/Pics1a2ZxggcfgvT7/CS1zL0P7xY8lY6b/
9VrDK0MzxvAjPST5eO6cWjJFnxaKtNEIWq9xUe0HJD/ADBg+ODaZjeufrDBvfiguqDlMY2G/lfRy
gHuH54pF8+t9l/KNaUVpUp6SSIDeY+b0EvJd3lnQeaxdmzyVME2wK2E4u9f0R9QghD3oRJHgXFBx
wP/TUyZSKZZhFvb+07CW3o8P+rQdJFx2EhaTC3TamvyV1MpTDPPn90OnDMZgfcmy6DI+oBEC8/ol
lOYVSKQizvCVrtixxvLTbziyBYICC7xLpOSvhSqkONttG+YwuOl5070wJa2MGnZCOGEE3wVNh5ac
4BfQnQPWiZcdMtwjgRG2Ftxc1zS0Rru6Zd2/CWTYX36vdDNb2uuVVgZiD85ZwHRmklq0yquu4hjZ
sJG2UvbRZUbz0alEEz4AtUicyy7mFz0/Y9OAcOcfzuRPTYYvzaD0jfnui96uzMRj+dH3o9uOZ9Bo
UGdNLfIvY9HP4ndHgGxPmD7rvL/YfVvYosP7LpbS5t2C4E70Gw7TR9QlMITsD5iLknUiB4e0qcs6
tetfbIFBYlsG4Jk+Hx+bWAF449vVteJON9brtT0Dh+wz3xnca9wR2Zv2rvtB6MMrAUgBQbrRkZJN
na1aySDpcJdjQT9tR/FZEYXUEe79CjJ2WAsHWmELRLCFGtjmoHISv3qDORnFLRM3C20ZnJLTCmq5
8E74nQlqUH/hua70c41z41t9ET3PqqZZ5dxrhfxC0yc35j7HQ+3osd4pMIYC41Yx8Vyv7BNvF9Jc
gBvaCk8raeHG5maRebyTxHLSS4UH4f5X7G2H8bZAZQNFMrqqdPcZCv+/E+kADE++HUP1I6Zi1faf
5hmoY1uzODO9Tla4C/1YjKNG+lgGCdqQZZ8Dfjk9ZIL0Lt/51ORt03fNM9DO07KUjgjVZAyY/9Fs
eKIpU+vYoy/LB4oy/pP4QEEHa/N87j2EB9IdtUpuKXDh60NYLDPrXyF7q3H0wY6gl8Ofx5092oft
JKX8TC0MjJvPGvrhASuJs7ArokN70B9XvPzqaF5ikzr4wy7D7lB0Nd1VOOc2X2jpJBFfw57ldH+z
HyX/S/1owZu8P19r92YZopM5psfq2uhPDfIJ8M1XGxGvNoF2XFCldbzkdOJnz77qB3+iySNLLK1a
PEyfR768w7nUm5kiaOiWuVSfUGi8z7PlLN4QDpXjodOJJh8zrSFQJfGUB//LDppdDpFwv+XLH0zg
hWn2RUi7MQEluKWIclZFjsBs7rVAztUQB7XJq4cy0AqX6uMArDNmlREndSfSM1/Xv5233HzjUEB3
fDMRwzQEBG5vDaF+ZB7lwqwHmOI1llw8TyT9KlDnNu5s8XZaXRXZevGbz59TcHsL2DuEPHXUXTjq
LwewM4e3Gc2zX4iZPFeq2psNigbGjv3pyQ4IgJh8cfSSRTU0glPN/A0z+pTIke9ol850RKq/WNhJ
BLB3W3H7MO5WoTdQPsUv5DaW4f3Fvhh8IVOmIZqgZLnStmh4m8oCHnQelUQojG36WP1l4jEaPX2p
1NGLpVC7HjP61hhtvSkIPbpJUOsWFC8sC21aycJsBYtgUG4c+J7OdNU8r4cJIEERYKMnU+PSqcn1
ENIbnySHvneZDrWnMBiD2M45GI5YyjpQ9/5FwF9R91NTjlbWzV0L6QgsoZVQKAxF8Ii8BK7zN/1r
cNEXiddVnm0gOpsa0hd7SyIUn9Sw2SFOwBH/b5NPFp7z5xtUWCSbox/Sg+jbuwKI9N+ZWoAKVLXZ
pFl2Fa9mlSq8a9c+f6ZbAbDibeO3WtuAj9nSukE/9malKCQV3PRbMrknJHkJEC+WLbpZWTW202xw
vQfQ0FnBw/eK+GVqUuUZDW51sD3+CkEYV5Jn7UCLD0jpHx90uF5mLxuO2tqkaIzxJkfcyozr4gjY
g46RC6wQGrbjCxMxiSvjsQ4pO4CgdeVLiVginvWUgJ0YKOVaxn16fiS/gwyON7il6h4IVihoBbYK
RKzE4CfoVxE4E2TNRRjqBVKQto/Tda31UZC7CrvdwgZeyhy5eP+982OjLh+2oiBii5Y+FLRClzsM
y+dtHY/Yk9UAWC6djDfwIflfIVflaOVd4b44hjZi5gPH7KzL423gK/qWr9POa7SQWF+945fI3dEX
6t1klNCuY0bpmi6H4i/0mGZ+XBjRMp9wpJyvLopJ2TQD4G7tD274SBZm6hh3xtZNTHZmXCoZF945
V7FzHyhNPeqa3k6BnccMtRYeQAuWdocBD0Ym6biVrZIAEQB8jO/mKX8l11zqi61GmJ0N7wg0VR1P
812iqQyB2BnhPDNuQ0mAAvHkxIs5QZLmOk6g8TWeLiO0KgqNFbhTss1xFdQfopYxJNLv2pxFsBaH
ohcFHt/prFIvqI9kKeaHHyqhra2voajLN79fn7dCNi0rhjNgqWX4fadKxYKqFDNR43ovkRnJPtX6
rr4JOEHPH5TByYpgoh4iw23qeYGaoJ2c5Pna4GUE0AJ3DkxvUEWdnnqMBXQIfwDYTY8PIeL13toC
YvcDBXXWGUNqbae0goYSP4siJW4BPGdVEOrbpikGxL0PHWUKPUeEGedp4xqqoQgCbGl3WVsb8uEx
ElB+qwUzwKp7TfSsn2uAtMshEWe/zhZ49IZIQGStm0uGh73LdbKmEVjOQv8hgbL6C6K8THL5MkEI
Vad4hMt5Sdvvq2Q9yvSA6BunW4JzqrFUYRmRjQBpkZ2vY38WenXV8csZ3Zw93F6Qg1hOzHNy0p6A
g2TtC/QdLAnHBsz07UCLO5LuURFF6PU4zq9pnBg1Jl4RfC4PLi6YUMq0M4O3OQW8ERabP//oFu1d
pEv8G9ukXWWOlUBVav3TD47mMZ0aYZW9mc5HYo0AZpHs5YpmNmuTJlPS01EYtdAFV213cloWGgAw
T+SQIvZVvZnwH2aNC7zoIq2VulHx2DCIuQi1Tkgr+mVqTjBvanUVN4SNwBuXCvEo2YtRmHe1njiz
6pvxQ/0E/QMkhY62YWjGO7cLa4G5pcR/vmklsk2IRx7CKDfLRFfFGodTQJ845zOnXCx3uw1jcGYb
hN7QLXTPlIINoNdA5VGG/sxXneaTSk5qFowvPj42evB/SeDdYOA9hWYyDjybpv6bPFiTzvlgAbAQ
b9AzXpmclErz7B+/SaHfWDGyrlZVx3/OKYSTxPb/+wIcIqK8K2aNQhDF7CB7lE+ArDRXrjhu0smS
/XUaRhAVeZeRt1mPDp8SGRzEVfnxQwsHm/w5OjniI4jIhPRSo+YA8KFl08ewrD3GR/LtlI/+6EUN
akGduJklZgqy/y0CfGfN1ANHNgQ11lvvrsCN/nbPz4buPdXz/Cyw28BweUP5CYnocTWv3vtCWrXi
Kfrqfmreuwd//OtXcIYQL6NkgyA7Mdi4r9knU1xorRVKcToV1mQLJ3h5IF/VmsXNpjDxxJKJbQHY
CQ9rKR5RE+MSYnjOzpAK7sKWokxxGZ0A/YF1wHRzXw4DfUy9GuAGulvkPx7B4+E/weFl1xmrPb4t
R02vAzGGJUeBRRJ7G+Ty4vv3FJrTmBPxbCaxt4pscvtExYr6NHNa5eCcEqCqxZ1aVPuvQPDezH10
UCWFqRGISc9Ln1Bh/Ekqjip6SaJ4gO385P/qA7VcCpVgwVb30aR7CVXCms8g6irHSPk/owrCy5ch
XFWPq9NRxZ06H38Y9CT/dQn47G7E0uJoucOT9PLFETj1zrXgP6+1q0gb80NeSyWAHtIGTcd3icQ6
HS1mk8/0Vqwb7oHsBnzaaCq6PxEfuILzpWzncxgTCoHzPKJZ3ZQuEsOh2r1qcCqdTfLfRhZPXg6a
hevfjuM1NczGS84x94KvP6+MiqDvtvg58OPxpHGMXpjKi/G+Q629hm6ribU4ns/7iBuaFQtzPMk3
upzLvEOZVtwqxhSCvXTx5vMfbbYwWdIbJ2ewt94nSDnN3cvESXbHs00NfT+tf4WmtSTFt32XqK4i
gg7xO8u5/WySaB0G6lwJpgF/h0sCbN0W2qgZmAqMIhSrbdFXwR6PB3Y7S/iIBzfPNu2WyinE61mm
JcglecLhE0sVIa18HUyI1O5nG2wfnmadRzotU9PHakY/jS/CbC7hCi2Ca+UZ1A7Vnue/eIlbT3AW
0oBr0+AeKNFvgc0EZHmAYyOp0HiLX044hE9SJAZSwciqPeC+TEzWZ7UkSsp/qfP+esot/gFLWhWF
yiuTj5JNj6BRb8aOE2R/FUbB8AIpA7qgHf9JOlSIelir5b/++8eZKVBqlSc69jPBgMtC+ZAim/PP
UOKctI/1OzGP5yoPdVfZsMJP7GvesVTfqROL7Z5GtvsFzmsXkztASCvaRxBQUxcuL5Cu9g7/STLU
gKu1jsrp98eCYHTcS39TrjyaxVL2BWPWSEm3lcmqqiRERf09870V4rag+ohwbk3TbWCiOhPYvBAc
JWPLsGWBzAUcESvu6TUmPWYxWLOjOKO6RwRpz8yDn9INOAp1BRHX6FGndL4hmiiSBUnJTiAX4poQ
joDiQ1vTuhZAP430ig1bWjoWsoV6wuwmsJCaXcSetwFQxXizA0wSFnjW36As7Ar0QAnxFh1EvTqo
hw2UxyXVBKYmDWXVQThlxD3SoU/Ms6LVg0J+taPS+iX6S9yU7JNA0hLgkee1QExiIM0zGMF9lQVj
N/r+SEx0c02hf1+zk33G5F+mN7pDBZQgiaHvGeBpDYk8miTSXYkGLbfKRhTIrC7Hl05wKYIGY/Tt
mJT5qwNVmHIppjSjEMeiu275kjPKcnSYDqyjjtu71t1ltyf101UlZ0/pBaGFmQ9MRQtSOuxmvLs8
ZDUP3AorAoDRaRaiVWhMHyW44IwHQYKqJhYTUm2IzJFHuKtcPA1rZ5S/VuQTaAEJ1A8CWbk7hKx8
3QNGNMRDX7jGCWwe1IQOjaKvGwda3AzTrzBgDPu9Linhwp01a2iMw54V9ikekCZilFYxcbzE/qUE
0rjJUA5wX3C1xPcrG92l5sIXU58kT9zl8/ZbDbgsY5O+EyEcQB5tbyX7bf90Ts9P67Iq30V+/Oq6
I4z7DdbTYILJ0jnDQhT32Wor/rktknTzDzZMjzbKGzPxjPpYoCVU+qXFbtrGo7lQQDZXHlJ3rf/T
noSbaWAT72GkzfIzHVSqpKOc1bYJwM/Hct0rPZphKOtmp5w2xY3lVxKGjGFLZ72GhGraZkc/2HYv
NDbUP7LXlA/8hF0siuvMhd29SxEWLuyrEk2xNLCwpPE/6YVCqrQeh7KqhpVK3o4Gff48hJG0afN7
AE+OHNYnffLs02HJp8z9RrU+RDk7uS7k89OqBi0N6CMJYupydVqBDFNcPL0KmuriYQPIbXPzrKIw
h1G9xM5L4c72DmoaXfYvJj76qxNeUdC9QrsasJ4wvCmoMauMW6NOPXvU/NgEvV4NQCqYZd/m/vGd
1tjj6R+o7nb4FT47ClKJ+2ZPvfpPzpP6d0ypoUI0HNTmZ/Qljm8Ceg423ClvenrDdlDxTXs1IJe+
Dr7phqoyhssg2zN+rXpnxg/UjJfe9TSnXoI00TWMHhvqoC+XNnZ6J/8c6/8M9Taxl2BYtdRev1qu
/nzN0GyqUPZtqa/GtqW0x0Wnn+0s/dcNSFG6P9OoTMyRZfkXQwaUH0kwej3s6i6+GURs7tuW2IIQ
PlQOmHpsqjOJzrKyPJwiMixqSV706rH3eYv0oFDNzCWGxnWVfmMMiXCMPDP9K9LhfhtViuZ5D0dJ
GQSfSdPDIoWHbBcnbh7YQY05YTgEIabzODFqrHZI9jWQhdA2Jql4+OQwcFyYci54q9Z1/e5u6Pof
vhnu/x5HeqnwiLLyA7sWb2OQBnFQgiLgbwIYqhm8DWRKyimGeJQo/jxOGSq4mrfR4+Btid9bYXOR
VmqM9N/f+GBECYgG3clwcPNncW/+M65MEPjAtMaVwJ4z1pND87KZbi8YhRPIB9DzmwM7k8wwesln
uN3QpUwGZeXUk/sSuB9EHJoAIBLcm4vO4WhEWXmqj+qvN4saIdhIITahUVfSDlxRFiAJKCUBkTLn
wpUFEQP8WkPy/v2FW8vlsNIbtL7behzLmrLqCfpp4/1JbrxIAZ83WdNyefMYB24o/xScgeqBIsDm
Z2PVonhhyxcH6HvIQIL8LLwqsmyO4aXF+6dGV61QqYs9e77FjFFI38rbBtDu6Yw7dxv0t+Dn+stK
DEETR118u3jIGYnucm8mZ9fVOn2kTQoOiqoUsNKTqwgIaQlL7LGzwHlU1sQfRPfoeQl5nyG82AKH
WfKT7Av0qDFmPruVIP0vNaOs8HlDctt+1s1Jf5xIv7I+n/6Y+6uvOFEiyKi9U3DfH1t5W8Jg0RUf
r6VH8glWdKdo1ZgkMjkmFCx2RBJnWSwwPTbmBjQIE49NgKmpGJpgQ99NPqws6emEovbGG1gyjw7t
bKx2bMryY1Es1KCjkcowLuiBq0bnOjgTkfofLGATzNBAEPFkLkN31equSwYAFwtgsA3vdzbCMES3
3SzEJFXgsJuw1yTdd7yDa8a/oKUIdwcI03E3DxTk42U4OmxvaaOA9otr1kvMjG6GF7/zjklhpElP
vx6ucuDwiuwKPobAUmX7Z7vZrPTdJ7/lh3jCqGBhoD32GN2q6LcJpa2S4uHciHOyP1CTLgPYXdk7
Uq5wzGwWy8u/IWM4al2Kd9uMOz0s+tCznWi5l5W3NN+Sx+5KUY6c+fEFDSZoquNhvhSRfD/r+N/D
JWVRUiJVPcyeKQOfp4Gn+4QEzGiWOOyytkiy3oNP8DpvhEx4A2TCeOizrrY44pEbb1HMUSBWUJtb
8V+GJYY6F79x+aX1xfYK+KK0Wait9sunz+A8LTTb5ZhtN9x0JL2hclk1/XxWWmzgHLzjtcKeUnLf
m2fPBtHJhYIfg3vIGxA3RLpNSG2dcAcfUMWfEM2BkEmSD7Kpa/8i1zNie9tOhTyxhKZSPlH6bz4P
7lkEvxV8wlroTqNmJF8j1pgcCSmxs4Ati+U4mghVd8GO+lysG7uiDuxQ/94fSix9EZO9fErMwfKq
Rka6IT9F68Hb9amLPdlw9SoY6x3xAgXlVl8plPOkxOHxea8S8/XAzjEXOx0RkfVS1qseOSYXv3kR
oxwBUPiG7JGvcY7G559BRc0VhV9Ycim/SEobGz4CMliHnqfipsz4jpImEKkHYQYbZR/cxGfmRSbW
CH+rcIBEuTMMgaafoNn+Fb/HdwLZKn064hTH84tmZ4NmvnodxWmTNXrnTXfMPR7TmNatel0DudGA
jdYxC2gUNdDPtEst8uTPHF3btngRMSZQQeiLJFGr5lMUIsRYPCJywf5IaobB6ikXYhGcKnYoU8Bi
YfqSaA47zMzJfmFLDDzrOuNUJF1WUKwJN0Za7Vj6uJpR9kCVBTOPL1qJjZrt+LP8Xe087ZBIqjGq
41nYpj2qRAB3gwKiplvrkmU8sZK+9TOd++toD2OI6p2P3iZRxU8FjIc+ewdyinZ+QVo00aU00of2
FAO+gqmm7ZZPj6uyXBPvpeJlcNkiNRsuSF6wAR8/yIGTSNOTgqNiwQTCzM+A/5+D+wECgCjJ4vem
Xy0BlMQp7MJV2mOfTDlkLik+eRdXb1hCwmrAFAwpucHhWwXHJaFUnLW3YCof24j7HPRZUP2k4Wfi
+vjBu6zbAtdMXanKoK+ghRISFX8N9jEOQyf27ee9CNsGuYwIPhP15pT9KRAZye451enzEW44gTDK
pvyhm+Hr32B8qsIoKh25gTPkmHsEZf9cN9eu0MIs7Dv7jaCSTAZ5XdCC7gTGXpKw1KZeERHqJ9T8
4gTdrGGjnsnJ6NJOL5PyFnD9Ft8LexsQ/72XcVZEvvh8+dijEmemLgvKLhA7XAr6It/qdgtzXAk6
stBU7QXIOMVospfER0tlNSA8LKpyWpegA46f9vvPogjCxH3Ltz9HiZ9RYZaO1Ryv++8w+yWnxIcR
78mVuzR5zYB9he0HBg8llavZliDE6n2TiNo7x2muMGodrd7xCs+zC4+FsjAv/Iqm2knINaFmAU6B
ihtweabA3ET7vopdYeVWK6thPZnHcI/nBmflWJL0an+kYHGxS83/1g6DJ8USExJYv3TD6pA6hOfx
dSYXiTQk2OoLP59agXgJ/9M9jh/nI7El4xONjl5fEVgbPOWMfTKFxBTKOPnes3vQAGZsH77Jbcj8
xYyhr7RMxefg5XDezpWh2VaqxYDxA2WKGWg4kuB07SYBSxgZBdtmB8lMEnS8KzWpU0uMoijsmXkz
Y85UvQikoqH6kOmVPSAYEe7FTeempSJtKbxdgQD1yBvoUHK0UBsK1lHe5pLRamD+kumOXnB4CMWd
lv+CgGb/nLs2J8b3qK4hXmQXKrssjAgVlZyQS/lojWhY5/w9K4s6dwIh7SF38IQQBqG+Ll4U0GBh
fk4uBXOpQC4P89gRSZ++nbGNl9a6wXORuID/FCXmLPTy1lQ/QOyftOYCKZABOuT/1fhDGsuPrG5p
0sFZJgv19XHh0ZIKI16WmhkdlDbUEHdzJ7XTirzCDwtzv6RxKIdOjvRITCI492qQLKMKAa+hk5O2
L1F6PyH/Qhux/eX/XApentcXvdz0hbNxU2hCTWC8dr2tmwnoBa5taOZzmsdkCFzmN0V67jbB18iT
ePD/fgGzRwJpYN08fKHBlo3KvYzRE59HuZDAhK9N3EQ+nOxP4l0OC8GDl3Pn0O5nR/O9Y8V2dAWo
5aZeGLUtSn0CMZoPUySIaYYJutk0abObfTNjDdagpj1sKzewJTn2yOco2OGoj4kLtRrNxxpS01ts
D4EmuANuQAbcZZxXGCJ8uwU/rg/d7R/nibd6t/pBH8Jv2lDw1G+Av8qTMXbDwI/SJxp4UzPw2Qzg
bgNpNdsdFdYxoPc27+km/w5thE/upNd43fRpZyDxNk3YNHy7C/P1dmky96opjqOjeKRlCMM8tuz3
RbXvMuBtrHOWPthfb79p5RpsiEI0IaHbl6+FpOZljV04O/7boZq4FSF+mcNgxKBe70fbMK3jqi1h
5vQH82vMrieepZCuF6ZS52BDx3v9VRhm7uQxwoQsZSpfs9gAraGI7A7DdCQJ6wjoSY5Oz+qtejhY
1741AQN5zUXy17vBDJKQOQ5/p+ejS2vJY6Eh+5OLiM2bJn3W+JYGHEL+vZVpZUcQCiE8I8XpaONg
3Xm55UOxosTq//HzTntaS/LvcxNPaTGuzBqXhY7QfpoBS90EwF6CEEMXk0eu52cGuY0t3/yZRASv
RDRqT9v/IbCuw1AVMeKOHVcRhELXDxVyVYvBpp+VBEFRvpnAj8ht/iQciE9u6oY7id06nqemBbwr
aEEjOemMYt/uMjIOM9eB6Ve1qmGwC9Dw44FppfpQXVpbo9uKRwNyePsWl+Wh0S8g2RuPLFzA2iHD
/66Fx2FpMhzpcA19uW2tOY+IE3ipKdrsgRgkDF2K11MRU5RgVSEI6bszFZpI9eObc712h7M8iZz6
m7c2x/nB1YFpYLfuJ7FoWEGILYY3QI+7gQceV6pqh4YDPNF161a3FHGJsrDv2XnZesoHK0U7qPb4
wT1SadJLGNXJc69X4FOacfr/cKrzekHhO9CxI2L9FbIYjEnAAuL2S/yhYIofnXMHd7oxBZxX5699
jE4VguHT1qF7CKF8P1o3N5kzeIl5Wuvjtgs9M4vSTM8i3FfUXFqQ9w5O1uLWwdUhfMSyhNnssp3G
ceBXC7bPmsL7RPPty+QR1cbA/1u+k958FZCkcDapL2jKxk1mBTPjb87H5H88cmYoL1hnRmDPsXv/
PiPxi757olQjGPqCWg1dKXi3me52n13lRLvQCXNSK2pC2ahAl8QuvWVkJm3YeTauR2MDgL/FFwCE
dhw3cse2k1Rr1Hc1bTcpH9qwVCU4qWf1p1AcsqGmfwmG5989MNpx1MuRKNCb/mIFi5iuGsmmra3j
kszhU5WAWS/lBVLlrg5XYpUwg5411OfJSuzRkurDh5v6vgoYCDZlD0LXLj5Z8tMocPk/g0kabfx6
P8ecNOVktDOWAcbuAx5HJ+FA1HSGEUYmWmfGYev+pSxVsm9GnNv+8B0DPOVqtNP2OR2AMgYXVL7e
fnJp7iDHabIpTcSJjnLd4dCPL46sBrG0TMbjk1Ar9EzLPqKsZSUouP2BjkLNTnYAST77Sxaq07xA
K9FREIniJbGL27I+kUJymQQ+i1mfWFp+wEfEEKK5JVJkW/kRKMav4U7IrL3j/rb0VqAKU5zWzsRo
FfXxA2KQmnb0RVSGQBcudJg2ec0uOQYcspCOhNhf7R9bKiXt/vweZ54BjLEkt6C07R6FtzKnSrSc
FVPjX1Iht2OabDRU70m2EaWzkMYNAe/dCLsMCNVJbzw1HLH0LpsF8WTQwm4ejmWesjedVwa5kd8z
DFXj2SwjCClnVqdVeKjHV+AplHvgFh26O9IJOE9gN3zsQd9vl783024O6+a+bI50b2d8tSECJb2S
ryvobf4UoD/hfnWnLgk1+6OlTxaJLpedmUG7x5/ieL09/Hv3AC3WnKjLD29olFnLik7ZKN0oLcEq
IXWnOfOmXm20y6a2bxfXz4BezaaaFMNtIs0s9/4LUOsL6rRfoC2mS2znWdH6p3H8GYsm11UY8ENi
wIzgo36Z8I5txExYw8mKJTiXHYa+F6yGSQsmQj3CAYIds6aT/v4iNdcmSbkUMTpnjKWCSMl6LW/e
Z31M24YjkFKRzEAMDbsSpABftp9sbH7jyA5WiegznZjqG3F8KjH+14FGPU+H0hivEzGetmDnyiVA
BxsnwpQ8vcZXwv2Mi+05vZ3bzLkkBy5VPXOY5R2jSJSCLXtdaJR9A4643uSHZHzfnzKUWDiWLL5L
oTW/ZDtwHqF5CZEvTNYTsMwD2ts+KtNN+fMto8xiXD/qe1ASOtsh5+zyM7ClYy2q60LIXSbjbwSx
WvY/Vre9VsMRIf2jBykwf3j5tyiiBFgb3JJYwQBBTjcJYbgJyQtop6x64kuRBoFr/L776pqTO7nl
Vl9gkkyvrYxW+owScVhc84M7DAvP4ytWKjfNYTuW+Is6ObyZVnIVJeokPJA30akb4iqGSvv/x9N0
QWZhMmOWpJXHkbwoBwaBlx7PeZYIIKaZdW1R3zINQi08PIUiRh9MVEV37nU4mskS+Bh83Qq0HgNW
Pxw/oqaCMWQz932yWKwkLTfjcZpRF8bzx75/t18di/QPmfqFhXx0N6r31HQWnfwscBfsbIowSPP5
K2KgzcXPWtPt3tDVEaMC3woMUZqBi4Lo/m3xUEphlRU05nGW2POh77X0dZ/8Tx7/xgWm4+v5Osx9
bsdQdidmilMAzq/eY9TUjG3vMfw4eqRgylQ/aAaNYjBaW0XMlWMTCOVtEp6K631he27e3f3jHeg2
VuLjQaimts5VLPl9U9BOnpI86SMSxHS7L+34/raSOizzwOpKnzfk37FyuGXTS/L1cB0bHtq+34Xk
yrjq5p8xkY85+fHrNJ3jjoX4+PDjPazBnVESNTEMbrcpvfzPTIqhpb4FssDEKiX8vm7hyZjfdUPN
5wQicX0aBSCIDGR1VyqU9qjzCYv/uyKettBZ0RHMs5p/BONfdiXEDYMHvvN8pqcbdBs8Fykq0Mvn
coY8bFsROaj21njHmWltYvQvhj67zJHrCKN9b7PIZ/ndg8AyiBM7XW0XgkK01dl+F3a9WMn+9qyI
sCUGczG2duhzirQKZFYG/ho0p2p0kUhUaBGJM32r2e5qlEQUalE0w9jqu0CVfrMPo7/b0DE5BkrM
8KeGv2uk7XPCIeAj9hF/cmZyTsbc+IYieHNQ5wK9ZqueZ5G7pOjU4Bvd74QEvcbFaabNb/d40lvf
pGfTUgFS/Y57aZ23/KodIUdcp51SdtxA0ZWEXg4E72KZFZEiI7SqkoUWWT1upsBKcyjRS2p3eH8e
UEjG6mjwx/PzBTuTW60OLv8/pit+dSF/Pq5cNtAvVFAUkXPFEOQTSbFpylaMxu/CTIvp0O4c4F7X
MAHPz5WoHXVA9W7QCcRKS9tLnkGGvuGyRUuijP9fv7JzD9tCOv3DzXgEosgoKpfxHoCOv3wyrj5y
Lh4mnz22Q/WP0Ubswcz7wA4rWewA3Ukv65Uheel8OPKjJoQBApUr12DPfuaBxT82pnjpli5L66/H
c72bqguKlHiZrmnwymeGpPcweCvng5qAPPSIniEhCkYznBiCjjSmTXU/nJZBfhYHQDDKlnHzTZuc
GnNCRtmFxNdQgMySA3BPeNYS4OADCcn7+HOjjWhT0vD5VUUvk/y/jBZExIXDZIFISfuyT3c2E5jG
3Lg/2Y4FG5jn04vxFYp7GwUitwbej9D9c/az8Ov/vjmV5kT+XVFVi+yVpBOvpUJUazQfzBK5LB78
lS6KbxvW3wt1l4ZF8Zf5tO0oyX3dY3LBaGsCwro+GIQ2oYmbJWuzUGr6stZjirs4XdmKusA9VwOf
sUpsLGdjCV/0IicqzrrPlLagdcrHSa46bzrNLxJT1mOOjfS81cfzmOVctk1wNw2aEu8NnVL7Te03
1I3y3erPvaO6sJEkkJGUgFJu0U2dqaZppr15D/UIN72NovjLmAbIiilBoXamaZ1IqlatqRElZkif
CXorNd7A4EQq38UjVZFnaztfhsbHHvGQeWYoGS5+xXZvo0o8zukIrEpIPkH/X3bU9jL5AEqTaE+G
oy4XcAUALmPaLAABbRlvu3AFhrqNfbs2EIy8zaMiqXFhcjRJ4XlZJB0hTgU1/goghLPsf/3+sDXA
O11qJFrmp9HPVGTC9AY9taj4/AkGGm//wiK8oM+OefQGLdT97qbaJRK9Gkco5mtH5JjbrV4gk75Z
44Ln2sj1W397LyFfjpyaV9/VSGdSa+TejDoxSsLdipw4eFNXXupa6/rFkDPe7uBF7fXgirw2x67p
JRvztUkhXlanfs5+t1Q0LqTrNcWPdgTwsCkcoSWfjqHmNdap6AnJ0hkBRMDfXxVgbQrlyEjrrGms
9TQflBMgm5tGXjBuFenJedz8yUj4JAboAkLwHIO8khMrFsO8+hUUd/fhKzK4EUdCiQB0iS+zub/C
q5aXoFbxkyCI/1QeCWm9oSMueyj9TBN8gDxAwfkTgypsz3VfcCmvI2tgzdywRwxyzJyWGYp3zO1P
wDD5EFYyfvDwLEYLOfw3Pih5tuN0blhkEoQ0jLXwNg82+/2rolZqjYmdCyTb2Slm4HgXvdj+EDTm
GjA3dZ7suQET6OQuOzyfN3fVJl3YobKuj8MyvMfOUrUL79KOMHqtSkEp7uRULzpTGEF2ddZfjHvR
Krcp5/b2doMOhiCZQAIVbzuD4wF1ImEzyFeetkXHWH7ELrF06kGDFpHleUtkWFqBBGvIyt2mh8O2
iI1j1xN1xgSSMBCoDZq6KtmwFj0RL/HwimZB3s8yKVwIjKH19U2/YsHSWaCkPDe2JNBXE/iyusmb
lpBjuVeIl7ppNv14j3E4bZi5jhrqmOa6jOGkoQH0aoSrP4/E56dHHE8RAVMXpPwdzvuA9Ub9tA/B
1hBoePBzd8G5oM+HCx9vJaXcKZRN7MVTYE5aPpdpNIVobafwWJnLbu2wZd+6xhrlDl3M37HJx/3I
VRz+aMU5BN54YZ9UU/Y1zqfQDOvFioIh0gyaA29cTnYcLkSDWBBTnhhshCoz1eqSjuaG9xe/c7Cr
Yy7MHTISnFjWqXOewMULgIzFCy64/eXV6mU6Ubct2yxs3WamIt5CAwol4miUhaYn4tpXsVgGvuOm
xYRPuUaq/XK86aDMdNIvjEnJ98+kJHBMc0slLYMkeZLCoHy+RK/D2XUOdQuUOGfaeuRtBFIPRDwo
PFRNStbpRFYjyHJcvyJNb6jGnxKMxqBBA5RFUA7SrqIC6JB4bgo1GnY+0SRhRZcdfLDKUylBcokb
3diEf0/2l11yGsI8nPWEcTKp5xsR0Pzq6BCaULTtdpbTJm6al92RQXDE9KLLZL5+tkGS90GK/WRi
lrwO3asF5km8rjFSDubxD0HNlBvCLBK0AZEvBa0v/ZnaT8eM13W0+mpE2FK1fFGhO44cU44wfQmR
oiHfljpqMovNgil4fiNxboP/bnK8//bLVTVkC0GIbfSNuAJDkHY9+yIEaRWEeruP12GC6y1NqjLS
2V/GdEcdkQSRbtLwLmQM4GWHhsB69NYoaQRg5zz8XyUTucICOX5R/tv2Fa5Ol2SwPY93aZi2otkz
YSdRGkZKM868DOziM6tp+4zdHI0jllsgdBuMh/GDAJcW3ZTNn9lH9Wk1pCNwSly2dUYJCp/VEudQ
eAbNiL+jNgX+FlAYaWf15KKqKlRrU9vgHlqBTla6LlTFmhjxLwH3zTd5TUNzY5aYLEytji13acsi
BO+dnAM6AK/YkXnJW4Or9+gGptrjDSIPGx7J66W2eo/pnE5ZnPFvmRlsqlxk9Da/qH6sUwptumvk
WVJ4Ojh+1S7VOqUlb1gAPjobI8wYI83lNpK6mvTJHjXEvYOpexDemqwNPcUoM27oL6PlvhE5O1jo
ROxBMPERQOy2F1zf0jwdVGf1ar0+h2d5llQsOjuDnMxUiX1xIPHGzwTKBvoIlUU7ulN/SLKX0oY6
cRsDwQwRaejGMAdLqE+wzXmsYbLhKbdy16LNCcA298rF6TTmajoxnVIrPJO0aeAdmwYcjMxGB5+y
FQYOtNOOPHkiG9cWLy9Z1uKlmjRWs9Hj+pcAY0eZXfRah3ou5QSAhD+MZzzMzXdAM6Jkxch7M0er
t/moDgU64hltkLn+m8kzcdEZJIHfqzTcwMIw2TDsY3ZFm41GEpzU1qfbkZvHYawk3OZV8bh0YCUG
y46y06n67xhharqOV5G5ahpRX1ArOKd+UV8DkaZO1eildMpEaBxcvFo6eku3ZmCxYU/mcnXzod/J
Gyo5MBRHHukjbM6ChIgMHu3ClWnWqwp+auTnG6a/jMk11A0/NmdwHXfMGdRrwTrX6Y8KU+U4hDZR
1F4onnartSNORydywWy9+c2O7cGUlxIKxS6Ng3voESuYTFu8wuRhWdQDuehU4LIJCTTKdxs72vTO
38W0RMMMabWddmKQCbJm2CAbByxkVe3NrM6DWvDCoDMYTvx1IX2s9Nmsx4I2obYTf6Bx3p4hwMhQ
9FmVcuS1zTgqCu4hJDM1Ar37RHjp0y27ZMKqpV5RmMMYuZPoOkqoKRHghSVb5YkfxV16itagRif2
pq3UgSH53mg4I+WaSlhSDXmZF+Ja0/ufuU41nihuUzr2jD582oFUd6c1a8X0r25SwN+EGR2MdUMH
rZU5nbyMSX1mgm9zP6uajNhpSa4lMO5kjDrOz60V4IqsR8uDqZuWMrnpvtyliF9itxNFb4L2sdvf
LkcYaIHZ0qBV7k8OMIxmC4owrbq6X99fqItlYkhZXomQeVDXguqTK7djdYS/A90fTVt0w3c7FCWS
FfxzAIa+oS6zm5CMedKT+FtfV5SSIez/b8kBN9smGSy+mdrN42nO4m28n0tOVTDc3+CCxTRY8XN9
32w1zKowibhTIooiyYkjH6ZRxsG8WkTFksAnV6u2Q6yHs5EvNqYrimEnH7WBD9cMppTtTIwIGPM+
VsiKMa+MwBKgOkWtWTXTak0rXRy/AN+4RRJskyRzY/aa7rc1SeQZRZ0t0mgPJM46YZFn9Bl5+xAZ
ND9o4iAMD1Ur1MKyX1+rrPxurVvUx6synV/bjcqpqVKAQZJnlGXmcKpwrFHlcY5f4ff/Qc9Bnsp5
VSC+HvpcKU4BHesEf1dg5MT5F+zxX8LSwBPdky5ugGX0z7PR+1QSrJSYCdjVP28B0YsBxyuTS8VF
C55ZRpRwFvdpPFW7Q2El8OTV802yAZ23hbps973stvLJ3CT9RWY1yEo5uB0zOd+XzD4d9pGM7/Hy
07kXpsD060Sgci+ZfK6iGPaByLXIywFlNaJsE/8DyEzyi0tiXgS/R9DZHXUssDNP4t10d+oa3hGE
zbJjIMMX4H1fkdDzBrr8oN13R0HHH7hEXYK9omQqNCFfhoYrS1gpZQ2GXZhXzdJF7RxF0bapkf1y
FeabcrABcToZ3RVKa9Sc7i6+UbGFv9J2VxtoEixNSgOpMnSxvQNfKbCvwr0MmbZmVNsLrUjAcxZX
HgDGqBLvXrVvyMdnoFXvrClqrmbOm92xaEK43E2d+RMxGTwWvd9MDvgzhC0OU4OEgsuwrW70FqZE
gG81ebxtw3RxXpyfPq2jX051mI2Pql02DvrHl3wgUgZDGyVCiC9eYNPsJR+WE5U+ifMnQroTwSkj
ggtH4im5oFsPLKA99vahuZW2qWE1GArvZpv40s4ui99keaaA/FMechz0sdi4cIG5D3mQNgm6xgrH
b5JNpbKD1dJSLtxcsF9OcZet/O1OJta9Jo7D0sy001qu69hYy0GTo79BCmFd6d+aFLfR9riJKtKg
zaDTzMU6V7NP9dh15AzaNi5sHmHRkDqgJ2Ru0VIC0mBIgTOHEyIXPqw64c6EhiSnmFCXNrMq0aT+
4nv/3kK+kXS0M+haxNuQxPPi2JSQk4QHbMgt4V0ZAGK9duCHP9/ONIUPhG3yQ2ZdGwoJoSGEs3qk
xSrtDzgZ6AoccI/2d2Ui/XpyjbJYNINWgfiI8lnoYBowKW3I89rMcr0GTo/02jXQDktAd22Jhqt8
PqpBkBm82TQ/LLD+DTpb0wk1ndQ1XzU4KP4CgQhUtiPeT6Ubx9fcVjDosnWnoJKbD09UkmyL7SUt
yOECw3DzLGx6sKXfS65SugKQF9PD4cgXPtvgfN6tU3UsV4TzbVEG31JI6sXW7tPY4xQB0j7toFT7
d+qp/fydl+hF22ynvVX1Knkk/FnfJI/V4GHZQkP6ZEq0n4jLZrb8QI6rmSkpzulxSlaNT4uenu/n
Pi3d7XN6gLEenPqkw8Z+5JAyZzCriIrjunf9NHXZVcPkJCvPPhxV+vPk40VA6s1xAeLhQhv2SM+w
vfjZiIhbPNoVkN+R9EYKoQCT5ztVLS5PWqqIc/RsrqNrDVoUsqECxEOP5JkEY8koTzABHd6FYO0d
ZtJNeHYT+BE9I1ttWO44KmEvFDZFszbuP1A6eaWXg6TRNjNykLYvJ94s2ZlSf/e/AJ48mDJXJdDe
3PD3yJD/UcGMa8se3LSszHIC1OfAFNT8hFrj06jl2WEh4zQDwqdwjNbMcwPduXjuYHsjQszqqg/s
G1BrNIy8PKJK8Ae+6AmO2sHmPndvn6ntAuUO8X8RkrGYgatzQDyccBq1xzsbCZ8iVjdZME03jdqW
tf6A3MguZVjDRHyIqGf+vwqsYKJzrS1Ie3YDmYQpkBT2pEnJRcxsHd9lTRIxjFXpqVhTuAuWdTDy
xXqc9QdivJ5BbcsU3SapLzZaOqVM2fUTMbeRxlfmUkBjXqs3+LqWMxoQCTZEuO2Oe1AaLhSifTRj
Kpibbt3jV/N66YZRLd5lJdCrl1rpVDq6aVpbqR4h8PMElyEZPK9qkXw2+lwfsyiyztuyhfiW+HdO
992msZDghczjoWDwKJPsyRASxPlQSZLRhDogvN8WcWEnTdBA+c2LZzPg7dIEU421thIP+NM6XbBD
lEYoOiYGuPIi+16g9h1xr2MaFVFmm7WakhhLl94Wry0eedrxxoZaPLFG0Bo0ZmCj4Pc4ZjUznbgr
n9NNvcuZQe+pHP3qPYJC2Hf3RC/2itZOvhirNuN7CK5h7p1FpIl4gwwCTImNmO41jjpG9o1BezQr
BaDSA9Y/023shucfrvnc6kKr2XgyroahbIUjcOTFrLdWGpTjEUDOjpU3CKvidRnBmPcO9JclN8Ef
uQkAQZ6Zt2TRZwXAJaCk7HGoJXLQr52wveziEphU/EzwzM5f0qlIrU9wIjXBJqmcH2jjAtJQxx8L
tJlezrt7pIBIEOlEeX1zSRzx9dL8AYtxwOSaC0L42hAyYjdsB9/TSDVEmUdHIaB2QHlFSmozBXyG
/rvFPV1yts+oNr8VH/NNLhCzTiAm8ne5vMwY/JDUAWIfQumlnvfDwPqS5Jq52r3onvjpYbdnz/yO
WyxImV6fmQcTbBav7VAAj8rFzaoqHk7RzF1YshYWtezCdHmIuG907/w1Ptu7dvFieFHiEcsvkthR
pPhrXT6GmmUK974lo0vXckBqf4EdH1kQT1sxvzsN7rWij0DfY2y8SHSkdzCnIgh7PBZarcNywJWL
ELlKQy/KuFRMEfswkxWeC1vRR1njVagGNBr3y7qymXg+EUepIoKE9jah696cqx2i/AIMbZBpwPG4
UX/l+3/mVeY4tEPQ1DyvN6gUUnI897fTzuNWWdbKkbgbBv6VWBOU0P5A9UnZzCAYOyf/esJcwPQ8
076Lh7kzzMGaL35rPjzeaYvNoL0SOe6Mh9AHXx5lP++RuQj7GBGN2xpG69PDoBhp8MhhuVkHv3vH
z0EUfQ88gqXsJ+qQMjnr9hD/Cm2pAB/TpVIJdPTlRuRbw3b13I0Mwi3xXFMqeTnXWIPUbM1HkXuB
hcmdxGUoCQUvMCPho6XoQ72LmqNOF7ZbCbyvtNtvSHj4ag+d1dthWz/pHAzldH5qKnu9cO0Zhb5Y
lb0JD6pa/CFea2K/j1u4T5SVUt/Q7OS3+DZCE/cbqLIhq8eX7pb3LEiIVUDMTlKdKlzhj+cSM3QM
YEGyGy/ldZP5FnYouzPQ9ohlBRL2knBoPGvxAtMVF795B82RZOndRDCbiurDBkO3o0JXKSNG10JC
vQQlR3Rovecsvq11CQ33ckbuTHBr7zPg1hplmuO2zvg+zBPG455UNvGW+QC39X9pbCxTWFU8Smuz
xRg35flaEZXptX6A22DgZ4EqQUvDbMLSidprWCf8B81QbdQzjseOIX6cNmbgn5OT8P6uFAN9jU4r
RR456sMiogVAOOHXOXfVbFhQS5Mt/y51ax0k63vC6axoYAMUpR3XOsxbk/SM9H4drMGPbMJ1PU/o
lCAwuTshaaB18wYPTib48XNXRIv68eMElMb50bYWSK6Iy2jJPLUMinXMJ8ycS1SbY6ckMIgDw52A
mFMvHaxTjY8SPBHG9wun8nnpfzF1cZxzuet6/eTsBKtr7VFrhTsl/igU6lGTx3MnF6A58k8x1y+J
U0hLz0FDgaF5K15hQnyQzYEITYoWvqzw4vTxqNiupJtkhfktqtMA8fZ0fUYg5nqbxgkQiiOLJfsq
I70OBMvUDn9srLE7qGPfgcx8DqiLYol0ktH1Idit4HGA6tv2bOdjKm1Jz0OqkdzgAHMmBb0wwF+6
OVmjfji3qQPEvfgy8EDCl/lQt4UT1CCkXjVR9D+9QXbEFWe4cpypJUnNsQSU9444RIa7u5LARjpu
oC8xvdzAIIJ10kvZ0P3PCI2i6NACLL3u7LbZzpbCyqKHe+H68jLhTVx9PfOhtvV7NhnpHVeMg7n5
fgcDAxf4Ad5pboR0A2DxL361cAnFGB2uhF3+zpJ6309JgE3slkJOTrV4YoD0Dz7fPGbHFSI9YRxB
YcWQNkuhYNPXDtMTbocp/dc1kX2Q3WzmyR3Rt8S0GWga09cEE2AnTVFlkJ1aCa5zayUziIE3+u9E
ikPjL8hTCi7SSQNk4aCG4FyyxA1v139UU9I1vQucrAFvhHn7UYFjQs/xPf2BNAl5A6E5uVAMdqkE
o3p1GD5Br5QPB51zFSFAU4PWOFyssdv4GcrbS/S9xfv7HrXahqVCpCm6h2oN8QfGwKlri3cAxJ0k
M0Jvt3Mp9Arkr5ttkTeo/Trds5bqf494VBvgZy69cViv+gpowfCb1QGUuNqVyFDQGISmomDrSjqz
SsQtNh8hgRQ7vhyYPXn7q1rHEzZtN2xNAXUg7YOA1ef+DrM7hsLaQWp63qLxtmYjDfz6LcEGukw/
/c8bZfMYLHnHnOpu9s/zr7QLIVfrZfp6sK0tbWrh62LGIfut4p/rw8Na6Kn1jqcIxbbm2/93Ypg1
72olm15Xs8tapcFYE04uNEf/UXlpYwbMA06I2Vzlm8/C4NCTpTlgsNmVDUMmAh9bXEdE+XG0pQH0
ULsywOe+DY2BgGZDy3463HgfHbnMtXXcU1rta8GlK5eowEcsAp9IkCMWi179kERlk0wJ0A19Jv7A
2lEQ4qd9uUCEnusvOgcrNAYeH47r7iHHYpMA3OUt7Qc1MjX+fWO2o7prTa1fUHYwO9BTll8oxlsN
qy0Sm2Pg2UflCtyK/gWDVQ2AVtIkB8MEsxW3CEBmiRVWoeG+7kogB+dF+f5RkqBWloHMEQJm6mW0
cU2I2Hrlc7EqNyUk4tm5x2+nSbvZop1RSrBX5eNTBJWxaAHdbq9hHem5uBfXzSC/+yAdwVOfpxsB
+lSxE7NJiPsKp342h9m9X1QyxN8P4+HeZF3glvSexQZQBCf0+gSZqEHiTXyE17DRPbL+KYXcfPBv
SBV85j7+zrOeRleX1KOGUy02K2sCTvMOmVQH6w1LqPda5lQFVwt4vLW+Avd+MWi6dPEmMEGKV062
QV9J3MFil3dSxfFrAu4AiClC/5z37nobmUm8d4Px2ac+UDKct3kWUYRybeQHDNoeP+iTtPdGJ396
f5hmCq929rQdf3B7pXTIPT9rZzTX2EDK75QWSKO9j9g9CZXs6F+NYnS8hjlULZFQZmVd4kLfa2Rf
VF+i7WClOPpkXNiQOWtlPYPdKrAqmJLQOxsRKUanuLC/+iRPvUC+nDj6XYb3q6MwWMXqgk9jXoU/
SWSHgs4nR2vUJk7n38+F7JCLj0itbCu2F23BCVJ/+6hCpvP+oRsAe6dmPwlPSkCrEr3QjqH2s328
/1/QXp785WbYSPVu5YRj2dTtAlehSXVGAeuSGsPNNzZaJvNOTXMHhSGfHrJy/jS1pC0ZvPT6W842
UnFZKiD9W72Xe6ziH1aQPwZQBiptrpmo4axpOSYA8NM9tIKgp7HZbYKBJZ1zXK+MwHa0gei07ZzP
l+Zc1hTKQNZAHDDvmDtfbQWbqgMUwFLR63p623nbPpL7X/dgR9FA6uQ83jxZvcM+qD1DSCzFVL2H
8fqwnCKtZ6mGyPJvGk01p957RCZtFsxu1dM4dDuOmRJUxKGDgmVGj+Wrze+n7vOsAqdL4ArTTuAs
1R+IIiZldY3jO6Aizw5QTKJwlWqbYY2PIZJQh0v7/SFMasg/3D22hiX0or81AOCmFnGigeOAvwjt
P0BZYqFy4bF8WEeplVuBkG7pDhnnHRHu/HpXFaEteJsBz5kD13PyGtGs1TpZE4DYiMr+LmEnAddn
doBHfeP1qqKrCE3N8iOpvA2cioRAgShvDLvH38sQHr/CLXOtqfoO9vfl186h5AIRaSvgGn5+cw8B
CJCRJkVlvGm+YdbKzDvZkR/u44OYxZxbQmJrESysCk9G33uHmL5ZoZnMcfvcr7X/o1CZ6lGbGiuo
Q1cBfMwYMuobFU+cR3mEXiEtsAVYLqfrq2/a4BgKNboD1ZJ6sxcE63cL6uuxLhXuxTEKEdX/4mZR
tsmNx3G+ja+BsGDmAJ6Dc2DTed8Cx4p1k3j5JJZoL7dX9zdGMjU7dHt8g5BZWjOjJCATSyyh+X+5
bOtML2Mejxb65Won2TLJzbMlXjdFVOVe3VRF4EU0tS9X7JPyI9fvdXFoe/Q3nxYo7WgCPn7V5c1L
k2FDGjierJoTNeG386WNUwPCBVLEL3DEW3yx597J0IAYoEHsSKj2bJXbuJrCyu4//jJz2gDtI1T2
Wafqhw1/WSj6zp2x1+BxAKpuYYLjrFWZO2Ht3x327cYOulMVXkYy/pF4RNfYQoVt3Z92IieBXZGF
NyKjUGZx3BQCl8u0PBLTpndioMAVfaELku5Gh5u0ENOvSSN4TzUh4/Yz/IysS6ATqg2l8UP4cXfr
+cJA0/zQcbeir1uXJ8fM9oSv79baXVU24AH/Yfn2vmhPmZyO6lWXpQS5p3x4luyvV711WaLplh8O
3emt2kIUeoe0XzuPwkQIpR3zm1uJgAMB7OGkyhe2uLvAIBYBNI0Xck2LzRSYHTffa7GdRfKAFUpD
gUBlF7QpVky/E4EoQuEQUl7gXeztf3WFHLQM8X4JdMmosuSYn0Byd2ZzqELN1TPi35IdfQmlolPs
wWvQjVT7B4M6LWX55BzUGkR/By9J29FwuCHIJwQv8e7oSn25CeJNrCbKrJWsMTy+KNqhL2Ofdq0I
W0F48DG01NpJny72c0dItTcqKvttyoVi9dZaY9I6ensbvyWj8pf3LmuzNtz7ITbYVGCrNtMYLIqw
x1TlVPWYTotsFYIfosK23bjlOWyEGWYZiVfKMu90e2uxGb1FWBXBo4BK6oollebNXPupTQpGpL52
qx0XNxvKtBkkBmw7FIOQ2jfqIB61gBRB36oRJ5L+WNFGAnB9WYDXU+1bR5f71bLTVdivfqIaVmXB
zpaZ8ho8ZY3009ZlIzZCMKnUWkk8POJf4/D5+4xY7lHvPVooMV2qrODCKJ96b3n7PWzBFmc2NXcr
1vnR+xfOa9JT2dUQJAwo46/maU8M+Q2x4uf+yLJqZTlcbw6kg/9MILntK236BCzBYogvTCfTOkio
wYKd+ljor6IyvqsSG63FBRkTvQ+ZE5KK7Nf68oFSjVHWPDSBn+OtoGapUisNtSl5NW8GWFp71GLB
7qTC6dQjPvlS1nKzoxeVrZcV4MH2Mpo6ugc72ge3260Vhtt9MeRleAPb7emVxlbuzKRH6ZDMUuZy
jYhmf8P4RJrvoVJE663EuM+4MYuPZBxiv4trNeUAElfvqso5SZQ3I7Ml0WzfwrWCXVtfugPAm1Ok
Lg66ULoRBHBJIPs/ylIRk+lYhNRHTrR4XHyNSwZ5BMkhM8G067VbIHb0cNMEEUlsH4LY/ssrREx8
p/Yb3Irw5RWYQh13yUwyRXKfnnyQfGTAahHuZCx0Q8jFyfnio95146umW5GOYy6Ri/dW3tbOq1Gz
U3MFyfXRi60cv7Y+H+1ecBkjO0/+jjB8WJ/jW2wwWySO9RVEUyXA0P0RsySb9Bt5EL97tgHtNEnz
r7ZTGpZQEmt9i59Y9+jEfoszxaPhIRuSasgGB9EY6yVSTysqZPah2Eonnr+YpSerlKghdjcZRJgT
sE9H3RLxNazn9kHZlYIuN3phl1+YoyOYxX1dgg7jcehBzwJ0SERgsqh0Fdqo86z2kjqH+3DI/NxH
iiItdJdimGIC+SXLKmlWK7GDSMJIkG+RIEEFMPaKlogScfjCbHJsPLn0JL+XoBV2z9WQlQGTvnf4
dodZvXkt4CBv46h29FScYY0uzvKR/1Q0C286N3+2nXACX4sZVrKmdFbPwLZWi0aBTfEV6WrDbGGO
ciLEjJW3Xj7srIEVaSmgjXW5B1JidjOqlJQ0HszKObEnMPmcZnM+3GQa9az/Rxe1lwXE4JmuANRd
lLs9EIxeKIglKBLDLINJ3xwpptkCd4EIPJMcwgiXxgY1dT9S5ojc9H2bcfzWmsPTMILvCHrqnaco
rfaR57+2dk2RkI3Zf0EX7cz7v2kBXAwFLcJmoubRSsD289SOaCATENG0EdeLk4DbN5j9sPb3v9Z1
EIOm5MyPwQHb6c9VnYx2LJskT3K45bP/3NJNifmzEKHC1AtWY6AL8H1MW2/ZbVvtWfSZqOl5WQ2i
wPORzvA1DIoOOyIZ0ATdLDKAHWpzpkAYwca6dUOxI54bFOoTcE4bpi1V1G/zewuw98COnQex1QnW
m/mhU99aK50/1BhB2i+qeYofzlFIyGT3s6q9qmmued/7IbqEvZCf0nCfnGVdulHYS6MQUoyLD1Qs
FhQy0sCAHVrAwF1qppUMP5UADKRRfkecLaNhvWbrrzJPCaYZw98DVOyqBmK4qkgDwkmVB5KzwrgL
GE+WpYUA7YaVIEqijftVAIJEYD4IgGDUSZ7fG9F5BW49Fbcd0VeCNIBAXI1fBmSrvFwoe5Hi7EGB
7R7XC+GlB2Mtg7pNGCJFFM0S2N6+FiT5Ynoe7HuAtQsYrClyGJ/b+LmWdFA3YN5s+0vx7LaYpq1Y
aM24YKzvKwZyC16VSrVgQ+Z8aGKFNeed8nFz9CRXk0hQr+vKxe98XayA7uyEaKHTJbRJbJ6LyEHL
0xCnvQSIi7BHHe63sKe1o6XCr52/toDqA2GqO7lDIC9UE6WiepG52zrzHbEL7N800QzsWVdm+9QN
LIRzKo8f3QUwX3xiJg+MzBLEp/xx+L+1VZCwbKDIf8yF8u22yzOBwwHU1SjvYeoBLaw4RHt8wfSc
648aZ+k6a582R6z8Zdf55R0Gu/d0w22tzuX3Itvv7il1RndXAABEW6Ra97FMsznx2jUbbAm7v3H2
woIs5glUmur6aCF66HrYUfGF83FBRdxR/pOApkCljnjXsztP04SxFsP7IvtZb17JyFLECUYYzoCw
Ixsg3v9LvdpKzvKUQsuxihY5jzlAxd3qz2ky11g/xW8tT5epR0uDMBaRO0Sy6ykF85zlCZgOXs+g
Bf6ri6S7VZ4rZxKJpnNnDDuH1NzXwoEOcTLoFEaW6C241UiK7o7z3w//DOVj/Eyh3Hrq7zKxxRzI
W64/8SUTvWAoq/UWJL0oAGJW28+cugkbqv9eZ4CQ0f7qbMd5Bg83KMgBoB0KxxKytL6Q6mPpFKRq
hcD2Xgkb+cFrqUNcm4gUpXQKUts/0CySdWgrfkOzB3nwn8Z2bKenjOszyx0lyOPVlbnjIuYWgndq
MLKt/XoNlj7xzTRwWMuf/N20VTUXs+bB54OeHIwswdmsCoUjSSAXzRe6MYckJpdyIrh9pmeyjpmQ
ERiCZ+8Gp9Nv9329VfrSleIyeQYJEdC7uxdsKn+3llmqbU5FruXa3MEDGVqv+YCUEU+f/4HmCAbn
pEjrWpvcLKXaILwOfLQ8wBJdOn8V8PuLjKOwn9RwPNff5yI+redylxyBCQfFtWs0R9qgRvhfjomL
gcZ+kPDpVR6i9fTdaxEODlkKtqsQ90IzW+M52T/wGA2SNopLkeaZ1a9laCxB4FzYrQdRd447ZDn5
+ckCVvlsieXKthnqFlhvGbJ8PM9q5TiK1LvgqDwYZRC32HnRCDTSodNQUpXImXbUSgQju7kanyS4
xmm22SwmVwuJV0VcSOCYSbOmMrtmjXgairbclQiPezKVBRsVhL6b1PVwMSWXsh+ZrXDq6gX8Fqq2
MzMAWbdGxO4eSxmRiPSuOE5N+a0JSKyGthjFKIASxo//VRwV7fktsI/Sw501q8hnJ7ih5xAJ9N/x
la5kWk/HdIPCRiazmQXEy9X7GqQ6kS8Dc+IZ9IjK9U30/Az/MGbCsvomButKEHb4c0/LdHvxiLfG
fVT+jcQzzzy8C1d86Znu33Tlh1P4v86xFgsWOOOxRrACFGjQUE0SfN2eFRISjn5uggeB8tHO0Tzg
rPxs0t6iHnYTYydt6reTbNgrefk9XDlsSACVM1oC70qc1LswlktVA4f8n493/mn+Zu0vn8wuSEkm
WMdUWQMjp/w0tRhLBkI7Nwxt8f6J0xJbQMudlxaRC8uXpufoNZuEg26daw8BCzROSp8uAjBQb8/e
LO1nIBA1tOk0AXheCWWjJ43O0j6FUtuhBC11lSvK46hJsybwcM71zTZU2EIxOhG7O5AJDM72GPeg
ZROd+0NFFuVO1+PbvKWg6+i5ez2wi8cEN4oIo+o2pXV+eEy5WqMiEgGIAH881oVmo/UDruB6EMll
SFcp3ao/7o89HbZ2vASVa3RFKG3YLmz/CreSd91RJQRrQZ0FMqRf11utCVUwz65zweAzjYQCg47+
vxxb8MkmTghoFqfLbDXdWv6ursSAr8eIGmCFT0YoGd6agg8xFPFU4w2X6RsS1oWjGBbayvz12DMV
ajbHsxlN4MqQ4Ma4m6xjTMJMWb1Da25MlBH85f5jeQ2P6zxdoa/bWdOxFl8ozXVivTDWrdxjNUTJ
qek9KYTkY0mYnTzTqt60PYdbwOKZIHbBfmHds6Nh/7lM4knIYkn2Y90cpXap7qXJ9CUPbRf5L2FG
KJG8QefsPLigpYpZ6VVOGT/LLkEJcz/llKQ3pKvH/i5QuL3n6SeKPzgFUn/G3g+xmzlr5HeX+tym
u7o0XQvHI/+HqYrT+SDVvZ9w56tkkII1yiGJpGdt8yanb05UrFeJ9OCE2Ad7VvMzhsHwLDFN6bKB
pWu6TdR3T3+8XZXwQqtLhTWTlcYf2lxU154a3UIQtyRmpCQhzTk16aiNpt3M4TDWeKWsJ6cR1Z8U
dTKPz7BaTpITMeSd/Q/3P84HTEHWxqEh7PY5+NaU6oeen93jvWEOXTCjM7CSMJ1N73vqrLZtQOVb
64KNK3WrAqk1C9b/9p1J/tYQYkOGW0658kBxrbiEWKgL+Ez8pq4Qv70C7E4ugOcY5ywDQLZoB/xo
wZ+R6Z7HF/pV/C1jNwUysX5Nq012eCiSnB5rAooWmk96H5qt895iUV7zIljScxkYFxZTRv5wp9o9
2ZTP8pxAaZ5yj75Lp68IFOW+FUBsiAMO3tl8M3rYMY6hklze4cPZNZsYc9ZGIxxVQ7hQRt/qoFfJ
T0g5RIjQ9NUDtLgnl3JukIwqVdA552rQzoRDCQ9YUOMg9SwEHEzkyjH1Gsg6KannCOeNS38jLnKB
/KuWS5fxukdS1a1vUY3791AIk0mGbkowcg2NvnY7PPPmRA/kmXOrllM7pf8H3+Ux+1My1hUCJIUT
L5u6aq7ejNHU30aMrsSnnFFIuUBeWZlvVcv8fSNFkS2LBStpqLI+AkshGjqor4vwhq2LAyIVo98n
iVCOrWPhHXag+Lg6hlMzA9hDy1kXbhqakoyyVNvq/NGQyEuGzzLFwnNiOlQRa6Ak4mnj05rpHoPl
nY0UAHOOWpFuA6v6Qs53LSWoizdwQH+BXWUfskQtPlBDJp+VTbsY7I1bgL84TRXYfbcTxZddQ0YV
d3pkE4cj/LQUNKtZ2sV3mQzAC61bs0ZI+KtpD9UOz/xBBLqGXaHlv1gRDnczD914e0VV+3FQS8wD
vVMh/R8SRSPkHaB0RhVDALrMCNficfBlBd4ALqxXLDZc6YwJJ8LbQ5xE0OncAQn7cHEA7rS02/l7
trx/ElJGqLeLGotzsiZLsv+rYAe2QT/HDRdydVByfCozyHygkouXjSChDpKdLsw4+F2B6cM0Fi+P
ItMW7HaQDaWfEFcZrry+ItAb1QPsNmJmAWOBHOs30YBAvKe6nzRS7Tw9L7u3xAqYYylx7mjnMLaM
ir1MYzi3FpyWQXeE6UR2XjDUwUKzeK0Xp+E53Lnp0n1TodLPzhcj5zVZ8wgVqzRrPiNieEfptC+X
OuGuicpTEPq9zG3z4+uHNHDgEm1C+NIJIgxk0aFU/fueFnG4N9P0G8djaWVDUevu0KowQiyx3cnr
DD2FxKlgFiqpnyY98oy5fyT9UnuAPf5J556eFf+C4CF76bxl0z4Us4UM2mTZI43lkz6FFg+ZOBp/
WFHtyvJDeAwV2hXUXB5m+YaV1N3TRzQ39fWP9b84Rjz7m4HTTo6etW4B4OnzVsDo39VLNysIOqhS
+XS6bkJxVt85VRRirX6hV7XqdO2U9E21G49nZ7o7vUAI1qAFKurUi5sTB+vQUjfL0fNYorvk9MaI
oLh7C3Y7HuFO6z+fGjxvAbZ4QqlQbaiF2Fv1mzXnISyAIt8Bv9Tw82AnyNCiHihTyumgT/++I4nq
IWujHtJ71nRWh0ycFcrSpcjEOZuibw+vzLTGT1sP7wFi2PTNd/nRgimOsotb5F+Zbv9qRvb4/GG2
g6wnEJy4G7te/XGzvitKUSOPe4e1/zE4LJOCmjIVYEYIyNCapmcaqMzb4z4utnKtVdGZYDKaKE9R
isw0gH3VTlz/EpKwf59I7nASII7fskf0/0vXd2wZw2VMm8rHwxLCb+owlKAx4KtHrn8i+JQqlYLW
jlTbUdSjEiA6NnAE8F6Y1ImP0iQvZ1Bj5d58lyKV1lphuJZwV5I3ORNkAWMW9YJA2YPCIFdOEFF3
hzh5gk+POfGUVQiS0Tv0wPnAAzF5/Fl+6oeIti/dwmyjecE8MpA4VsrJ1sMVC0SPlpp407eHr9he
ZwPnfzn7UsTD95TfR96pcgybmaqxa1OMmfLx2Hnze7zjj2SGFuGhdHr6zy9VrJrDGCrNrj2klGDn
I96q+y5QorKDPPFicus7K1SvmGAp/Z7rY5hBKNGQeTNmSYDHmR8Rr+mlUV4GQhqR0StdOA4VTRnH
9SwaBVzocLpWs4kR2IqWAzCLJuktM3cQfrrjXrBQH5FUqXBstXr2vKUeZprMjYFVNNkg0PaM/T0A
NQcnm1KCtxWiZGm2s80p6k4hX1GGNHLpeTVlvaK3y1BdZzhncHm59ZCaIcXVBqF00SWkRPI2oG8f
wnusg7//v89sj5vAk4IMT2kDqJ8l4lVMh6quTl4nhny9t/7oK6lcbmct318ao4KH4svV+RmVoytc
YBEkfQJ7dHU1Foqavvmj8DZfziGH7oEDO+ubW9sziuAflOZ9XtkrEUHq3ZVsituKHfIfIgqOtlmG
ew8pq4Re+LG/Fas94uKEqtHhgPKJgVUsG7eA6xiB9qKuNVp/w+guy/43NyKQGqVxcjzfymCaxo9y
qjw6ll7P7tVOVvpxU7P3Nc5/HghCvghu5M8sLWaJfrwRoLsC3v9qqRo078RMqWcrLDRCG+IM69f3
PEyHhTM/5KyYGqr2Lw1A3CQgJDVKZe8vMvEa8Fs+5d0bxMTxHPOcwO//2E/n7nBDyloCYDG2VC+t
zlOu3wvLPjx8E82DO/WTUMooT5xTSj8p36DGgPbRlbRaMbRLMI1xrvuOTUREDaZFEZepLlZDrF7C
hKouusDbN2o9VpukJRpJSC4Lf0nwHQAF/Dkn14a8osSgcnN40g52dVLp+S2LWsqpqvXJq3+Pbpwp
pIp2y+1WT4GWGOreOit6aK5mHsQ/3RMhgEQi53bJ7oaJNfyajfJsj28OMp0tN6P4yQuOm4GlvQx6
MpKefWMWeGhirVI41BSeVLd6hjWZEUPoDuH7i0RJN+YRLDRZtWs5Rl1lGWTUl4aUIdUfRAZKFLXe
DYPhgceyFEzUMeMqMeO0PIgX0AHqre4y5+DzKls751YQFT4pEdmJeLFgjKTIMuU0wYR5FRS9I0cE
mMzcs5E1mr5rWtaXNoQLyEezbdrGZemZJ5XR3tFpqIfqB3MxJrhGPrP1JWBSQmGO+VEpZvsLqfRs
3lXEfDnWhSOQP2EC3INqzE/QImbDRuw3DSnScjevz13847UvVygN9SdAdDyl6ua84KB0GFfiFvvS
PqipbnEXW6AZQCD8zf8qI56ePPOsls3rUnhpGD6iPLFDsZX0ULMD0uRewed0p2b1KmKHPZx57He7
b5cgWo9wkGQ5kO8//70eUhq5xvLp/lVJh0m2fA4ZQYoUTsJiO0KMHdxzrUlbT3kL15HybgyA01PA
Qsk/uPXDjIthWc2INOyaOrU5dq8jwz6aDGLgxyN0PH0XwiudfZYv2NvVW1qTgsum6o4wKLt+n/IK
thdCFaAMJsULhNoSIPjdJKC1qwwBk+Es0a2Eatcp2u7fxc0YUaO2cbQbVLMFgtStI6KcXHNd/Xnu
zvhv8bZhsjntB5R1kgHI4Fx6unT8Jo9ZuDp7mhqp9/G14yvE5BxLvCEYqoVJVTnB4TSPRrYKzodo
MDjR129uhCCLmADF+01ba5SufPzrBc+hUqs5s+2HC0GOCLDh4UkIqYAWQvRwJe7SXQZym7BhEB8Z
Cc0NZS7n3O9I+tlM/a+SXY9wcZsaJDjk5OmJtun63XCVM8q4X8zlmjJxEt4bp57Y4UnsGUW6LHKE
7w0++tIDUQ5w8kz84Zq2+Pl/RD3Uprl5uZgv20q1Fv0zJtTHvMThVdAvmAS3TABrmhK5rkFNoEMB
sLbxBtBKURrviFmAjsVDzuhRmbtI1FzCKwJXeB6wPxNEXzv3JIliP1so89FvoCzdoMb4xO/ob5JQ
la5OFK9KG+NrDOXWAB9kdyQozZvL/cZv2UstpG1iUlMbTCTBzj6gaFqdds3qQBKzH1xEAbpShmfd
vj7NOzOn8KkYodGkaDxfayl/xliou754n2FYkz9TiS27sxafJZH15LqJOfJ4uagBtFE1rrXuqOoN
pfq2Wr75M2tT/cUC6D6KUojoiCkRuPsCJKBYzGxJszvAbAVCpRURhZlqDP4zJV9dwl6w7sdQlCib
NSTIXB9CulVCCDfabC6D2lrBwGhq8jkDZyCjrvCN9mmKnyr2VjZPyYmwXq9rl13CuJQ3buzb76Is
cBNz6lZMMDIhqK16FNY0PebHNEMmHvDwYV+hs7fcMmdDKHvvG6A+ryvgk+KOZMmWlHWZ42czKS2h
ubRqwS1/WDo9b3tO2HosAJrndA/a8ffgnSfC/TMcPXIITRx5NsG5vStQUFJDdsg61RLqOLAgs8sv
a7iobwZxOe5LKvLw33owOP2WaXBoNfyuyYhQXvK5+tK7rNoAIL69svdEnSL+OKyiQXVQV601TZSr
2XODC96q8/NwUusxoMlcTFNreLmakewv+s110+fCPpPPEWFixtjXfAJS/8mYjB0FsLWIsffRmwEW
WiqUdNxdv465EDDISnaWuGbKtFha4D4mFQY68K9TPntw2IJ8thyf1R3laZCG5Kz1AxXqoWb1lK04
mZMySOqNblGugEEUQylVrYxZg/9DGKkiGdCPabiU3VJCCapEq98UUTwdngyYvZxlX4lttfD5axa7
YstJTDX6cQF2wPF60SqI/CayOOmE3TU36YEuXjdck0W+3OF7+o1YmldhseAJ/31JBWp56Mx7lsBz
HxVMKHO4yWfZiYP1BwgUssWlSZqXBRZPHKTkl4RQ2SSXo5oDiFye9s/bPrHlc9zqUbA662Z+RMU/
ls0jyH6UrhJZw6pj5QMYnZKr8Z+e1nR+magbo7MTHqG3tu99yZK09VDGdzfLuh6BlL8kLyP4szEt
/0u7Rzb6O5OeumkrpBb5Y5Hyl9CgRKWKTMkECh1J4obFR407C+KDMknlX2uxgonuEU8/G+2hFET3
RweQ/nIOaub0hBTVuV211B8rR2na+lHRCPnPf5/E5aiscpp5KN/10sKTsmPbv/vv2lANTRvXdwTL
0GMpIgifDXOMq/j74B8Q5MRflawbR0aC4+G1VY+LV43C65th4KqIX7colnJzph2zI10IA0zj4O2D
JRnBbJfFLfaU4jtLsd4LwF1MWgoIySysu64vrGqezUVzgKE7q52xa9K7m2kBFFMeTqGpCNCs7MP/
A3mtdxuj33lZlYKoWaH5iv7LRAIS1C8mQLaWaM7cpISpVnzFP8UkEyIhw/Z2L7hM0H7M8JMfltEw
iGLzJTi9RRyCo38vzH1AGkUCGhHVEqt49D6Is8iFxKrBIMi/JBfyjTsAohgj+xdnhgTr4+3OGPLt
UK/sgjWkCjk7oDNvGcqWsokTvnAeNHUGz8jWxdw0LRbUNSUEwJC/EKmaPwgtwIer0QYxh6/gppzW
pAMuykoKHwDfQMbkp6vk+Zp6/mmULsRLfRceYwPMmgMvFG8uGNgdVGGWZIySsy7sjJez4S+jh7oo
NRRYRjTT7tji0K3cOZkN6Vb4afpS7PxBNi+wXT7rHRbuQYWgmRBk9bHUuqy8XYiBSL0tb1CFBIXH
PnyYgFc5xeZNyM31l/YIr1xWaipnA1OAeycAV2DEXjv6Z1CfnR7qAVnxE7fXk7QGqZFhTMjSH4o0
SPTgFg8QytaGV7gjxyg2jtHJueC6OffB5xUmnOUMXrF0EYfWH9U5IZdFT2g5wJHy+kHbQAFk70Xe
K7dduJukhWmYlfft+eTWeX26QbYtKfcC+GwKXnIlRBaX66mKwRAvte0QQFZCjO38ouKhHamZMncF
gD+dm9Kx5yVOZNQsIiivAl1or9RQfRWsfXfXXDFA4FgbmvU9vcZyjVzA6WFw1gFe8VLd1UIKxZlR
a1ZBkaCQCsmlQmSY2E4CONN0XaQ39cd6LodZ5uWkXz8D25mu1lAhoTEAa5t5hfgluoKRMbaP4PY+
F1jTaNDDvHy8VDLgBt2bA7UnnW8qcQriJjjug/d5KJq7uAXUmjHYHf0hp4Blxp0OI8RldHrzNcVh
mSJIML8rjiee7UHxVMh3mgJZwJum7ZYQskUOqJKt7Xt86f8T4VT39X0cOoe2Jr631+RfOLqeL9XB
aDpFtcEbR9Lox8EUWrINkz+IVtFE+RuZYHv5n5w5UJF8wD76FOit0EF5lftyLpRX/FuT8PLUbwAA
HcO+Uh8mj4ADtJC66LFNfhYfK9MSVpImQ2UM9vcFIQWMcQe69wB8MQqIFba5pzvzMzzQR6dCqq/l
ucJibkr/CWU2VlpPSgdJ1We4pNfmmrelTxSjNKwrgMyBEfhWM3gd6CaN0graAEvb2MWB1ZRMIfCp
xQCq/uEh9MfHHCB1BQZd6A1r/TbyU0NAoRm4l5gAnkhUC/SqACCCOj1wJoMKxm5++wFJgbLBiOsI
Gu1sj+LEUrt75hJ6sWYcuH8OI0OBjcMjeUtSHm0RFuji03HaK1WWqdeGqGa3hG+VPzf+Cta85REN
chW40FtRmYVbSF0W7Uu33DFRhkx7h5E7fqwlLoURjPzlQd2gp5RYaKlL6c3UbxF58TO0MyJ5C9IZ
bvJpv0KIOl1JPDB4BoPaeJpuNx8ktsL5ZMQLjbjg4F7x/NgjFSKFWMlcPfjG6Hoy2GkvKCy0qfud
M7wanW6PCBmXQU04B38o7UkuvrUBgYnRqFKy0UAZlj20aSAANKHc9NO7/mVsFZMSo/YQj7YiE6AN
PiGaA4jH2kh0/kHtJLlN8XrQJCQsv5QNX6HGgwO/zTi3X7FfbeN8B66UvFcgFXTTkHiUx8x5Jcbm
i9Re77btxlepT9vrhGmntWWRLTwkhsOl3Mc7DPfwA0PpTMFERmTKUxqQdLtUWDGTWSge48L5ZtMk
Ec3nCbO7quTH1dY68tMqsErEuBjzysIN7GktP63j8K4CTu6v9afq5sObPLbtH56JKcIXku9TBVvD
t+VdkM4nIew+6OiO1FouzaU5iN5jdDyUYJkDZpgQtIYBJJVv3bJSMI1NY8JCVNLIoIshD6oYICK1
oeOBNHruHI/FIy0FKEvf+lnN73RCG4vQ/Nd/7m/DqFf3sKplsOUGWDh3hNNOfDIQCc48zPg2PnQ9
rPfzs7Vuowv0iPZ0yG80bz9w8uz+ruw9Cq0GLAPdMnZ/LJvIhI8qsKFg24wezuF8iBvck/01iU3T
FWq54NjqwnoDj73S0DwpcI1Sepjf7WCtSu0CFc0GSDyuJfACjutfgkRRz0ZLgeIbY+kabYS65EL9
7RENPi24o2TDKCb2vhvFkGYAbGE4XzU9cFCuSv30gRf4GUOJ2othNNEA1fylC3YOBLfDFN3yVxtJ
7gTq85buwWSF1vt2JDRuF85qLGYxCPGdwLdsYItj9BQHe/5lWdg7r2uqUOaMc6A/XKsa1UHcXB2I
SRcbajmJE5KWmPCb9RLhyZXAivbnl8ByLgRd6pEF/LLThEgnsw3eIBAFSpfNFbtYk1oKLbgCzYAT
Y15Oti4riq9AielhP8gjlyx4aIw68Ny7iNAcOIhW9cBUh61EPpb7LmnIASspDtaMuRouxDaLc4wP
SIPvo/HeHVVGlccSdzL3MartQXwpbeFiTWg+ssXNgUSYwP93X4vR+ZlGscIWA41266W40TgMLECm
hJE/Ir96FznRWO+NG6ysWnRp5PX9zBwg+5bXZ04rSe2/H15xMvld5Q19Pf7zkrEiUi4n3hc2rlKC
QkKGHCQ+zvMcFW/q8NfTe4mUVGX4t7tGJQ1nCTi9pQfi5+Zz67oeWcaj3mF6uNhC8fVBCcSuYIh8
oyfedLBVd5+C0w3ULPDWzXAXfJKH/4aOgJrBRh/YA5E3Wn9NdM4+vOqZQjTYU1tnNGNQynU6e3mj
SW+Wvvzp9tiurkQwhv3ZPF9/yxb7u735n19EV76XWR2au3rkHI98AR1vStWB7U+iELmLK+VsPrbZ
4PMdXfKBzgCH0LEkfKgBuUQ1zFlAPq2nrrvrrKqmTdQtbZlz8JaFu4gXNnZndho+aOpIDFPicrwh
GZdWxd2FArmTGPQmWKhdSazuYaxJ0d2S5qQqniPnzBIdf2Ub+ZQEhzXxHE+zeOCxyAaNmZODX0Hk
2Pihdi4U+UAHfw/hRscuS5Cmono1UczDGGHGeZoCLzA0HkkNY27gidfmKFmmrhMJBv1Z790RHyf6
dqKEkK0kqvhqfXyPyDpo6XXZbaMM0DowjQHqx6kx3wMM6eg9b/G28wHNao0/lPUMAeMQxck2PzqW
B53PAgI1EpKx+chIKnk0ADx1ox6q5m2p84Lt88lDvVFyWMHX3ELiW1kKbW2zK3jB/JW/YVsywmdX
BQrhJ/ttlix1l5F6jespq8n/lFT4WUP7PkGDcZTAFO+BD4fDg+wQG6+mNTovjs3/GZfmijEZLQvj
y0hw+20mP2++wd28RWz3kbDEJUgtltv8qKUG40SFNdffj073mhCB7Sbpe5o0pjaey+Y7gx2WOV9V
V35izWvuLqV0V/PEBRSEjr21pSauxM7N45StjnTwf1asCXxSalweA7pTD1thjyCTP0xuwTnYSKVI
mmo4CqUgQs3SemG95wh225JdOCg2YB/9De8D2sW2pm7VxK6/Q8sw9V2HX3R4nIMlVnnJhIoQMKw6
pmdEN2o/rxLUTq2tbNatovnCErPFXU/qAYvcyDXpWwS5fZWxmOKVWeLypR5DaVJ41nnqBFWZeRS0
Uk1KFIRvQu360mQG/cZlPzmfhXoSFlnHMBw3xtI1kal8tCwrZhyvUOztdOaIZlfIoj5iakpennn3
kMx+ks+aW11eIhZ5/iPzOqcnnqYy/Q7OfZMDsthEKmoHFDjjNChY6mbSWLvOJZUcrrM5RdSm+Ysq
aRkRdm1jGTM65vA6f0Vjg8AlpOdo2xcudsFfHe4Pv5pxnVc7TcCEZ4mVqQBD5VObvXfY5+F5Fvwj
twWyuDhT9+cft/93FrmM7oHnhNfg9AZVE8+p5KbTbt4VYFkXQMY6BeHQaXu7G8Dbmhtxk5D/qxev
cXATREGEVRE+vJAtZsDFqgkV1OcOHlaiO6Hy9F4wxPTl3Wa6oxxW6YT0t2/jaDVCG31xCQWH04F2
cFTn3SUF5L2vM5JyUcXqsv7IrepBUfT2dN6SnXIH7ZG6i2mEHBBP2GENam5JNlZAykRrkmJ2qNnV
a+ZbQgJ3iSylK+iRTi/Vcw6WU8jqXt29UL71j1QzQoKKFxCb/OJ8NHzZZgbU+AVhCJK7KV6/OmY6
LeT8qSkHfoeRKYWUuAI8EMlruSsbgbd3EqGREk82D0W65mRqrzytu6jD81qPDytEUFPe9Di3CD3s
QDWjNKIc1jnyyiQ8cy9WAw0hwD6JFecIyqg1GP3iZN53u8PD+JQi9PUXG5HTM6BQ6266XuQoU7/e
YpFFazULNnQ/yQ9zvVBaT8LAOO/zQ3YERVoCyHZhT9JHlggKfdGzQRsJSvRjfduBVMjeexRH9yUk
aKhD1R5Kl35EMMGj63S6GqVBFk3CLx6DwYHt0WjMEdLQRWr8bz+IA75w7G6rcmijsDZhZegFwgsj
7Zh/1fQ35E6vwsl59wlw0OxdvqzoLHbV3UytVXyRKHgNCt5sXHhURvp9Du/tRstXiKt8mwT1CXrW
oYQQUqDSCIJ9na0G55SrzyiZS8PojP4Qug4iw85e1FgcvC6tW+GVV74j/lCa4wmb6kGwHgEEIgt+
yEN+BmX/Y1hEkOGA9ahnNaaetfipnnnkRPhFQtXdNzArJIzUTxOgIp03pKoDJdrPUYn+p6lIsQlu
0lzlU/TAPMIV6hatnfvbXI8hOTUTMfQ3i4f+y4ZFdo4OVxV+x6IdgT93pZSv1NXN3TxAUa4VM3Kc
vOekHq+wcClt/eyHt2fY2pRsnrXLyDKgOL/iYBNAxU0l72eW6zKPfl00InH9R8AVpDjsOmWvQN2l
tC49krGK9h8EsPpmYsBruglNltqcfTXN7kxABA2+Qn8DIX6sKowwujt52TMVKNnI9T2fucIctNZt
Wx4TGGg2QCNgiKnHocoOaDQBTGcnc0pTq8wbfG8vZ7yp+IJeFH/7AUh5giXXoVPhlIEUMwcssqpA
ShVCrkwJP7kqTSDH+9hy5M+fybI3gAs46MbLc58u0daaGSJRKk1hxXcc5z95Q/lge7wTtSstqymB
UOy+b+85oS2GxghHXMiv+y7y8xTrR5k+wtrpOZrQR+wKW/57aW0SMqpP/CrhzOjFybURygJDxJ13
PuMBRWDomzCWUE0CAO1sMItooj+zSpFtkFCzAnzVMxRDf0pcPZQUYLEBJ2AQpJGgDogySqLEMaNo
1ga5YXrjVS/TyUm2fA2zut4/n8sT4knm6JPW9cmTa3O/xo2aAB9jt9ID/0ez/hNckakKmNqfmJUT
8Z9GSUTNVn9KfMMrnm13nFWGxJ7K72jCSHbZni1r56K9+j9eXBdqoqfR+yhptJM0t9S4xdSSCOGh
eJGYJ2OtOVV01MtClJ7c1mOeVBLGvxdn+ISp/1ugjHf4I3POvjbsxupTz4TlrvsBzPJ0YjSpW8km
9yiMvWiY2GeA/T46HHyw+zS0F0UhZo7PFVgYQNTV3YIIDCt0wHsZZLfeffyouvpiTF8Xh1nqo/RY
0zAo9C5if0LbH/tS8J2GxvjqE4wnmg3zxMMUiy0qPzE3Q5mAuqT4WaIBPkH/ffitIxkLPOGhiLMM
ZzE8NAaZlSwu/LaErBKeJzR4XzXcsGR4tQ2pGr1lzE8UOXL98B5p9xzl5cgywesn4aJ9yoLXUvvy
7KcOBRFxi4yZ9OFgjqW5Nj/GNL7zCQ9POq1jVzouXCIO0rXcFDD6bXZ8/NOsLr9rHaHGvdAOrsvu
rhMSCoz/dg7FKE3CGS2ndhJjM+CcwhF6vPh7ySnnyEXCcxi4y4kJXT3gw2+oZQCfVzMnVzoYOT1B
PrXvLIvvW2rsV7VBjoPCNsETf4U4ViSMg9uwzMDPTccw4HFlFSMECU/dBVApA3vOoLu02F0ZGhKY
BGOiK139yeAeOboVPuohtblesBBgOJGgfBAYQXHwEo8n3AmBkNEjP8TD7z1X4px254XhPhIcLUdn
v3RsIjC4akarobDK86kVFd5dUHt2db6bC1jm4K1dulJaE316EBbdHvGSGqh+ZE9oajAk4UbqD+do
Dn011NSP+izwPUVQlW4fwU2XSNSNZ0Tcw3rV6/SyHI206ui7EVtJLTuivCHnRMZw6R2mdf/Qom6e
H70wL9iXnPwqz2AG1Xt7NRoDeYMhHj2TMDdlagScvzC1JxC0qJ8L3zKQW1Of3E+QhvH+TuO+Pd4q
LIMzwfsObKyS/ORBePc1XHmqpPlbNLrqe2qyn5+mHT4iGAE21XgBVuH6MJhGQ7iSv1JAnorgBOuZ
FfnjIQtJr/odSOOGgRp0SAiSdGSWebWNZWgfC5q73goqYpKqPSJgdPK1yh05K4CopgoArXwnbPC/
e0WuQfq0Ii1VEwFvax7u7ejGWFsiKYALU/UEkG5VHJ6TWWQjGRvs8WrmqVTF002mm/GjahCOCQjI
2Q5v62tCn6q2k2oFhM6CRMb+314xsnbfA89wnaWHd7ABnGbR34AvvELh6P+IcuJ5UpLXtPg33/QK
yxZ7vI6dvHG07xD0+wWTy04zigRGfOL7KJtel8dkgXf6qlLdzGuYtexlQUmGpGyR81U9ospg++i/
34Yf8Ot1BY9HahlMVq7G2IAiYI8tgpkIRJearLd0pAmnSQMH/Qo3eN2H1ryQfRtQ2elFkmTkWlxb
PEPeRTPjgcdYzj2cWMlzLIrVVSM+bBYgUKa3kWQ9pEu1muFL+jNw7WW6Qmw7oEdkfrL9IF7IoF3b
qgw1L28iZbZCNrjKwKt1Y97YZDL0Z1PbP9X4U/qvo9U+E/LmQV+LxkzfLuYejNlP8jTXz3MLsG3y
N54W25ELdaucGA8zmwB3wW77g70hRBpBQQ7KL6wKLOByN+OqvoO1cmyXPOr8pv+gB2ntZtN2TJtg
jNqeV37emjg0mjqN/7g7b5s3ksEM1j3jzMBobVndfqvMmimoXFhFevdTkfOsdbvbj0pyh72nOLI9
+FLzqcmSyZ3/tEnCqIFETonQ8q002LWmlLAfgpn7iOUGIFy/KyDAt3VIoR/NSdrLPMnbqOlIr8vo
K0hiOk4T4SZa3JnBRgWkUgAJIK0ic4nSFxfYrfaosYdSaBkYMFI4W/cyz5RwheAyJCSwCPE8XWfw
FlUdozRm4YEQb9/vG2dhQfP5dap6fFFUFTPQyL2w0EIvBKVKC+AwzHij4aYHBvaStoZg6qS1chRK
AvOXl10TLUXQxd/aGyVVRRm6nEa7kSCjYJgOfr8XUT0fio+V1XWitJqgzP1vJaMiAzx3N57Yxxwb
ZmEZ5CrP5ODJkhD+U4WFiz/0CiwT/6f2eSz1WyOXd0sS6AoXQsGZO11pOXFhArENRL78OaRLZNYc
cKNiSauipfA7al8eKxKC02I3xWWySOV9oyWTEtHobDdzAvvc1oqXDG5g9n8+UXw2AHW/krT0a8Aa
SXLzYcr4nb16TfeNhtDTRxaSnX0OaoBYxPSmDqDF5TWWSGwE+DiBl9pHEReZ41r4OiWZV9TJyeGo
qtRibi1HUb2jdw8lcbMbLoqFfAhUS56umhUWoXHmIqQcT6Imlbc1BXD0IFEEsa2xjTbrPzBSx9rV
C6SDAziVagLAiSu9oB8ON6cd1fD1lhUKJacIEbiO4N7ILQDaG5EIQ2eae7r5S4H5deMTm1SOizcN
MJmxasnH0b8rSveTr+M26hDfgHnZlPjl35p8a34ipyE90qXhFkHFzBP2aS+Nr1/Oi3VZMpYS8M3t
BdN3XJbC+D2URmwln0MpqjelFU5fmhkKBYuHfwFAS+OnjNkuDRJB8j/pRjY9KK/OLtNutBQdNUOf
F3oGxQle//RxGOP3Kiwb2nrNGqHKatYeIuZfidS/gG8tAA/pUmBz+q2zjvuUXT3r7givsIdlzC42
CKJ49F5/gv1PwyMhmqpVSMrqrns9FKmVm4cPjIPaSpDJDt26B3qXTOdZxGsTILHtQpHOqhL3YBkm
RzT6wMKGTiyqXeo9BvhPdI7BASoLjP76PO/SDrDY9HN5jU1UD2xKZChcHSxKh1FxQNJZ1DPMga1l
L7m3Wmo0CQhYsgBFGJQDubDAVZBY0+ztoFfu1g5XTdW3PTEN+XNtLDk30swFH/mXmPN5CVwdTK9i
Z1ItzgfakAIA0QTqbLT6oaBBfGujuHbhQjapGcAHXf4pJwgp0Z00Nu84PhUMgtLrQaVOByfaLglo
PIuro6XEVXdLeka/b98v/S3b5hUxDVL/cqk+KfX8v8cNTagrTaLfVzcNH8PdLk5zxMARseBBaFGp
XcZDW/phIqMHu5BhQlbWx2F3lFecMEH90uBHTYlPl4YVftAI2Y57+mW0C7KkrFXVpPCHQYa4h3J2
g/K2ZkEKqdz5woM6i6ALCd7+S2ZbbfD5gvKYZhuJ7q1NrTO3V5GvBG/oLRojkH6ieiapfs3YtHry
IE1QiMmNiTqx3JWAuKc5CoSJmU4wq+6PNNHsMeimtdrJQd2usgKPjo3ShjGinHYx+rdgGZYy8M8h
r/Y752eso0YaL6dHPnKJv5mhLUYaHS3gCHXjE88U00FnRspHsiZ9jOeCxAazCrR3njJX6Hk28V7g
EC6FjTsURkWD0eldpz+4PGUSKL7I3+jzQQiNK2nc6f/yfUfkaY89aIiuTu8GiMj6NAHK0CZsFW5P
MOgxy4s4dzpcN2rdYuOfkdtIYU3OEuSIRA1DdcTnngOsFr9I46+FRerDs71CgSSC+9mclmebkO7m
jutuIzac/ofr5xz8K7ViYEHwcKJs15ifsSAJhgUEpQoJPJtFMtn9ThsISn7gsXHsOAgFXOTL5Jrd
l9d+N5VgOXWmx/R5F9Pr7Z044ktNh0xFJrLESmB//MI4aLxwHyzL9e8rhRo0N8oW4YBDZocb+yON
63/gLh2BtQ22V76z+JWvWkCLAFBK15p2DqqZsevLHZiav14qTLJQqldcbv4e+JN0qGXVf2OLSe51
siCKAAw13nvZGtNnQ4BQcNSNfYoo3VSXy0XM7Qwc3L2BQ+blv0cZfykZeocF0CvQB7YmOwdm05zS
njmuwuroZKcVIP5kcEKoQeKZL1eZQo4s8j43gPaPYA7fuIn/OUz1sbVK2WvTT20vfS6rXALIy495
+94ckEmTLUhWthwtjNikkKQTM1UTuyqTtuBXp+LR5wbKSbqiUijSanOeyf9D3dwae6TnslEunitL
fpEg5SPAtALRT/CbYdDLNRIZhDehKR8nsrCQRIbP18PnhUHXwmMzw39XiLkKjjBZvh3k+Cz2N/FV
jmY+6Y0tjEWxWPHvUemTzalReM+lx1M/j1AOmqRX4sRfwocroq5AV8K2DjmUC8cGCe1TWvsWbUvO
xGMhyBy9sMgc+lKE8np7r3skhLHTA1VfLapKNVXJH6npSxpbrhFtEwbDLCEf74FHs/jPlRpKAtii
LejKrfGr1XG8WeoZmcvwvhz7af8rvd6fM5oe4GgRcGqnavdEs+SPItLriUxFYrlOHW2sy9NfZcnp
k4Ppov0AjmlheK47uJtrUAV0JqFAxia7zYslnYSs8ACIHPskURoDacvL4r+wYQZLM3Rse9ZD8ToV
nq2JcYAHbBo0xjY0JwceiKfbqw6qDSj00Lc6MZ5sMeGs+deEzNMny4XKRq8r6U2WX/xEJBWSL6Pu
vvtLqM0aiPDQAF3p5tT/hdNPIqBYcsKqPDpCbl292yimDSoKLSFszYiCwvaCLwtgI/mdOi19O37v
Rs9PvtfB0zxiUnX2XRb+x8XMunbvqbuNfKefAzYX3FntI6muppjsznJn2R0l+aJ9vLLUzGK3KExU
UIsV143ub/o35KGZjyWVjVo/g0V6btJ6N4USdnUUqJV51bCKsFPpUTtIN4YSGEBfmBcTnDDoA8RE
CUabtbYmnW8LbmOoMxgqVAchZ8dIPW3f9ZWN6itjZ8tu4H9RgbXkDV52tC8bcDiEjvNXlmDaaFB9
nSF6+/nyYB1hAQUajOi8nmwPA0bNTk3DsFw9rNzn0UU+5MSPizhid60X1ORetlZHO1+S/bvG3eBK
JtH6yEN8S1ShBeJRwXwAppvE51wndjZGGDssUUVTacKWZkC6J7Yb/i1nzPyUzFof9sgCu6i8CU4p
F8wa6oAyIlFwIoNWui/4/tGmiyqNd1rTvlE0h4UhFCDQfrmWfoG7X0Awa8HYdF84XrS2PEDnmuXV
46T7OvCfRqXFpVKV20SHgGFdQIp8GfbuTeOzeT3M7oFfMIaCzhO/Rezjr9n/shWRk5VRV7dfB0+Q
Mr1ACQknkLgUgsMW8uIjsPpe+JBTSpoB1Un8AQJxpL957NIAeYZ8Jf79bRkuVSoYIi6PZXdgdRgL
WrcVA7ebbKY74AvVZjloSJE518tS2IgRx9ZmlgLJomQzMlwuAmPzy2vvIZMgqypT07z9z/beRZFk
i96KIjrJvUsMKiqE/N/yo8n1cSLOMNDLsdVy+74SZcEAV7g6WKGVRoUYPuG7/zGtAeEFpMeTO9IW
TStYsr2rsRLj8Nr+/SxiM0Mw6EQcEQiPZll8UTq+E2WXTRUPf5Proj6i2OVBTjH2dfpxnb1ARa12
9OH7BkyYXUMoKrjIbopESO7J4srLyJ+wa1814e1X4Uqe652GNMpOtEjTTHZog01E4QtChsocn8Vj
PiV2600kNxIjsg2NbdsfZ/mkHmyULsRQWMzWA7/K31dM/uzIe1erpR2Q9hijVWYjGiSbbMLVh30g
dWjYCAHWQkn6hWT/emGoS1l7b661pxDnfrhrTRYkZnb2kydq3TD36wZfdW5veB3vNgeU2NfLjAjF
7aWer2o58hTbAchGQWShDzNyekklJSBz3TnDKOIVtcvZbQLEUL8Ygdybpf5Jm7TQwQedS7nqpnKH
1z34ywrmwip21xKfQTiP5nHTyeJbYSsXRQnG4qxd2nUBYQxORBW62eEM6of2iUAKKX7FeS0yhvm4
maKE/BDRgHprGxQnGUMk3G/yfhFM/iN/e85xSN9y93EBJTz+O7RwermBJDKOoAp1LOzd38b/h4OA
M+ksLAmfJvtmrsLHSQD+rIeuMM78OePuG57QsKfcNm/Y/D3ZapumfWix2zviNEnVvPJJ3CFb9kdf
IlSqawFxWIGsf6jgkPsvesrvzfVKoi/H3ehqgmXX3UqZVGRPZFPZKi5MLXdAUHEkrXF2oFaAgn5f
cbDO0/LBAo5KHpTWcowp9gdho2CkegIlXIHwyMC9B9yvjmlW/6NkqgBxLpvWKqR3yUjYr2UtEmd4
hIzcbp9HvjNKXXI4Nw+Xf67bbEDekiaagnUgdOMuLmR7s19m/1ukKphzoXyOF8UE1HtIkwOXRAdi
X4j543q6RGS/x/TNiA6y0kyxEABO9MwdejQyjrrb/P6yW3xnB1gaiXGQbP28yMRhdGDdRisj0Wmq
KIKTYGcmnDrDPjGE2A7mMOeOGiN0gjc5nVX4KO/3ktzSs0RHVkAlX/Y1tqp+unA6z5A89LVFW5T1
n4+lW2AinFZ39zw6DF/nz8IfPgGAnFHw7yGUvWUW/WE6EUPQP/xROi9YwMR0EhSoIEn/j7nDQMqo
kbZJwH3dB3mbqdhKx7sVI6cdIlFfonJXS/7bMrBKK+bkThgpAxmcsri4aheF1j00AssKtbtD1UZ9
/17J/s9R+0tZuzmMBDHrlD7Z6t08PD73xCPhM4u+qoGpVvyUIgZSzmdl4uyYzamm7KgmM+JQswov
BqBKzbFQpgy5lF+MUp5w/Csi++w8rZLKu8Oqlb1bc8l3jCA8hlL6GjcymTkyrFr10fBWkdTw807f
14heKsd7xwSf7wObBakRGtxA2yYNHUOol4M2ecDV1ECv7arsI+TJ35X85G0jbllVFN99+vYpiz3E
3obqnqZJFhNQKJ7lSuh+K4axqOSTVZHb92Yb8SzbFylwaMcuHywDW4VwM9rrwgInbj7Crqfx0SJ8
KgkqXcJbRsrj4yCujiTcQzkbnCjQLjx9GofH8GnQ6gKXYfz0MMNYt187Q5Bn5ZDAq29Gbg8HNp9r
im9WvhMiZN3ttoj4zEL5BVcBMfEN7wmFZwsZblq+nfq0zbbv0XkzpBT/e+Y3+lxVBniWQcN6yF20
cc/nnfSkLxXK1XAW9XljjxRHaCqrBW4v5KP45iGQBMS1Y6ZWyLU53zV4G0pQzXoT8cN+FpAxKZof
a8ORhG3CKgU7F0exk3+3oSBZo6bNy8ArZ+6cCFwCwmsNIhkf60JQfXrKBNQr/sGz+AOobYgVRx8M
OiciWE+eqyzGrGFi/bLhIeZA36J1AhibzhtsAhhCiS4+CJtn/kEFl4qbiucsR5QenE89GHAvfE2d
iY1ORioDYp+O5rVtvqj7tPJh9z6i4P5RU8FRsF/busVz7mW0sqpg0DCDPb/4Qur7cO5K8wKtKf8O
GbUnyzPafZKCaKttquW/lmtK0+X4v29upOy9ZyumFGGeXlv/uftE/yI10LlQtrjX/fk3TH/uBP27
8UFJHUbLpksjE4MWXhW9ftn3q7Vcv1Z0r4feK7Tix/V7EU35V9DjV+R0W6ocyT5qrDZmUZ5Mn6aL
KhvArKuJmy+R5Nb4i97WkQq8DFHKgsZTIixHvAd5RLFStrvYW9PHhlLbTvsEOxCT9hPSiCZvf6id
6osflonsqzCNTt1rrpGonz/QeVBU7x5f6E9jf/azeQRBKQulJouj1f8Ab9X2MOQhxyPHP61qc5h5
PdpJt1a5mJSSsz4ZVewgXUYSLg1lbmqMjyYjMm5C/5KM7SYDpE2CDL7cHwVlfe0cZfj8T9Za1CHF
d1sWO0beFDKKkX2+VEr4aOShQUmLYsEgIWC/2jH2k1QuVcxc6ges8XF3qDcGL7ePSnqHXDYvjwOT
t3Q5PQgpJvPgKIUFwo7VYe97KGydXC2PyIbGO0m1AinkNcddbqO6ZJFgsWgzI+zgsHnLbb++iNRs
LwhRBY4puHad2oY62Fg/grrvCoWwkhejlcQ7O8Y1d8MwhnVaXMf94Cl9ztawWw2cC0dCRIFsTOQ+
204dXV3CWMb0Xvl846610/Kem6Ket2IekaUi6/QiSXeACVFBRCcRiLxV7KecyH44yzLE4vFzKJwF
Cpdl9Gmo+Gj3sfTjIZ9YRvgMjFVhOjxXLIZq1kiWkOStHy9T4r0D7CH2Egb5wGOb4d1RlCbIz7h0
6sWJPeHakv9OhkhJ/yglcUaSqjTpDnV36ehsvEBy3y37G9wzMe8r6YAxiKYFf4SdhhtS2R90M2+A
rYtl2Yc6CZ3NjW9jI5CegO6FVL7+ke66/6pbSQsy7TYavL9ZFBoHO7Joj/zHQQHd54uXPZaq4kpv
d3yfJCH5jwZLs9BvfRTwAa/y7KkmQJYhPfC3gs0AhM8KPBZvUOUOOjLcRQHTrj3LpkhDmB0MslV7
hc6yX4tExdMOw9IbFGAwromaKrKruK8Nqbxi1FjDHVqDV0Mkq8mAoutaV0BpR/nO4FnOLRCCUBLZ
3Cq4M3/QS6DHGUhavb3W/frijbvWpDSjHBHA7m02X6w8iqv3lploIQeb0SncUn+MGLE7AzWUZ+jy
63SUvxZTIw2cS8tTB1wSComF2qpAA6B/ydqFj9RrN05ziqRBIphZhON9nCQSciFBNQxfQMN3Kebh
r1J7CX6T5Re/68yDzEkD97TWlznD7waWsNKn+/uygRUBAo3amVDA8VvCxQZIf0EQZCtH/xx4Kp5h
HOJaFhFvxG0NajKKMzv9tfV5WzMl9heo+vA3zz6+kLcJ0Sr9eetc//VtxGcujmZkGzyG9HHgI0hM
w1nsrkclACBcoJwOJHdPoHOiZn22Bdx5V2F0DhBur4D2uIhXgijUS+36cwmCcRVWZx5f6iLRT+dm
q2GUUETnxeXjmUrO/yp7bgshargimVHDkPVCDr39pqjInryFUOv0J+p62d7q2BVD67+A6Pp1ZSYL
ntOgLhESHoOMbf0mwL4RqF92f1IlbqjB87mCy3LTG9Ti7R7CJfO0FtXt23kYt5ZjbOVBBFuQi0TU
FcwN1XKDkGkGstoHhc3s4gYxoBw3aJskKoc6V31c0G6aK41j3T7nnWmvUwBafHhJ3nzTTmM+Kmhc
QdCIwZO6c2MAET/k0OuDSua2xvu9Ko8u4hpbJMei5rW//YEzHWJmNknh1bckI75b/grJrUKxBE6/
7BMg1TPGORzRuMlFK2H1ph/M505SOKkR6Ume+xjBRFpMAE+zMtzQYPlI8wmUS7j3xiYI5C/do95V
s4cnFqAyJuK7gK4AaMvigHTb3N2+WY+l8RGLA9LwORfTYKljqmv17MVbp/ZOkuhVp5F9sBQ+luKT
UNrKKK1wPmr5+Y64FmCib25YNuInt5UvVHPl9KGLqla5Z5N0uDanLwM/ea/cOc9wuZSQqV3QIvTX
I3e+Qi6CxJwOmGb9NZptDWJzViVt7UZU1amZxpXuIbKDFtN+H1Q2MS3G+8WwFfy5v2Atee9efBh1
64p1SCshe4//jmnaAoyLRYyE2rMcNG6UbJFyObxgo+5IXmTBkdrvGet/wkgYeo+k9HhpaRtji11r
t70EVFzfHHj3+Uuzx0rWinMz/8GlQH16PfmOwm6y+zrQA3pFX5WkEvMyNzo0K2AlsUCf4UTZ3QCp
pWBJbbsBE0IT2Wj0F8gb0qz9aQboBXGC0bepK7tvkK0ptUx9nQfn1sgXa9BcdBySwsY7IFPRdsMc
rSvT/Dwcg9m83flC+BdMCN1zYLrR6b0AMxK7LPClYWc7hR+mVkxkaOQFSKl3DuMunuWorxE1I22n
fpJzKi+ViPOn40NBBsvHLl/2IVRSuOBCPbMiO6Pjhn2ou6VBiDOKhXQSntO9fYwySSdAm/aQ8Klk
uMKoMoM7s7K8dS2SruYWWML3WBz1oDhEHy2BhzvWMLandzxf/IGfojVGMYmckBjcgZQxu/bbBNsF
mGwa+iq/rplivliNEyOyoJxpPAI61MwqgmfztvlWv2m4LffrLdYPt7RMpwAa+HDMyQme9oRibKcN
rKgL4bTfySoMywRsruaqEm7OlSFIshRYUAyTf2Ln5s4GAqSvb48RHFOzK04wnYFwXgYZYxwHDqCY
4fWYMxJqQaDcUXhil1AZlycTzzNe8hqCo21a6c0hZAKMjLFCNOZNn0ESsU1BxqrMpp/dsk77vme7
LLoZGpnYc1w9kHKsQBJsjDWhfciGH4IQlm2Q+LSc55yr8COFYRsAwEqusi098fb3fucIOvrdewjp
gDYq7t1y89SpQYQTj+KMgDaNuxIQLpKCTXR6VePDyBFfmQdPM3+PL0tjKLABuEhW7dOOJSkc+z4x
Wvt6N/XR5fPK5wn+ev2TYDv9QxBmWXxwg3gTRJU43tHKyylYa7thW44Q1LeLzq85ilGpJJHSJ2M4
ru7CrGDn8pY3moOEim3P3Fxo8X6jKT5giGMjEa7HnDO8faLBg3nwkJsd8OP4wUcQ/OUv4ZKgnuGB
rWspiqUHYv9d+G/0Tjh5k4ciyEGDah8ZEKa3td76OiPnxcHHQsNobvr+wTjvIm/qPVjgTJ8c0P/5
JwDq77uOyu7oHw5GTV/wliJzZ6jdshPwUodbJbtW946h56WNFbmlFkIF/7JRh1Ew4bphdMmeUhHO
iZTG+bIQzuH04OX4ABSf+UBZp6GdtUEIGkJ0mRaVBsVLPdiTwZynLP1y2Sbuk7vOTOLYU0MaGD6i
OUjU48yj6s0Xyk2W0E26P4RW+62TL27NTHsI6jLL2DV8SoLWK0k4J+5UmHZckUvbndO4SMkJoV30
pi3gvuWID9IdQIqyWRDIOGESDXkx1mrX4yG/GzudpsYZh6zezdfDxuLzpUI2NCvi9ZxrgkaijIXR
agVel2/kUiynbB/D9FFcuuz5CU3G9RB5qCowpP6L5lGNjREuaBfKpk5jRZbp9v5QoCHoXwpf2qHp
FhRSfF8LJLqeBEl9a3Kj1x9Sxls+IdselKAVUTabTEP1riWB0NMZnA6DnwvE1a5NP3SySsUSTN4a
yH8A9J9Tw7tF+HtqWVkJPPALH4f0Wy/Pu2opdc3f5jgixPgJR7WT5a9YLzjuWZ/cJtUsApIuH61I
Ozn+TAM03hVzR+3tUNSiYMz7kk9m0EHr8trJUi2wNeHT+GWdisZBsIwB/5vFH0kKg7o+i8z1GLQK
HDxGK4Xltg/UwH3WDT3OzldUBCD/wO6y/dayTJIxYmBJEUrOt+DRpiG5T6N0JNjPe2IX3yYOs9wl
2icRltlYsbkI22ZZ/1P1T5Rpt3WcFqrgcnCBJMXKKyIIio3zq0oj492gFovHfP05a507DzpGOHv4
VVYFAq5BgvMeKQ3ZiVnZtRKa2Nf+ojhETcdEh9DjWj5p5W/BVSAddrqkrUswbWY24jiTMJkyrj2D
Og+2jxtSs4f4mIQo4F12rtphHV+Bk2nfnpsOUF4p0qOoVwicojNXZMMObn5HjViPq2o6o0aFFD5m
lNLcQAYkpUhpMNUSnONC/7wci2StJ0YRKx3uFEZZQhRx7J8Ze9jxUYah4br2yfjrV7SgsAtNfWOO
ewTwmocYWv90VeIxjIrUHxdExccCBkTC0z0KJvwUE1J8OlPjkY0SfcMpG8gr0FwylQq4nd03bRv3
ErYXHkEaAoSUUUKit/xTJEouLc51r/ltNXKAODK6GdLlyQ0Y3tYyjoeOhD+7ifl5gabGa7ZuY5Ej
4NMceJTIm9kQ7q1b+p8bli5nMZEUDWi2nlLgYPPew+bXYHSESlibGr5muEek2bLx2wOeb/mgy8+z
f6yMqd99nXlM/ai2VRJAtXFGiDhA1fQfhT2qvX+iCjahQ1GedUEjCF3B7xkEaikWkRlxkfVHI6Gb
MQoGSJdx8V12eNBDccq4DGG6YD1Zsc6jxwFo28WkEGH2GZhVkpLW3VOdacly36kKH0kv62o2iMPK
T1WQMXvcKIVFQVY+ObGXd1TxHF3xITKXrRtJBjGNmXXXSe1rSIVvPqjla2wbcp+VclJe5KnhGvBd
Wi007if+iglm57CMdSoLnAnCS+G0PScUv7VFkTQR2ywzyDYcqWouc03/QLKFsvVSDZ/o48/G7LYP
Ryf+TqJJ0XUFyzGYKDPHZjZu0ulTG65aImaF12wZcm7DrgpWOWY6VhOe7u3k+//xbAvYkQ9115ar
W3qiMws//M/ubY/Hlq+C2zjPdpY3XrFY4udXyU0ztdMmYIGFiqLrI46hQ1pkWpUyBsrFEMb4ecmi
WHk8TZgjYv45i9SuaguCZQFtv8MY08TjZTzYkQiOKd3aYmWzaLqtnF1nwW0io0mGboVklHB2HWoV
yJ4eDUgFq1438lmHbf/9nyHnfJQkFov3rby1rAQsyCcO9rYevqlmPNTza459PIX8KwrQ+odkcf1N
pCDViOAH4pJrwBe5KTHaKajLNB1f2v2tc0k02coJER0siV+483rDsRZuyf3E2YYUtnDH3kot8+PV
oJ5/CjAwCr5laenjNfsF2XSaXFSj32tFezqFCxlw46iRipDGizcODTjhDKzliuE58nASnZntNAGi
DsNucNLMICOCNR1PF3igDU/oKjSR/h4Wj6sEnlti17wpEG5CPXdtLXU5GTRxTWHlz8R5/OpId5WK
i+oRGDS4x5BEvPDVKVXbmbuxETAw0FL8a7gCYc3QJKZp9vP3/4qbH1Qc1Q7eTpS9CkH/Zb5AhHLy
pX+JqG+WeayPZKWK1SAhiO7YwT0yHx6t6ZSBbcgfMrLUFnWgC+wLGHLQmpfGzXLkdlHkiVrmnnah
plAyyknksp1hzM5X4PYYjuR24P5X21TqchuOr2RuGHQ7Y4ETAsIxPfGoL8vm5wdOROTmvbyNyk3v
qQtEUPj4jNspY64fsI++KYZLDwAWjmRQo01cJwoiPtKUmYjhhTOOXpa5s+EUvi6Q2QJPR+EzgYmw
oEYsCTBcwB/aQgnhkfjrRM+a79njq65bnuh3j01bV/slE2HYkSfCR9+kYfl4+RgTADrve3rRmIf8
dYGSZq/8uGlQVgbP25qAishw49DwQppKq6QweU9Tm95VXLLRUxfmvqqkv0Rgz4LCQUVUk0YuQaO6
d57P8+FnR+KD0YTDpeAjeAMiE0Rqtq0LXDnajAYPY0rhgzsLhoHF4gBynpHX+qPq1E9zGHOJ2Jgh
LA6ZuQhC3Zv9YtnAJdag6bg5s7i9JIbwCl7HIYRb6h54lQtGx4hnOYwJAk/5GJpMtsm8z68zAzhb
mcjM0pyKwRJokwvsX+pXnFoJMVxJ6Ft7VhWzOVMVbHNVNDS6JxeXJYkBpeePVJaI0Or6qTHD5wPt
1op5VmVitEuHEGTI1UUA4UXrmPkb+h29xT95+xjR2JuwSWvgU9dol6VixS0yRwvO5Q/liMl2V8ZA
/oR8Qu/yLGvo/4bdC85C5VnIynhPsWcsCAc1WDPa/+IZ9tE5Uv44zMUfrOS6SERIZq/k8HywytWz
v8EDrf5ZpRfA2z98CeKyiRuSDZm9EsfnLjf+ZUu47ortt/vb35mdSPVg3BWpMESnw48brVDdxMwE
4j71oj/yO9XlW/lVsgGPQoExS9oWtK6f0PmRtpb17WmCZKlocmFnWOZytfJKKM/CljHU1EL5KlNL
HsYmcAwPQwsrf+Oehg20TiSZiIRhByZzy1ASOw1m6x6j53+rWPCjAYuqtFFRz2vdfbUs0mZDSFbM
nO3tKHE+w5WIIQTtMIu971/0YjH3hx1ybLv3+t71v/J4GYXowWcbEUBgQv/8XDncrwe1nTlSkoxf
Mz32criBNq/6JwOBAg5bAZFQcpL+DtThgs6s1obxutOzSAvDUSqFHuLyCxkFerArYuA1xyVSH/Ix
TfCZmJ9u3zhiPV+xguebkE8c0Cfvq9V6T+G4dv/dXTI63xq+rBNwLMj2HTN+3ISLHShvQbA9v1bm
TjJEWQFJyYpPJEL7qyEEHqBnhpHxc1sngrTlgh8j2KeUKRthhrINyNdp5Dki+3Pm1zsMI5JHtsQG
ZMl6KIGJFy9wiOsHWntoelri7pMX0EBnEb9eGZSdxSeHa83DFsQcGMrpCk7WM6U/jojIl/+IO3Ps
684qp/cV3NwOGRs5VdF2vQpE7LyNWDLxlgc5JxhYBz/tG04Kw10UR/OUjV0wFHYLeJf6AvzQ3zub
bUsQ7eS3dB6LA3trK7vcvVEKntHZqRtFSZyhNoGRq2c7HJtwCQllnLhygOEFptbz7kThb0pzTXIM
qfb4WL7rjwGVsxsapsz+5eaNCpce3d053lEdW0hUWgyk86I+boYxRcJtXjvUv3PAE2aXrKZLTPcC
mv0LKf7U3kosnHq0POxfrm+deQ/alzR9tUqY/wW2HhRfXLvsHLDtPIopXvrDB0fNBKQ2lYF2OdIf
ZqnNK4KxM6GbpcgXIdN9yUhe74pTdG44g/r4EOMXq4LFsRIke60di/A4Yalu+6fK1++2zqGlX5Hq
p8UnxN8A0xGebll8jdbSyeTCXmJII/rMs1SgG6mz5+2lEWvysaQMoJXOypAcnpRUmcvKa3NB4w9v
OXSr7E7CyKZBtMR97E1Q61V4OBxRmZ+9eZ+9VDi2UjlsC+r9BrY9C+SOl6DOed45tOcRTpjGLgm9
R3Kd1ddGjvbeFd48ltAQN5mL8/1IQFGnle2PwGOvmChzxcRfVEWFAW8o3sO2J7mBeFFAiXScDrUF
oZSS1FhZB/nawIZ7tkulRs591lnrgGX1vZcRm+vPvnAaUloUmNXQHliZLaGkHvaLGQEPyGNe+dnK
FFp1JeFVeXFca5RP/TvN6wxlKJKzN+9we3i0naJPa1WMn9YFV6+g0OfT4yh4SrbPZ40jkYADRwhS
Z9UhdLn7eFD0rJWp2DL6x4jSrvLF+nNCfyKpbMEOP9QoVjEYN5hE89qJ5A4bSptHO4sP/SJblNtP
2yP+FIGl6LyQeUMt2J383/cS9wZSxSGFGsU2nTDOKFVzIMpV0D1qwhBYC50T81A/D5jQqQi0lrnZ
CW17Wt5I0wZGqyTm+TdJSywpku4KhWQKwilXmTCgDtev2BQwD0y/dsM2uQri6fgMSsx8KEOHKZ5x
zTdQhR0lLZO1G3NV2t1Qrcqreiuo88P+IkQwTQ4Bpv4zhzJWu4LtiVmjNVFv6FvP/LmxGgr2EXA8
b61osb/UE+Nkb4dsbvrOByjHYl/M5yXj0oLZQ7csiPmytTyYtfI8lDKHhx1Ic2g+pNO+ubDgBUmR
+j03fKrND4AzBwi4b8gkE4TF6natGqbl9b82T+krDecdoJIR5ifWD5zQaofEyeuSeFQ4DAaXMbZe
xC4N7u4zEgBu3XQ91XsdKPDdZH2tUI0IazOUZQ0SwNaDm1wlAAcXU1jAYNW9vyc/SvOjdwN6JxD/
h+HYHB5/4ob9bT97UddtX4q8SEwprlVOVwBcqAhMJJ3zTWEsXXiJlWZabJpiAewr/LGhwJW0Nh8J
1a8BJQvgLQACrUGa9+mLJwlM49x+C2rfH4kbeggInYBXBTSNQSlNKFofP5ItB0hNjGa0qVoUJOsH
ZCyXR4hFhx7zV5XthQrRW0NQjV8ZUyFVsMtz4iDT8rgmT3hHKMEFn4Zj393pMyHXpceu/hnSBDx6
gHtLeiyikLnmSMI1+9rDXjk+qO9dhsuKgr1waEvGzIRtWhfL1JvBI9WCvqXULlCBqeRmC4OGA4Ju
PveOgoqeTpFdhfM9MUjr13ix+ucx6OBtdvfWkPkaVth+vXMhIk98ayU++oiYHhFs/aZR2qSXmreZ
JQjpz9/SzzczhWLZTLhzCGGwGN0ak/tstTBMdX1tyxNhZAbodnnuNbKiWrhRDa699iJ5QO/2iYwg
UU+0ph+cocTs0ZAxubQuMdUde20Uua2Uhh1JV7yGjmiJcM+jtZWEZK0wDBhBwV/lOZsXcKKzGNnY
HLVqmLtQ0Abgjv/MWj3ot/6P8ojsIkhsoIFOvms4DSt3Iew3OIQNVYaU68Ad483NBzSkxCl+7y9z
lBpB6RDmdVPcSSQMp5Cuog7LvnSdHJtU6UCqkbAH5N5iH/sSC8LErwja+ZjnJ+X/YNUQL8JuIUTJ
QvqlcKt/CI4daAnuqZvVg6HFsZXdfPegovNeH90okygjmnwQVi0W1I2OrqZCaSPYnwq5qmSnEJHZ
mJH07vJEyvApxj462KCMXdUe5IwReWekJoNLBekBm4D+kI0dHifPdJkqxqkMywY6K0OfGAe1alX7
EswtsdZy+fwLTu6OmnNRJFtaaBSa5Qd3oHR/J0QhEvGMdAVJUnYV1yJOLFOoZqjSx4wykrtEshrv
HYJU48MJDvrTA9t5XqK0P21Inf6l2J9bCFs6vmnhfyPpAUAkwuzjhbo1t+4vVU3GC1l27tV0Z/YH
uz8ionHfXZvzfwMQL+pv/oTg9IDANthfR7NK99rWTvfToiQ1aPAjQocbV7KZDsrXZ9VQj+afEugX
Skz5VaaAwdE1tlTy0TWgX/WSAtaARYnR4maZSBPsRr+L77XlwfLSw5j4nVWLHatn0UORBSDBmtXm
T43qQjGR2JvPhe3W0yKsE0ot80VgKT3cwE4mdaGIY6H748rdQjwnYkDIxLdT3PLfrf28TBqVQBRo
/po9AlOvErAhty4wuv/bYHw1B4V2v15Zbulz2mClBd5BtCugQ85IAyft16a5KQJDfvyz1lHkR/0h
A5agaL3aaL5qOqTH9qx6D17PIB7wJqF++1CjU7w0R0T8mld26TnhEg2hdymLqNN1BEOQVNddrm4K
cfh8+g0SH+49OTzutE+z3Xqxt/CjcCu1QM7C8Rn2dHMupT5EbC4TRYPBBanwz9D3lOsyG9OqXXUw
ChLmrqU9LexhYr2F9/scmjr3e+nAYsURqoW/MkuH8cybJ3DOhN7+NBcmVWwFYclkr0LGWqa1bLxF
aAJN2ld1DDssIx/A2LSuRtw5B2oWqWx6K9++56kAzmH3E5iGCgSIc161NpeiKQOMGnyCQYtFOs+r
sPUK7U3DRJ+eVjNH3AoqQ3DQ+ogQ1GbHUPpMVWMeEHbb7daJxv400bgubNsh+Akos8pYqe+Gcaus
H6MITekSSkYpvgh5fGtkXM6FzSax7l+NwPNweEzfkMsizP4wHpdj4BMZ/kgBYs0BLmu/Fk3y0YRs
jXoxGqoDaPUcmaT7JiODRJE7KtWgHJB01+OW/9hdj0/Dny0Uj0XNbNNRvZ/8AyIlKs6w8KHQF/3t
l1zdq9pDQNiUhFZwk8CbllX97XYEY7WFlEd1map8N58NXr8kQxiPky4nCq+wGrncHidK/5NEQRaI
zivm3X0iMRM+duDwdDQldrUrNvyyQS6H4iVkmBozhKKnA+lwQ2YO5U2uRP/iFGg7wNWwaboxh0yv
UwReQwv/Hez5XVqSUmdQwrOlfjSmFMGMtcBVYMi0wllaue885wPaJI+kaZG7X4Z4AEJkU/Ou9PAL
bd4DLbFqDA0zEMdHnwn//5WpPS3N2GwvncVSL/u8eo6xhi3f2agfTFVKS6PQdk87qqBC7zfz6MF5
p8X0JFJjc3JnjVOYRBPj+gyWTLZBEJ4lS3fHtv8Hvdj/lHVAEKszgevnQa59SJlHTX1kxGM4RxQ9
4R2yUWN4MMa3/YaiXBKNgROba3tGzfhOEX3addYbPwIA61UEiZRvhbENJvkcJAkI+iLBcvNjpO7I
Vle7Id4jsBpek0558qzYaz1VvhEnh++6slqQ+E3pqb1QBY2ndBJCnHu1J5TW+z3Ql2QPmsy2vmZK
d/3NxXs9CdKlw1w9dWhscrLNqk5tptwhPfu/aSesAPv1KHl0V8PtVbqRdHh5ktdyNugijyPwpnwv
YM8uQhhkq9bk34TOT0piIn/F6ownVRFR06TCqvtmJmNXNWCARE6FXGZiDg0jAX/h3gy0MOvblCXD
4IV6HAOIZr64f58gY1+O6l02rzTv6pugiF6jOUwfqvueFwktG9utm0pZG/XtLJAIjXE5a3Nzqhlw
Tm3bzb2aJSOfTVZ+yu+jyTJ/tqlJKS1zE2ACq2v0cFfRgX1GTpFMKNwwf3y0hrSxHcZEPqDEjbA3
r48fAKDfqbU0fvUkHZ32u4Bpqk1d8K+sX7wAcrP8kWNxGECMlwi3NfqlwR44iioW4xCGGfDfxecq
WHYdEetn4ptmct1R92pyCZpNjxF0tMlnoNUpUHB7MGd2xGH9KuiBlG2LOTeiSmlKMMUaGkuJije+
Xj0nU/xKaFcfEdmAnNbA0NBvb0Jc8VRXUlWPBpltOlvWR2i5VgEhIgjhLB/QcSuHk/EuwX8LQ+Pr
IJ5X+W02oQUROscDXfMphaxodMgqsinAfSCKMJkfmnzlDZB5bJdt49UcA66lrz8yjQC6KIAsV7QH
PmbVPjr/sO9EY3Mdp1HNia5I71nNpDns3QvhNKSd6o8HGJ3wMRRcFqldZwRjw6VvvuzoNnimk2pf
PPKXE8Cw8uRjAxw665I6XZQ/2vg+DiUq0bZb5jvnuecZhSewPNpqPaJRJUREmfXHIPTYPnItDEb4
drIEO9F6BOca6TT8JcR18Ob5Uh+GigYQqMQAtX7/SE188Vmtks3lDWoU+xqYiYOmfAsEGqr1Ic66
EixPlI4gMM9q3FENWOE5fhYDO0HIVBtFOvixLwkNHX2UIW8AKC6yWi+P3ztD1gvBRpfxLkPfDiKD
ePg34xZEgBFFeWJoMB8iRwagQ6z96plz0qGzwy8WDqnlsxhzObey0tTmQVMNIbInA0zZskjD9YRp
apZ1RW+h9zBhHtb+A+y0fOoETlYqV4OLYWz/aAtJq8OKQb8YDM3DOMg20uhJ5efQGGMC6nWo76Ee
w3X4mNoJZ7GQVSwBCoDjoo5Ey5HXnZMRLXJkf5M9hpZG4qYKy1m/x44yBWJ/I9lX3rinF8W/FiiH
xMyGD2jr0qQk4X1jaQAzigfo4OlXJRJzn9nj/+ohMy5nDBPvtkJlSOE3206DJGJ9PjZxaGW8FBZn
rUiRTk/5cR6RBnFYiDrONM3UryVo8hDQfCmcO7jSm/mvcEAOA93zNwFEeAFHn2m3F9EpEbMcpNHF
DIDJn1DoyeLwfnENO14/w/QelP5R2dZJD2YdiMWGFPgUkChrj5sAdT7UPxs0TLf/ycrqF4rEEw6F
KdSN2Nnj0wvDfneuFq1xkOJzGgav+R+drBFnyZz3PgRutjQobX4RyK7oTqwo6sdPOzqYzl8rE4Ib
ppa35/QhcSiIwR4Mzgjw/xGfaYqVt6m/ApwHv14UHh/DNKfHIkavHxCxZDegL3bugmCaiCNhipPq
Mjf9FeV/EGQjECFGcVmnP2UCKsNk5uHah1dNL0MgjY4uA3mbXnN1x6t/EwSxUNdlZXHxjSnZoBmv
vuWD/xkGe7mXIU4RBgnJ2FyqtQPDQrhME4GmfmBE8oTw/j+T8xDMm4PTT6DHE+NAntp+XrxWhix+
Jie8NHSHB5No3uvtviM39nieMXMbMRs61lPMAbnUn1mNIhhnpc/a4n6KfWTGV2PZRQSQlpd1xrKc
SKB+qixKdKnjQE4zdq5V3IeguLOzcpPPMRvf4kmswqlXJM+AFXLDOiKYL6payjyHPzTSqyTQ7YmJ
6eUhhvnExUKUwxmRyiMZNRhjAAR2xer791p2YQSjAGmuF8/4bgEVn3WOoKoOoa7UJ9vuYTVcZ7o4
AVqEEiz9Qg62Xew3KMA3xXlPnW8rjJT4OR1CGM4aSjiJ3M6Zns3bXykdwgwAeDjmcLh6xEX/ICr3
ivrgqb6o7I9h5lrO0uCRL+TVWe8ouELfPQDuYEwSfpcrxqbzAFTL7KWL8EWBd7hOIYMMkuYbkC6R
DIU+p9rmlyiZgKHDhQAeqrMqBnKIqueRHXKuXTaYmdqx6dpFQvlTqoMGhmXm6qNbU672lmn6LpYj
dBUdF/zSIjjH2GiMre4MQOEoT3bghkcSyzhmMsj0l8ghdnFPyL2NmKrCgfoy+bblBYXepsEYiysW
x7nOPNMUSzMk31GIrMLEY8cTOgxjcnRHQ3VcsoLwD7/XhC7DMbr9tsuL7YnmmhHCnVu+89M+Ew2b
lJbucBf0zNj2Ikb1fdVJ1Jv4qXKqY5+jqmmD8dMzF9MhlCyUYU1rpGXpmSco2o7fL0puRJ59w5Od
2RhjT34oZgtUBkxpsvOHTb8AVfL/1kqVPzjYIpjtjQR/3W5CnwtZ7Hswyecm20vPQz53rZ4j07/W
PsHvSXG5gEfAY3tJoVwADHaStRKN3IG+e22zyZOXIdUW44t+HS8pXmLf7sSpCMhZ7pd6s3iYHdu8
m+vCfUFlMBryukwW3IDXGHHcNX7csMTui6ykDuIWZqGsU8i/IHoYt3iAhgAUsLCAPQ0iP3JmiFvX
qjdDO74Txg14DzQ7sFMc7JWKvN1tus3n2iJGMnFe/N9FkJqJPlpJJplfLAUTUzMO/Nm0ug161uwE
RVVOPWBHOECBOfm/fy3SlSC5rhuvpsuLuTVk2wHKc4+aJeSkbPsfKnFgzIqhavboXJYV271kJWdM
qRq4vV0QUN6YAuf+DZufrUoPD0+SIfpI0aO4tUN3j++dRzt22dBfkdQBqRYouYsh3tCo2QZlAtl7
iqlscFHfidppR+V6Od7cu5fg4trlCBdTKmfzcbOicQ7jK2HinlMVjPBKmRH1Zm9+mp6E+rriKzog
rZ3w3YZINQiJmgwG3ewZpK5NKWzXhE/4n+KZI3ScpAaNtKVlfwD3Z0PEA6CL779zIdv3kl6pZHnD
b+pKgTHAvIdnyW61cbiylc1lJEITdLmxvJChSZYNkC/P4+B9t9/xQMNwVURUHmdL9nLEWJPcgdb/
pY1vy5NexUum3EzUbJUOWUm6lZWIzjeRBgsfpL+YzaKIMBOAMkoYrwkdyAZQyy0aAyZphPI+NRYp
kaKKS8xaRen2wpQebWg3TIGVUgJA3Hk5xDHpyjiY3EpKokd4EAtCsmGwFp7dcnX0KGZKv2idg2W5
gx4clGPmYuzvTHAh+8/cOflcY0NqET/m15C91LAPAnmsN1pKkdOi5k322xugRAmg+qSGfHLi6vMF
qXPuKS9Dsc0ldJ1jfy0ZL7+19OoPyaPvE1bDPAl6lwhFB6Zh2YESKj1+sP9KMkJKYTQmdbFXGxfK
WTqToXdJKtgIRtb6nvPEurLRdJqdnh9jIvNBAT7oZjMwVFUQmF6JvJ/x2mxwKb72qjOYCNuQvwOO
Hlx2sdu71xyZLsgbknQcoeWlp9kCY0oRiHXaC1a2conacti4XhLMj8JkUICDxTHeilBxtp9Nklkb
ltRLBSn+KrYje621jjC/yFRQeTQ9QAsDcCd1WIudGf0r74uGYAaooWT/qLQYzbO8VJTGfVXkjDLR
uapWVSLKTiGxSLDua4DLvnCLxaxaxaNiCdhDL4MzQFuOH5Cb8u5db0FEb2bTYT5ZGARIb2hT3EaP
cPmixKm27tqp1CSPq3905GYA3eYYgyZy1ZI/KqzZG0wabx1Z8gYwc9RW3vkOi568WnSI5yeOTRJz
FOIWwNQMsuZ134PrmQL55Penr5TmmFZ9yF+TKPnGVyTee1XSxkuhjhxMLqRHWJYTrlLSf0N8v/3Y
pV5K+m6Ha7D+ehg2wo861gSpRil1jNaFVBjluPAsXphS2x9qELkgj2DISBYuPFZhXsIpLoXqG/jK
KWsuK2DLGQ9ev8Z4qg/PL45iU7CBqh+KiUdlVQ7JkDTHGrTv+2Z0UG44uVEIFiTlGoxZPf52urdD
0xcCphEylwZseYy5QqH7YgCAw6bty7fRq2ZLhmqB6cA/nzOHIh3V6iCvFnzsD6Q6OpZKJBvnkGY0
4txE7xkOjWkSJjZId0ms/Vj0R0dkHX11OQ9A8cVR8YeYecoW87k5LdnVRqu5yYPe2aFl4IiWYVeH
bA/SSFDkA0onAY2nMcWRrXaewZwxnxJ8a4uZ3z2K02iT1HJQ50FDsaODKEUbWn7ItfdierCp5P4L
kLsDI+JxWw6udPdlYeAXNCj9wuu23L89unjYD+T/nzoF9hvud3bLyIDhpsjPPq6KcRBAnVd3ozZE
njCHhxvOKj20rObQbzktefEovQ9HVP9Jk3D+OFWtIqQ0OydBJqh55enSel3WZDMe0SALDMe5D+qm
9Dv5DvJfwMt3ORbYt8HPapA5uDSZYqZm3d2BJ7bbWwELFYaOpx7xBQNaDEHBT5eNwxlXiPPMonmC
BKlbfbt2hjO3wknEAjr1nEXgzLVOiw/XFxvN/x4KNzOvhPv4vxxZQf+uepnxNLC0rtzSGBEgVjKc
CSnd5eCuFYldZIPz5S61xzJ989+/1kMx4Fk54jas6S0gcHvd//iqF/Fu7lW9pb/euJqDjQSgWZ/K
6m5IFDUfeAGeuQSR4gpq0Djjp1yXpKau2GSgG/lGT/BvS9gduKjaFA5VMhJa6NydVyHcvyM0JW2r
Rj+TI+96qOSITAoiJaf6q4Ppy2dF9Zt/y/avEiUfbksGUKsIWo0b9gnpnWyTWyGY6p1GKdjgOcyO
KZSXF5ttcrzi4lW/rPfIONb1v5/Xwd5bLfwtEU1yOat5aGG8CR9ziMGcsmYVv9va1pnd7gw9yIfr
TfxEQGlGhedVPcEI74MqZhoxcG/flM0NyxY9rfhww1EgXDIdcdf/1lTPJHo+ZR7hvITtwIU5yG7S
w1zYgzdhF6pthlKaHz0R48KUyZCpOwvC0DUyYSge2Sh9kVhJiMXO0GlzxiaR7X+cUTeijJXZNolM
J6qG/M9urhiC12NNbRyuCf3BmdhF7E3eedJn/X0lqbCMXJhZMtTi8zGIMrXn61QxCLFUDpL0CyPl
MLNtc8Dwm1QYEziFf1Gzeu8ZBjcxzeZqpfYXcFl4hoS9zJ4WJnfRBqcDBGGoqutOw9OyMG4uirrp
k637Im7TN6arAJ2jl0pMrZy1xP2wqIImcA7tTwgc+WzycsE8maipxf5cEw3lwfw93AnieVFGIlg/
fH5im6GZx1QtZZfC+JpFjQix4BQ3x63atMDYhdRRCdbTybyFMkqb0QZR3RxcD2E1EAsopplRCnbV
zIMBqTLErawInN4dqYcTl1NEh6DSYc9e0YJw8V6NAIDeKgLkCPE5j+SoWoi0czvku7Wu2ah3o6v8
LkcacHxHp+CoPiRn03jrrUx6QFX0oVi3tkcnjcBdixVu8mJl70L0O6kMlnXSD7QTdAb6Ym0RLL5o
ZmSSjhM6l+B4Pvx5mt8IuBK1V5mOet+uy3a6uQ3XvmNS3e8eY3NWy7Jw++dzH+4/u869GTsyvmGG
el+WcXglMS4v76oW1u+iN6unlQYuZ8/8n5d6AX9mioQlb0vrqJm5rby3hdlHA72LJRfMTYjlX6QD
dQNZSlQ4HbVALsh8AWh2hqcTshayFqfy67Y8vgYvmD1zVlMHE0eFy5zG0k6GEbWc/nNN0bvsiuII
TRKlOiR7d3gzhhBgerTRND8eBLZkUvawTHSMFH5/1f2oU0UCROOpJSsDTAVuwFFdsxSKE8URqAm3
uk7kt/eqyhdl27gS29vm8/ntflATBr85mDWNs09ElIbJwHpNo+dReHsBZyB7aUW64C5KBs0YOS2U
sGlBS7QYb50cmnEQUehF4VDz+4bt+XNl5YtP9fZJYDIzpPc/O0gE/SJ76/wpAmZ2YGcXDYxiFdjf
UVriWaqsYkskz048/tV6g6u52zdO7P4qDF7oEI0Xa7mxtmIe0wbOzqe+lNCoKrMZoXd8u6tI9Tcv
NusoVOgZqKinYSAuS9yKLj5P+F9fYYO61mnuaeVe7rLXp+IGcJS3qjSoI3sHIv235AtLAiRLjBwc
9e1jIlp9pmrfUDWS801jNa5+jcMXDmrqGBB4VvfFVtcXNlGSjTMT3QfsWNMkkqymmkuB6qyimG47
egna2bEFRZ//8Z8Sl6yd1YsoMj1frqsG0C4aaEndtfAdyjhWhS83dJgjikISJLJXo/aRJ7FL4q4z
vIPiOYOyLNJIooyvMockZFq+DwbTZVJKJlszs2XiX3WXAqidNkOb5bGJ+Z4FzMU7M9ctNWZ7QtFf
aR/j0n8mUdeaWl3IZmvVuc+fSr2kDXRADojkwHPYnraWJ8yUEJAiBN5/rciVEDsyZ0k5J0/fTmm9
JoZBi02VSAeF7FEm8am0GTzoDzGUzFmOO4v7tDdhX20+CX6VxSWIbJg04BTyak1a9C5z8T1pob8B
Jk52r8xc9aYzKMUmNZqoyHMIGke+m5bvl/yvNn3674KQ2UyTPMrY5Be5BzvVyFU8oTwd4STMVsyx
CfE8EcqX7ZqX0SUODePyjRBIHYqgZYfKkerHFE3184D0U5deqgzzvS96tMPOU5pWgVVUM/BXavJ0
R06fh7ct+vshnJE2tAV551PIVL/HPl5C+EjI5XDurXsIfOCw46tN9UwD1em7zfcnm3iCY4u/HsMm
PtqdkyqcmUHcmXdvadEBUQoaQDzIbWsKk6GJHhqzXLWGbzpNY7G8lSvwCArElbk5lKI9BfpSkmYp
ofg5Uk2u3kgskb1JNMOTUGQtmxHr+XShqbpYOE1yiHe0VWlqf7B9kOpOltjTx51P//jG6f3FlTbQ
2S36PbaRRCmxU/vkToxWVJmU2RQy4YGPwAv0KS7k2rwp11iZ0YV3wQPpFlFW6kLeaDGc3c+b0QVF
OVL/sI+flFGlySCzzOgpSfDarpPvvJUWDsUYgbJUdbTZhe1+0W96kWK3qmp7cllKWJNOdgL3jNBx
oOzjuEvjIkbopc3nCxwxsQUrhLhh61M8EFov1qipghcw3nDA149gMFPzzPiR6fqYWRpagDmGmTUv
Rdz8+xyfnBsBtijiqcNs3TrS9GxJOYqu+1K1H8ZXr8DB3adfjNsJkvFlcb3+AVDqIUjcR1aIbOhw
P39gm/NwUDZj38IpdWnDf6A9fhKMx7dqfLCdsJUxBbVUORnkPbWtv6PmcLpODZoL5C7DzMb3kDwz
qX/zkr/6mYs/YxHp+mu/QuJ3KNK7Fdiz8PPp2Tl3+iJnRQBOpMouvEfCCTQ7jDQCZ7DrLQPKC7eZ
6eImaey3kluh31gH9SRnNnh9Ti0FKSzN9SYyRK/KhcxBf5IkwVgydaN9Uin6zBN/ugMGRwfc/TJ7
5zqD4QJYPVTOl7O60vRKgHHkrye2JzWJL/JiWPjmDAWAQrWvJ9aiyYM6RBBsOxNjhT3UJhrxzkfS
6eQQgKfDuoaR2MFNYHAUP75fNHXNjy/3IAH7g7v7KnmyyR6g7yJkXxhiMwe0EuZ1XLzgsM/v/81f
LZNUkZdZn9b0XA+raXlwV8T0CDEuJ0HX4xVD8T8iIf3ntSqxYZvgIiYJMRRv0eu2hA5kcKHw2eqC
gDGgfNAiiyK2gteMzT4A2aDkDNYrCB20jif/Nf1LNxDd393DlKEcjgoGZgtH5YOMceW+78s3a/5H
4UPD786RXfnE8/Awf+gE7cqpgsC4CZ2gTlwlGMyEfeQDxIDFPWYrYL2pnZkaP/pePuEfH/IHZOyQ
LLdj1QMdJKOPsY6G9g8GNh66GCkjOnmKNcvD9ysQLY4/BgDTyuxqzyOfgAlOvtolGIOaoZBmTfz1
mwLKXX90jmVMUvD9QsZMbXiaR7VOA4jjctVnPgQzJvgoY+1umo78Hgx6hzqB+CEcR3WbaCzrhUt3
jZtdfSaezSvka6k/7A/jn0UWaWUVtmnPTKVdVsjsbzRDlCuWjIVsnYbWnQDwqm91PAThGJ8mwX5F
GJPhFlfxhEDrA+z8gzDacm61EdIqzZ6PnTUzTaA2OiKI2Dvw4CsVsLVY9vOvMM719TrlTWqHVYY9
h+LjNqdoUn99p/4D1ws1wRtVXHCACpOn0Q13HdnbwLLqIsPG5IU9JdkG6n3QE2B1PAkTvwlPJPh9
Sz4ohNHTaMoZF1f9bBWOs6BL4cE6OQjtES3Mw/Sq6bApo6PPHUzgbcSt/NGMrzRwMePRW7+FlZpB
F/tJHy55evm8GUa4Cu+DE/9f17/UVUNI9lCkheW+p/1VGr655MNQFOXP0YI2pSNG9hJvxHEYl2p5
a5qsGGQokcN0T7KS9RMnM22k05/hukHiIJwOQjvYOqXN2ITIs3xdvBTDv+OmsE/O0btWeh4wRFpS
GWRVKsWjyHfK8X+GXep89ErpU6qqb+v0bBwAXfs/PhqndmPp4yvzVcGjYs+NInGG2DJsLM5L9hFh
uvWRip1y6RtfPjfe7aQ7tgWO4GgAHUZ9DJTJe/wC3Rlm8YcL6H9wcM/WKhnIqO7WUQIjcPU4713F
LGW/PazEIC4KsAG301BpjtWcHgS3N4Tg/HwYLVSAFhe1gN1Amm1Vij96YR4M3mdFfT5C1KSZI3kA
Etr3kQxuSkldqXIaZU5PG5VOF0deasYvLR7091T6qzszGSzQ0RgN/iYmnjJlhvcj6r9pZtCEznJ6
KFs/66CgksuV9Ktd1nI5Mnr0RX6UD+jllXX3l0Cjv5bmEb4IQRspZWtHbY4CSqvDbsTQgA3Ri/ez
JPqnMA0mHAS+XLsY2FHqSxcQp5HTNwxS0g9Q2brolUb9JTult7ACTuZBVNXGCcCCZTUVPc7F5ZJJ
X6J7PfessN8eTdwzo4A0XMVaTNXFyaHBAPX4ffEJ8vaqqp5jR2glq+qr4dV70/Jzk21ZxAUPqP7S
OIjI214c2JkBd8c5XBhxudYZhkAkWp4vIhyHVZPF1iCH7PYpYUGJBCnG7Ha6TKI65SCgXM5yT138
GX47N9NTzuTbaMhUvjbO0XRAseMUBgL07tqdukhnSBySobhqe5fJ26Tar+jRc4b3C/H2WkfcXjVm
TF7P0E8yjIR2Ryphj9PEfC8WvyJG2DVeNo83gB42Wx6VDi176T/RRGLsswgHbE/wcL4lxZWPMJJV
2J2QLfLzOAdXBDdBUvKefyzJcAfuJ7k9zpvbJngstjEKQmJqZFilIAW9+cXNMTq/ua40QXZayoBp
TIhxWGQN3x646IkyRnmDpQsmNqnstFYWHZMadiP0fTqPc5KKHoIJrOe+ll5bFaI1Q2TpxjdaxWHG
EzcG/bE7OgXKOoaeos7U2JVWxPO0C2JtwBcGqU1e+rgfd8v1p4ZLmsZ93KIjPvQrtKoJRkJz/qxb
/4Oqv7Dqq3gnmuGi+87vYNybMNa/J+MfJxIS3G5Vz3a7p/zvZqIxLIhAAwuon7FFaP6gM8HalmMZ
wyjBfYKIcdQo6r2yhhYNl3AEba1dpk66IchrzXUwPyYlFcPBb0PbAbal2SxlG/mJ6mhyYlW3rzU3
u5i+TCzcqIbbF7sn5botjbAXj4TSWpXH68YKHNAC7fIb+BtNaJkQt2CTzD1MMfiSGX6AZVkA15cH
TmkC+M23VhvS2i1+0rWijB7Sq9LkhT3Gzb0mx0ThubcxBsphU2gkXTfQX8+ZpVuTJwi26X4sT05M
BQ03Nl/fHjDvtCXvDsEF2wfHq5ER6gBRHB5GwEmUi9A3RMkVGDefhiCC2IYasdmGQSabYtjNZLg4
XeIuP54vYGz+m2w1HrNrs6OFFzaeqp/5GX9IA3M3VexVS3kVpHVHVnmE6KWgfxDv0FUxsVlsoGjE
/pJd0neMg66VGodiyHRlbu+Fea555la6YLav3CFJaQDzVSoFTOlAVem4X/NjVLZvORVff6ccYJ2h
JsQl24gt48E9QqBkFx7akSN7XSB083wvxrmE4MCoJJRY1BQVwoGDLFfxRqJCL8nTZpobdVlmEcLg
WPFuHoz2qRPYfhl4FDW+cz5YrlfMPyXb6ONCADILv158OfJ4u2nbg2bllJCMY++gOpgBe5Gpl6zZ
sakzWPv4CNNbp0mpgW/VGwbl7J8P/Kkt6KCfwvq0Le0iNljUOmTaZsnnxjAkcrm68/LhpBCMMmWM
xPRgzNuiku6DwG4GsVP/imntbG47KGBYr5e482W3OegWEkC78NERgZzBrrKRQBBuGXNmqX3/RvHM
KXrDy3tkrYVAA3pxvl9gKzOJB+KfIoQ4/Vb4gy85iLE/fnFxhsC0YN6SaecNx6l6O+fzSGtLJTU7
gLFsPa0gp25YWW01yYOKOUe4RTakPV5AcHWhw6s5XD30XjpmB44/FnkeSeBnwBOCsmhfu4OemONb
FTONLdVw28TlAg3VFL1yABJkebEzO5yp/CpnOqu4Z5GF4NRszdyN4DbOuwJ4zAbhuJ2rNAxI8Hv4
YcxNZ1qeb7Hygtgp4jmcio96yXLD4i+/W2izmKazcqi+NntFPovmiA/9Ysfy5wX/AXm5EBNe0RbJ
lHAivXPIWqOh8BhVdDsqfnBCLgeVdh34navckMSTl+hyXCZZpI/xMfnF01doRpdxT1TnXOd3gAch
jAhDR0i090LhmIrbidDWr87YpP3F78COvKbIx594IOrDaraVt+u8HF4Vs3Vqmg/Ta/bzFf/SA0R7
nfYrjVoBQQeZB8tIoLjlWp4LOyVyndJrg6d3m018yTSkZgNGBiSwF1j1r2H6Lu3/PdZjT79GQ314
ODIRpXkeLHbtD+YOdvgpUUX/QhhXVsvt262Uegevj35vzkECp5mZL83lhQkRa1Ng5NrBZAxxg6qU
OCf774B/dJNH4dgAiUg6r0LFOdJe4wBvsNUilHGJExQlJYU8g0X7mV7scsDf2qfA6O9VPTjgOq/a
XJywVxeJgqrp0JXaz8zDAjZUpcNMlnM3N46/hGjZ/BNn+a9RmMaPlVoR6uHe70sbflT6OHs362N2
AybX+EvwhJ/bfxh9R2Hw0rDRi1uM9A/0fhk78qBGEwGrBwk1j4QApBTAd1xgIMsM8ouu/2RH6iuX
M495AmybnaiWA/Ty4t86J2KcXVzcWsNZSpqMPFFZRB+9S34tTfgWNxBNyv3pWxWzLRMzc1TZKOhe
MNfbUAAM7ofvUtwMNfcW7M0/ttKEHTNm2pIOUdlc9h4OfX3hZhnwB/Z44+Qm3JYHlZWMtv0Zl3tU
coX6VdNwwQVXFLvIQPY+K6zk6VMSErg+GnRxEz48fbsMuwhD3sGUasx7Ba+ageF0uDv/67aVyC0a
bt7Op+sljRWf4eqktfM7jhPGiMAFBD+jIHczg2FEfWT19kz3ceMDKEb6qVL7UdtjhFaIfkMN/p08
IH6Xat+Vmiwczi8265Si4XiSlhxiHIJAUSlfnNDCgXvlVveWVT6xEe4ViJC2nQ0TVFUguCRMGfGs
z7OJvI+nvrn9SwrzboxMwnK4Iiwm1Ai0vaRsdiVxYitADNxNOHfJpZbuPKW1pXrMU2K4XinZ5jU5
ww2LzHwIMjJvtGOjuSsJ9XI9J9ZkD+KKdA0ZFjBT26wTl+P4A5rzrK4cUJKXVNcKG8srNH/lt7+w
cMtNwhX1E1GHvzO0l5ELMfBBapofzyJFvvdMamqKsBRUOLTGBHVSbI2VPejEt8gNIveJSj2ExMNI
9SJ0OnAdNLoNxpE+yMLtbnlldFxC/f9CqjhvpuAB2otIuChLqGDXj+mzKdZ2wcXLF9HAikQOUp2G
ndGBxHIuFaCSuhCt3oBK2RJa7M7V40QraZvuNv85PZplCu5wgV+wQpzSP7ZIqqta37IyO2s31F2s
GBloRS6BJ+XPBhVQoMz9M39k441wEQsEnN4NxxBoNox9r13HLtau2YviZd/GQufWhEstQOkDyyc1
jbk7QA9gcFzDfOEQF6mb2VwCVnUfnVHQG00Gz4dN5oyz4fqnxZrE2BCYX+u/fD5FqX+YKq49x/5c
iQeK/n9fPe2L0LltQnydnrqHtI79MR8T4HDfpSlcNsHlMDOGG2L/qJyjIuvRtJvUFnIpen/Mx6ua
VvuQ2F7IeCdoZG6j5k4mX4lT7VCNJwXJSRJ/eZBHFjaiXe8m7cDjgQ5R+NBY+c9aqPMlE9GU2CVr
GwO+meEHoNZWfjDYpSGOQtU1DAP8/Wnc7fPhw2e7PtSuLELE0Xnd3zHuaWojLdDwlWrv+ljrzLyb
iYXvBWZcsThTeGhMmZKQ0Whca/w6Oe9usNfYwuLDasb9Xy+Tln8m87RCDwBrCUaihwBVVh3wHjqy
fd5PJm804Jxgpvg9zg0JEx7u8+F8xCht2H6r5GmuxZOh9LBpUgCncze6zZdKRfsKXts2xta/0o7P
2wgc9t3CNQrjZA2EuNfdDxSrVYjtaAJcMICfbzO09O50s/DJJK3ei8NtegUDvHK7+ISZJBPKPZ0J
NY/CafLZLAjv70QA2JYUqzsXRsiUr3CIl2Ti91UIKN2ezEUBkn4UoRmd0OorURIodhJvahWva7Cd
YhnEjOecs7pxPgE5TXrs9Y4jvKhSkCDc+8OC1rsZwN6oNR6vQ0Q1ljRifKY/jekoBn/5Ld6Q7W4Q
u5HktXrXHfw1h2pbbA+M/maw00R0VFjWJwof0R5stCVU5qmA4/vct8uu3/jNokWRUpLKSXauHTO2
xejh4SzRiqIEHdsnhDV2OIzSrzoK2W9DDFZsGEQ8ia5j4Ci9DT2WFkz+/l0pWE7IIHKBqZSiHs4G
fGXCDzNJcA9CYGv2r0BPUpMLP0LiBoZ7FmqX8c3LLRCqPZ0cA1HupSBtO0S/K0dxNaJbnpDIRlc3
Vq2i6+69N4LPLvqPG6dOBfm9D/sYL+8kQ8fHHwClvaqGtIb/ZIl8Xi/zCsDAKrmuyEa6ZrrRxi4D
o2X13c/qBQOByQXxxNfDEJqYK6cbSAxJUzJOZ/7GnoaXr9r8FQPlAaGtsYyguuGktkzWDHNK2YuM
556ATLVkBzr+C/qlgrrDgWtAqR/0lzSs+26ECP5NzzhxnS1SxjUf6MkzgVXsKJdw+/HJalRXJ9z0
51bP4oYoPS+fMjTmebpBSwIrnGDHXTxJZZwWMh7/EY/sGUpZHlyQmBIKY+Q03kHjZMVDv1LAztIi
Iv3g4IvrS03mtceskOrZmnrjz9S4tlHz4aKI+Geu5nKbkEVWjoswh+LE9DDOGOE1BCnGQfHkdKmF
mCLk6WqxYOwNwWEew1wtYKh7UpCEwpF3r5r+BLjUvGrzEaYW36XnPlzJHSIOU+m1BNMde6/4KQbS
3LNZMFGBd2/eavl33HkQXlNI5sSeKq9M/qsmmJ+CP1ZBXOeYmfStLEd5RltF1ak1s7qnCsnqEijI
X1uEmhvzjIx2h2iEEcMjmHD+9tpHA/4qfhPpOCHH2JU1iVpS7Rp4ko+JzWlmo68f1IUmPUVkZbgV
6UN79OEJ5SKcV3DRZzshftxVS33dr08BI5f9eB9f2YunCWq+rjBISZq6ozuCAzIN0Wiyn4w9yaob
+VneiqZRHW+ydN9i/5ekS0y1exD/L9qTWDGO0smRC2ONQvk2fcVFL8w0prlajk6ShTLoGbmAPmIX
wonHKomofiiBzl9vDbbk39BpleIrxXZjcruNQttLs9gPRElauWLn9GxJqn8LR4mlKSswEI4776Wf
h7MelL3YiAaBUMrSoagQwp3neyL1T0ZarPUN0IGPZtURaQSqDnVtJaPsNUMP31IUDa2rixrbtiKX
K5/GVflW6JgFflkCVJqyj5ff4AHYGsiV0CkIbxYFqGDRWyI4g/voL36xoYVBWiMkpyTxRp0FsIhe
0HOmyk3SyZnobPQtLHIWyQW3MMQBYLVz1uwiXBVvihb8N4tHNI1dCSxOPwHj9ShvHMzL9JtISCJw
rnKZDO1Ki9v0c5Uam+zRmbuLj+pF8KYRRn+/6C/f+5YqhjT0okqkjhz7Hd8pkCEpfziz/gQa3Xi6
6VSx/U9y6wCj6G0m0MY0vkP/no+jjq7a5OcucpaJDXC2a3hgT+WB2R4wU1fNnxN7oaTWUSEDArZS
jyL6k3KZLPLFDtsrFRT1PBVonY6wF7pM9zkuq5xLBng3QihtKH19Y/0UXI9mYcM8WqcN7NKzXnS7
ERe4fb8aRNcsaKR1Np71IkJcgonOs+vdhP8RwuKK5u8in8yrOcycNe0nHZojf4MLbNquFRXgIoPT
DkjCgKN+4vNdcHki3sI0zBPfiKxG+6dvaPxofVNsyYRXbm5K42s78rfUkkZcRM55/EdIGPQMUiFI
WEQlog2FU0CXfVMmr/8sE9IrxnWKN0QdTgJ2+yQx9Er0/V4LieMk/8LWMVAcKJ8Y0GLXmqlIjE/U
kCDpF4vcrqAG5fAZxDF41Auz0PVk0AM/4LIwQE6vGMQoeT0A9gr/eKSp5mLxzshpTxTkcJ2e7k8T
wxhMKIkr5UBdvymSJEVOip5/ZSnxQngoepR4wgMLNJQY6b5B3vSxhR8oFo5ONNQQf/JWyklUmNIJ
SUrQiueT0U6Vq4b/aE3d9ymplNgbIE/02rJq5HkOC2EUX0Paf1We+hOxhp3tQUFph2OGELMZUoQm
Mj5cXPQMBKcKUslgJEzF/uqY2LOToNcDhPrY37DbXAjGPpO1ndfWs3nyov+wacyvvmbeHGIYPp57
UF2qHnIFmiQQHwCNMH4gcQ1S5OMcVt6mlGDxKKAI9OtwAvRJ42C+yJ9L+tp8Hh4ykn07l7viD5HL
/I0Tjuqm+llYSVf0atz+lr6ftd5b0IUsZjViCrEEy8aPBX6/h+3XBFWTAOhCUhJ5lu48xskyxP9/
idJ+nDp9HZ6sF6NIvINp/sQy+j8qWjEieVwScIjFQkbLzAttfAAbzz7o08DTNst/XqJ5bkCvGBOF
n3XONH/ld0XxKjh2RjP75xzzHt96IGR0qV64w7w5SEicBPGH8Np7ABeC+Wqxaec/TZLkvJKQws2S
/mpn5RMB7kqANK+ohCottu9efovFSuWubssukInRv3670yNHTFkzJg/5gvinkiSQAYIDNzObeJyh
TQ2DTbn221zlTungDM4XTZX5Ujqj88g/B3QKiTkB9n9RAJ0VapUBTkALz26D1cEDHqnpjsPG8LIT
XPZx/p049tZnBBsOjHZMcv7L4pttxr+HbWtTOyscyzsmKNRDX5A053m64xL4c3UPTHJ9ac23xKoF
LRhunCUlcvBKocrEut3kl/1XBUfmPe+eoreSPzhtD3w37D4iKKccSoYEF7WFkGn9qet6lHFvnyqt
zJOIRSSW8HLdSpNvOb3/AEn5wLWSA/+nIKPPd8XjZpqMu3l314mm1DsCsM3utXH9ZTTDW6d4WtqJ
sAlVk6rmNZ4r2GR7mkx85MAmYb7C3xgOzepR1aW6/jKsmCQjwDJTsnsfIHu+hurMYCekKLXht2AA
4fPre50oM7vqZRngx3pUcPvs1WVREYLqK6e93QnIXwcU74Cuev+x/uFzeWbDu5FZWofYh8hb8uvx
4HyuA6TMfsA1RnOxUe4H3+XUz1OnMhh5dci30VarRtjWuuFOCPTwJMq0AS43279s1btNFuhizBaO
AAJVy0jUaq0vLQ8lHS7pZMyInoGenIcnOom2D6Nj69x6MRuyudnomtPwqthMBT1yQ4x45ggtO6a8
6Ur1CceB5QVAz+bTjRBGQiNLUjndjiY5aybz8XfZRlxWW7Q+veHIOHq5OxM/Q6xNx/bB6WiAAUqQ
8LdC2/utRfiuhB4cAtnccY9eAtXSvmD6uuIe1vG8/1D8KGc6WdKR8NNV1A0fVvClx3/oB5vuTfKE
YFmU4x3UJiVeg5FP3dRI+DZzQEw+PlDA4zP4ZIpIvo0yvaQRuAZm244tmaHPKPw+OQN4T2zdVjPI
KNPD/wmTu62D1axIis4/ZqaPTY9OZ7zXzpy1KWX17+dkWe/0CGErurc05uysN/wqvChvPaPBUOTb
sNX7H3IRuGuIwYf6+BHoALpuyngYAlJvjCH20EAmklh2gtChaKvQjF8kSJhPHW2PuUq/Vpamc9Kg
4d9SPQjXl2xkD7oOFvijBEoT6m5fv3n5RscbVUtNuUOtFke7XTCpLIffWTyYxl2OgVW0tBX7Dfxs
6RcZpbZVnPRjgLFU3StInPkxt/jLDamFV+8uicGW+Lx0U2n/q+zLtONlRj20CI9t51h5gFSqaDbC
w1fo7ASGDKe+k6SvWGHtBWm9Iy+6w++jJquY3XZU2AsuBcNmoaPwaU0YvSzYaZKPCrpE0yYeiwsL
LWI+eRHdQSE+MsKH3buu7kGmYewYW35oLhdAjnj6jqdYZRY/b1WdsIVo1jTiz5TglccdjyGaM2dA
+ddV6X2rwLvrvvoCnilGDy2dWPFcmTRFe1Ee5TSO18LvF+g8dCE40c7huv7ce1ufPVDPhkXPcZkl
yMImnW375jEn+itW3qo7ITnVtyTy9KraGWI76QKkrk3X2ZqfKlBlzZ1AQYXCxzpKaY9nRTfhdy3X
GwnjfBRBSLQSyKDrrnibdECHG6hNXzO8IUCiDv+hLkcVkdymwpFu+D2AQZ13hgjvEu8yuzKzNDjj
EF000LtwMnsZTbbjjNFYw9RbsQAyWLOOieL83mmH8AOjc8k2rNx2IwPLXB4Bbn11QW/1UYOaSqkJ
Xtxo7mPeU8+JCn6922OKDIfvDQ7jjzD6W9y/zLq/ze6+bYSbK+baFXpxnzWpTdmNl6AeCE8BIQKn
Gn/6NKUICjD1U3utDY4awZvf/r9L40TkcuPA/cusRmSpQsrKrLR+zVBK038UxHZCYx1qkukTKumD
ewFkzWkLLFRcfwlN1QLsfF5naV0R0MQ2Dsq4Yn6VMgpLRGe9ox1EIzJbRoWlI/Qz58w1pJmCJpC1
jg+1AZgFq9h3ad9YU0nW60F1c4ebFNp3L8wr4FQDYZMhM4rLoAvwwSbs4RD2H+rAN3lZ81vC3wRw
njX/MqMrZgrpdyynCfERJkMqIO6hpeUvnjuqWk5KU5dKrXHjoDczTTmVttDD9OOaI0/2yO0Fb6dO
sejzeJJqs3/WrnR2/Y6E4+ZKYkOilntrPZ8Fyq4k1N+zLZ80Gu1wGV5PYlLExJd7bkzcfWNmUtZn
5XZOlZi9wPthLI9KakGAurqb9U9cTh85WEnuub9wtmssJT723RbiDh+M4n1bFoQwz+c/Cck+9J8J
iquFHEHXV3cEMwqowfAG9rRC4l9uTjb3GpsqS3s+TYXRFKQJ5yKYwuqZHrfMvmnirGBXR5Buo4Bl
FVVKAGZOYV7GgI6GfYQOlladdW5fIQzMkAWBKBloXZ9+0MKct9SvIMpR1mSCHLr26LZ+bI7V5xeh
jqiSF/kSOE2Wh1BmKYrjm3TVx0eFK4QD5RBFiQjTw+iyQkOE+d1le8fqfhp+aJDxUt8fDq6D+WAq
TbLZuGScakCndidV52I2gLntugJV1oQTd9wNIa+RAGCXNwGqRxX2mX5ClQIxuXOkry0rPM2iyq/N
pgFAP3fuvSYBDqn7zSCISbbDtGeofxCqPjUvkv0DyFoyYGnFf3KVxygp6RvBfWc2+GJ/35F/ge7k
8hiYz/QvFtBozybYzqDTOYWeHKT2IvVxb1pLHSNv8u6bdiVuTOm4zXYDBAVDOdXb5OkWk1XbvvLM
CiKK+XXHyjyQ0MCwcx4NaEc62TVrUrWYkr4lcScHLZPQ4ysDulJQU3s3NSQF/xcWewcpwOEn2FFO
lhx16C+lIEI1Z+7C6OyXJpanxgrFTTn7+VRlSQ1b15JZ9sOxyTNnGkPkuuabJfP5u7cRK7FLPVIE
SA9XnxY2hVaZsu7LZKI7CizQlf1b3RrBO16umXuCLmiXFqRK0fFDFqtnAqjYzOwcrG+zco1cBzHd
0/MPzdfn7eKX0WiTRyF9ACtx1NwW0Zki2Y0av65EpZcgdzUAXX/ejZH+EeSnAAzvElQi1wChO23r
huxSI73sBGUuL4RY03wYAZiN1xdBqNJYB1LMey3XrQpqSS8rqlLnbNI626WUPfniltFFmaUdd4YR
MIT10X2eQuUS8z5X/QCJ6D6pST0qnMtYebeiVTb5c+gaGeH8hC5mEqK4UxnXZobbpw4fyVZ3u+Bc
oNKUDekFLpiPoTxdPH5kSw2gJvKQaZksHAsaqYY8GdDxvqRiNy1z3NljL9G8aBxwUTMydhQn3msp
neDKQjKx8ygsXWP0/aaw3tolV3A1eVbss2I9mkhh6ydAHtt9Od8/1QiwQsY4glmnE83cxayNeHQj
V8zTSyzNVBh8nW/FklZpxwDeIQSOwBdnhL2CZyZzgSygzsty443kvO12sw5KJWbFSJoNs0GmdjGW
cpQu6Te8eLG1QB6nsjlEs42UHgSNjDhTedf2aNRb5ZYXv/K4c3wg0GMsKXA1J7CcYQicXFjT7h1S
gGl+gP4BoDhN/sWMBDSJYwQ0v407268LjOvuEurnBh7hwPsL/KiiFegMtPQAcMw4R2C+RrgPcTOu
y73ZpdPs1q3ahU342/bzYio9gjMhJNXWB6TjDuPUfG1+IPFMfjWAmDxhUcvYwsBHttQVUWqe7peb
fYJzDTLw6dPVw4UPoRn06a65bOMLccKgxJ0wKTy5UYOYEZUl9znpnqgLfswsa7tLZV609hbpfmvW
LFsdDE3sRBIAPpX0vkMwubRp8yDkn+RiTcF96uc/AZ8RQWqqxhp8zYBsY9d4dxhpI7fTb+gG8kci
vvy+fCnRyFlTUyS63QpKB0BHBeQGCjmE7r8BQlxJC1CzIGzRO+BgzvLWtjllXASx9vl40ljDe6fm
3upmdnV3Eyyy+0rydKbq0B773w3Cwpt5wzz3yhgqH5crcCa9EOTBM+62q7REty8Qqw1tfWE/+RlR
CX5X+VqvmW03tnCMSUhUtj9Ly03QPJhaDuNC84a3jlAO1zxApn1b8jdLm2dXb225/PjUOrg8c0mh
cYZ+fTOR/Y5GWKBF6ZijYRBMrkeCJoHYAx9+p39b7+Hi8OAD/xsFMCs5VI/Ae7MBy5SGrgPUubgp
3EaCERAMH3MoYuMfp+ZRNQx2L26rgIWDxjZo2q7AdQRdUFN/RnDwZQyYg1m4bv3nS35SHqwFLyu6
Pwo7rCrdAM+4q2nkI0H0KXBnMSZYwqL/EssYY6+Oq1aWwaXz+FuuUeFjLdkyvZuolPYREJjGJDaY
ioOz2SFcWUGZMQhkJj/Y6IvDhpyh9poFVxMfSrduyp6AjSMRK1zm9muWbEz5rFXnGGpy0AGCdre2
KNgTv091CyfDaKt35F/E2Y4kbsj5eJWw2tMlt538J2sPSsI5qmkFKnCHu4jIIHs+PdDFg/B76paL
322G4eB1prfDT17BGyYgF/mLDCQh8wehoVKP26fb5zlrgDWU+Qs6HruYy41qN001vwmCLRQu4goU
jb8l9WafTvdcaQDzfRd+h47I3QuNsEj8iLGmgxxPITgu+coQYB9kapeyqg8jsLaHAosgPWnqOaJ3
rANjebGs6FUurZn7YhCBNJeE8VYY/1hxTidmc9B2qihdKcLaTFXr/0hr9jdJoa1TXKXIC6E6m8De
L6DSYlDTdnSonhC039pDJ1k7JHvvyAd8YBEklUTQGVbuFTUMPGy++ljc+XLtkxMlmTLQpZRXgdYw
ZVTCfS8e62NVmN/BA4QyXQ3FzEo9VWp9FHPCFbYm0BEMWl9/Tt+vwd75jmT/OxicWCrp4tLoXabp
1eD8DU8HijL0Xu+eSqcZWSq0ihBJW+Ys9DH69GwDADK7bG/SoOaRn9DkLsFt9uLFCalo14N3EOtc
hqouP7G3ZsrhuWwYM2aECmiCqsLai4TPe2UCGxbdbHNYUNMFYUqDHdVr3gRwDZiQ325EEWydE9f+
1VV8INwdTymhnOWnRbLbCS9y1tHh7MmJUhedqgx5phHaTAw2uf+Er8v34c0s3n/mqxMcVwjJ0X5O
4B3xizNqfSwSjm4oD//L5tspRqLSK3yJi/55eh8/jh6TrSFWqYxNINAKtSSgvhpMdt4wlJNis/s1
2yDJ15GyRE4oOlOR+QG7CVcVMp08red+UajkmNNXE7OyP6XHPrGJVtQvu5JjwqO/t+2yImdVBx16
1WEO70BlfFTMtAKlMc9M0FNfiL5YnYaHPuIQ7SdUyqGTi07NDDdc9nRlBxIbUwN2ws2/FBn8vOUR
MVe9W/Xh5UkKoqkyHXfRpU0ccl2ajjc9lSEB5GwZnXZ/sCrAV7H/21jB++MvGls4uN9mkzqdqAsz
OnZDSXUVhOn5whsGrBd7HG0qW5BcF3lUNGQWyciGodWxBNuuzsnP8ejnsywx4XyBAZSXetYcR6Rq
TjVaOdaMfx3ssoZaPbjgXhXrhOvuVoszNquCuJ89+Le5keP5XTnzfUw5GcdUYZ7e7lRXGuixcvTm
pghhUha2ZXKDx6YiZbaq+QfibzQ81/MDoxbmS8D5X866/iQSwD+zdaeBWj6X1RF0/Vrxke6/GR13
5emHbxVfz0ffiYdQ1TvmS3b+RXKIQLHzPGmTCHRIoEy3pu+kNbfJPTuy1x8sLIMP/HGhcsH7x++e
16pez7At96egNapQkY4hj3ciH24Ei42UHQ2MLH//RGxY+BA6hRvDY1grwyoE3KwFmnLy82AXYLvT
z3okWh1ySmiTlV4ObEyeRFAu6I2HCuPNVKqRbzNUZJqgtgdZJRUOG88Qj85fG5Gm22kybXoxz0ct
bnvfKBdCymYsDQA6mWhWoxhspqvlLM/u+XnEZJo6BmdLhGXT14OO2bxVV8MHRPAIbuhCLxMj3F9A
LZ7c3I1UqRsrCLyCTDqV7pwuwMvwsJ4hn2Wln/hOKf5pDeNGAyGMKjjtaI1lByRNWqphg17elrBQ
qDU6SJ7QAmmVbVPjsBueOWBrZ7AHb7VcPXnDIwzWP0mQ6/ru7xUPijJP0yrb7quCHS5Ux1GaetsP
v6tJvnRUMFkxiBP19hU8UUlYCGwJEzF7YmThy7w8f2Gjy96PsMZ+v0daXF16NGQRdZM4niwlabi5
tXOHo5z/7GhiXqgUlDGwDHEMv5N9oxsC7MKXkZKKoM0U7orEWjOMwH6RGajdIRvv5WmzUvStz6K7
cf5e790mupJrEj9c5UD2EjxZpmZ40n3L+RbPsQGLkmK0lsrD1kkMGuxcviZ8gHcI49iR3tlKHNP8
uLsBYQ4NxTPc4dTBRXZs9TvOYXhCJOr49YiYEOgU/gRJ75kCsWivjxSZfCwTEyVF9ofupw8yP7FN
yhTYKvgsxBWg79ZhtrffLvfykFkN/Gp2lBHPmngplUf1qspLxNQOQnDkoQaVK1c4owFN7Awwlrnx
eWefM3/OL7xCsaRbqaKk/ZqYXH0EZDLOxTp8YaLMTmOpapPNYjkvcDU/klKTsePFUwa/D+VLPNc9
UajOiKjy4/xu5RdztnHFqly6u2L//9zMFkRmyOYde6HtomWA+0xnQn/mEeqyIoBoz/AC2Fvk9fHS
wSoMYTa9NWSw5ohfkivK4/CLdjp7bMFuCD5+t7L85V3im/ATgvuhj2ilLbO3rkwyjpBLo/PR4b9F
iXLLhUSpktRpzrWTFh+4NAImE304ASJnMTBbBOgTwQbarUhsrqCr0DYqonbA/lc+PpX6A2EJUzuB
UNvaqYsQx0R3SxwB0Cbt5C0kKDbPuHUCYQPWm8uZH6FiVypnnOmwEif9UcFQkM3fw9ZngzoLnlou
+HfqJvBIATD6l6ElLeGjgF+L34lPPxGaVbIHiW0PXgBDzR0myCiLSUMu55Ev+q1n3JSmfE/gxSdx
PUf2MU2n86pwetDcy4WsUzt3l3ScanbeV8eaqm0Cmre6T5AZifoWHttQGaKI3J1Le8j6YCQyHfXb
kK38+y40Rn7ttGjNlp3KLU3rtASLowBuo2RIKE1Pdjqgs9X0LzBzP+gzJyOBv3tadm3rTmkSrRD1
ksIiJofTzvLJ6B8PzXR70GJVYH4PQcOoooLLAj5lqz5s7kyXLfwsjKGejS0eJVZ7jR7Z6EQtIleV
wxmAEIl50/3h+/Uw21/d9TmaMYFGPScLM6dSr2z0J+a9QesNnUUNrtLN72D4T+7vQNcIPQfJHyoa
a/bWbkoKPoIM11nEP+OVrfOQ1SO1iv5QI48o88trPJKs2jiL++UAh4vBUXnWYlNmBeztGSdQ/cOM
qTCsr1g359WU9I7BTvjggq4Dr1cPKqndlluwQX0XUKf7/dooCj7xpG9x/3wcV8GSA+QEOTWW7x5V
oJWuvHILHXPrstZCIWATQMT9kdhi/QfdjInxkYsfH6zvZmLMf4jpn6eOEUHd6ToFFoWA/bKCc31x
BG47SLR78PIO6WvCE2z+LM5IXVhgYr4ojlzTqNgxbnDOBwpkyVMKiutU7Dbk19xvIWsXPHeCGuZi
wfdi28Ts4fI4NFb/jCIX5PdT1cy2XU314OABnCGa1rkO6YimN3sjZoLLRQKmGk3KTy4g8ZUdxX/y
7doMsHPA97/93SIjClyvDWsqaY6ibrA3wQWTeXTLxq+ydsVKMuYRJBXLeXZC3fRdg5roaivthA1/
40nBbhkeeo6Vbq3SB55SyUu8x2Aq3P6Wz3LAOcwiow9u9YwlmgfjZRunum2uJEghw86nwllFxhBF
F/1Zy8s6N/sTujZYJMPh34NBQUn7Wdj1FU2xZFLYv28kmgWD3k8d6QtLAb/GHT/1NTYqYxVj0c1h
8d3K4CGTUDYuyrFBzS68Ke4UYv+tl+o9ySbcgKJeiOlJUoCvlZNjybcow/WbaJ1Rx1+AqzX/XvGL
bFsILt2uyj0FBfr3bV+snh4oXONpoZmNwYH4kmm/xvWpGPhoz2kjIkLo/UrfCYP3BRKJZokhUG3E
2RkLu9vifKcpCk172ZhPSjVlPmdKP4dVjMoFKrjFUCNNDjbTkpLJMJPy4AZCyi/mtRo+eSrEiKMg
OvprSDrCmJqOVTaxiGnes+AYOv6PRK1kQV+0PTGPPuFQ0t0hKVYqjqH1CQMNJZchGoBnkp4p35NR
C4ssnAlmnFyihCyT+ZrXjHy2yvyRC9k82Ur0Yik2ikj9jqEvrRLmOxbKBnuSL7oOCbNB9KoclKVw
/DfNIV5P8aAytE1Nu82AyDuxQ6wOMn7WaRxbORqH1FjNA5nGQC3brscMUVnde0TPqy2VgadRQ20A
hbTtrMuoSfQjeUTavcjdlficKYn85Syul69dOFoitfDkwIeiaJJC9hBRNldCr3dEnXyDHF5lTF2y
RPqSACIalqoo/Irrlz2BI8ald/QwrOh1RYZQnJar8G7m5+J4Q+zupRZ6oDKxsBkgK/mIxUMMvJGi
MWWE8h6+pmY2liCQ3VL93qfnY2IzyhFKtkhOl7Yn7Eg3Ay6McxGlPt3vk/DaQ10EGU1j8T74yafc
ekKMiS3Qa2M4j46o4t3esEH2Il5HhK/4yzYByDow93vRaiudTFoE0NQM2TToE5tdtt0P+bGQHRBQ
wthwY2lJSALFbhT0bXc/eqOB9+yvdCVqkD95wrWeZM25hFaT1qyAPmOHg5YgOCzzqcxqV4ZkvHeP
51cpalGPQOHrHB1BWnWWr7Mz3sQr8XnqPEbZ9bJoPzGMowpcoRo3YGy0kSTl89SwZDm6EcsqztUe
EOwSELJiJJbRsH0Kd544NPXob87L/Qge/OgzOhUTXRsrpIN/D1Zn9n7vKiEMxCOlHI9jRlLigTX0
IziiV5ZkpikWYyfAlj9++f3RcxkasXczb4ZJElHbHL4INWJJmeScgZm88eErTeSM0WkJL4OJomXv
VaH4l8xLXjyxuoIWZ4ll+8e/G0PlSrDZiTm1Qdc9A6Z1r0T7NErZhmeGDvbXl1VdBv0cV4tGxHOJ
8oFinZSAaUakrkZk5mWKUQoSMJjMXxtV/GiPjwm3P/Jf1L0bjjb8KmLIDBsXDmbqG0rnrfnpCxxy
Vg6mOZDxpgpPdsB6gTkL6IDXgGUiseIDF2kNLsiagK4XLDjodd/i70Sh59IWBOwopOFgtGaPURMy
4/6VW548uYbBEVfYTpS+j3AGRKwBH27IU+DTvoK4ElkuctbALKuRl3kcWqIhD2cETIaBKl+w+my2
Dmf1PIpVFjNwatqLqegx8GmV6d8KO/ZPNZ6/Ug3fQsNZqlxxZFUckGGmNQi2F5hC2I5r44ptLXzz
4MzlKsdzjJCccWQtMiYFg9z7pfqevpcImv3k1Q+F2bQM9XXjJt4m1FxAJ01xFrPz7mm0+Il6WGxN
bLVfJQnyuYSIY9e2JruCkbxrfwFxrWKIYRmF1elxe1eROblHppDKZqb2dRitwyaNeH213WThpsjb
kHtz9501Wkfn0Bbou8nSRwNCCiQozFR0QwcL88lu+O73ZZtvh643VMiULSeHdRRO9oO4JMjz5ohN
FGxPEMso6/RTHy3EmecYqILb8iHTQ/X4oJ9IBbdRROJOS/CnXpMQxxArD9ZHZ3nL5atircLh/DpG
QSE2UMqUk9Bc/4RNYJp/DVj9AWDqmYm22XWifnSc0qqZK41q244hg2WTVrzYz9QjhD7r1qnIrG4K
EbgKQB78StTKjq/DNpUfo/2G90AAd0/Yjj/RyLCeDpx2E17pPGW6WOS4d8p9bbgf6JybbCOfL+fX
ch43juUB8heauw29RHi1cbRrENsc6FonxS6gFIHcoDBvsHNa87Jooi31GO8Qynt/Z3l+hQN5b6Va
JjosB5KzYeU17pJ30k1BgLGj/e42Z6HbrwX3kucrZ01WkrnL3vHVUQxFArDUN6S6Vz9NeCwjtdsh
UUZa3NV2u0XwTAB4C6Dm80G7Xc9gPm10up22xPV8AJNJz+0+sJOD5On7hBrornZArfErB2G998Qu
s8c/Vm96Ci4BK5RE3mumfL5g1zuMaHxbZyXEt466ChZHUA8UTKBe5VEnXaE29P/hFk3GxyIgOrK6
1asi+h/5FbC4oTWWg/luyEUakBGHJetac2BhDVYvZxLKc/6MvNsdoYJv/BzxLgOtslzKv92QB0ZX
ePX+huKod9NcnJ+mDAVwgObM0sijBD7IYZ1/ahPm5S6KZxAPROZW+cUnBg7I2RWFSa7qenMmOtem
n8C6nHe6gTIav3Jz4WntH1OkRys9qdYD0eGei8v800qIvHtlcZSQ0IL8EeDvQEndV5K3g67gG1Od
h2qWnltJgqmukKvr0T0/Vdk3AB+Y52zLfjdqrl4aNVY1P0EXj2APRdsgBgpez7SfZirzT4BQDciR
F09tHL59ZtkylhwYS+nWW2+DprsqaEeWMOGGttdyxbdiFAt4E87BkS2hE0DIMrBDwjyOPRKSs3qO
9lIHUT/tRURcorKx5hlE3rJHoSEc+FD5NZUWGMKkOzIE8prh5BaD9RT4f5oiyGt3dWw0huMuiEwp
YDcL9EspAH0zwRuKFiMmSv8JR0brqSmsZKCFgM9yNlSL9j2L+Pkb/QWSW9Zb/cT48VviS8p1TcaT
pf7rNNuLJrzZryvYRIkBsNfImu44dXd14IpHeTzsoM+/XlH6hdfbaPJlZ9uTFjMHrq2x9UqJjcje
DW7vGg1H589aGFSADz3Gq8+PusdfvUpKA5cr/ABNEZ96LA3sUXG9gzWxcm9hXRkR8SDxhX31YS85
WxW5cxK7XAmUdFs87VhavdKz2k89dJuspoWOOyu7YaaTba3vzKmR0idr2+mbVvhPtUZYLSKwICf1
RgnVJA4GbINQBsakPRRG0Yve6Iyif9N+8DOlaDAQTvK7Bp0IoP74WdDXBEDJmHDRMFVqytOW7/b2
YALLhRc8a6/QeOqlJyB8PrFs4kp5wv+cWiVf6Kv8a9u/4+1e85DXwkYDg6biG79WXP11WWcXIUW6
A/xS9PBEsxUPbIrFbTnxYCaytARy30Cl4WdsPDHbkC2MhSem6ruCTZ9UNBVjH2DsuChAHdDroemW
XyaGHV2hj4JbtDRU8BPkiQwqsrlWMrV0xMUixu4fx5ZuJUZpEMS9gMcDJLT6MUeq0DmqdpU00r5x
8pZGX4dlDPP2OMGWzPdTNNNk6jXgUlDrNQ0+/m2uIH+0LJ4mqjfBkbOc+Yv63H9Pqp3r37AS+Ggj
V496/1Tv11cIFo16yQ2x1aiMryZiOLGp74J2dFUILVtGdeMK2sWN51x59RDl6ly2XVxQMM/JHATT
5rCXMnLgcFZsHoqLbDO9ZXrUFV9Q8V8D+me8fngAuwBw5oR1lGquKuPR3OcLbomu73tuMzofPvng
qxaRYPsa+gZvAimIityQBtB/uB2HUmLguIzsVoYKcBWNh0KY+eE0oIvafVNjPPDR171X7uVr4FVx
qSdTz0GziSb5RrFP6hV5GHADgnUMjFGbQuAK9vJDeaLyuqu+DamKGMJO+DVt7AaPOcK0ncnBwroq
LW/oTDbRbLzGUxHypzpNEZu3q5gqvB3Cd/sUg8rxTHcbHSai6sg1Ufs27NFDDc20/k0h0HOICve/
LmYuOPrqqTCu+i9xyWgiUXMAnpnm3BhT0Pc83D/iP6RCaZZL1G3lmikfjnnFp7XVrln2jL1fh8x/
uL1Z/T3UCT96UJ0Hq8A3118zaJewnDKZzrNSh54MR9YkH9HYhn8nBELv0ZN0Mcj76JCgjyqJsdXD
1K63ltHwI8EahQ7CL464x0rbAvsRYMNdJ0838wZ7L8GygNZdUjg+beVk5KP3IiMBHu60ExFzLjzt
pIDtSfTD6iPCwtfoyAy6EuYLrPV9P+0dnhlMi8GhOkKLaAwBYvdD/XiO9RNmB9Uu46q1J1EGYVNr
qd+ssDzW7XCvUFhz0VumeH07FOcTBeLfUkkkA0T1MzZDrR8TgrfKT8uM+MFwQ7kzNnyT/mleyL/Q
fCbejH13hkpeJ12pvbTkyuE19Ug3DCCnfiMk+GPSsVlNapRS5E/6VinE0qQUtOTw8byayIxayzjr
1n++ZmdVPBrvTpi/B0D82DVhgw5ty/isDEa48QIKNMnFK4USRxx/utruBqjiSMFIosFSjU6jGzt7
kNMrEBKC6kBxUPoFnVHUuBWCVhj33hhspgKDwoDp8HjCPFLoza17+xNx1fX9bzoOkoIdn7fp+JSF
Z8vMC00kltjMYgyariBmiCdBnq4RjEDnCKS1LRE9dTWUb2sAuLmJG4W7Blb+1hF6lSVK6le2kPKs
HnKs1LiAbdbk+a2BfDPPTChVFIUelUzWEI3cOsBhQyWZ4OOPZ2v0Z/LqmA2Ri+T9VGvxDSwHrbO3
RjwGj2CmUNnyalgQjbNrnZaYk5mpWKxqENM72OObAiApIYodUP8JbVORUPafowLgT2TGllF0gWX6
Tkso3rbPiUxxfaMX6tQwNNnxUmS7SxhwY8rUtR65P5vpHaJHuRGK5MahwcRvJOohLKRYL8XvVQJ5
NY2vQxDrDeHzT6dm4svjRAGmSluOfgLP8BmcFisO1Due4Fy+lzA/dM/Ey1G/WhcDZeMO77lE+2vW
4QgbxAK7fp4vKS9JrKM6ZhYTd0E/mm49tP/1AkyaN279eEeqdkitDDKagqE9+JH7Phahpr8hCZ67
boPWHqjKiWc+2kQMhT5vg+MMzC5dTgOh+t0IUX4VkBYnGOnrqDP+qybF84CUuXPAHByP3T3ZPqqw
xYwHV7tvmdtMSZJuJgl3ZCGRCYApllEZwFUgfftibZG501hCxqg1LHnxg5QtdYYz2QMHLMwl2Pnu
WGdNVmEyOAanUwZfVTcg4OyV5DVKBnytwqSvNyTkK9JmI/EYTlCO2+gIEKP/f0WXfhEOmhz/KitS
IeEugrSaR1jiiz3Mv1LdE58/qOxWwarawKa+kJZhDyPX8mdmMojv4GnJcj3M2zqcGYr7rWrXQs/I
7lEl8rOby7eK2/beHPOas9qNHqcGeh3xHPZX61Xg/mnzfP8IA345Fg2ED9xfIbvokz40F5QJSCG7
MQkz6yubW02IHOVI77sW1g/VTEI3GluQ1RYErUYR2IyImC+aFiK6kLFAPGc0m4rRItYren30uvcu
Z7537w31ppCQkh+jMYIYWIbFLn4/tZSxgC6RA4s2rVztsin2ZcdrpPCI+0Pyg1XzfWlkzm093hca
Fqw7PuG60OXuKSQ9Na8eBwHCxnPdEz02bVhldmAX+egMqKBi9B244ignLn0Pv9ep+qvxbK1k3FLZ
OSD+IfTYRbvmrktT3mi+7hswRGW/HB5/vaiJuUCdYyF5u7Yz8bleubWYQRBd0IgUkeINfkNW3Yfn
MVWWtyyAGv7940KQcTxVCXRZMVTjTYeTSzBVP1azLKg8038cpIih+GuxVP8O3mlnBQfZPWvCCOmA
DLGZb0lC4ksSW5Y6Mo6u+5u3IiMZJlfLoC+qPpGn2+fchusF3kstKtLJuD8okPXF8L7ha5ChnUDo
VYBxLL2h1t+xKYFrPcXpvri0OWKLrdpHVyLg7S0o78tDNV0ytuFBrX8ZRcdxBquVvzqVCEnrEdJ6
snZMVYFxM3QcJEgLPqxus7GYc1jdxik3CdjRnSsmjYBgdwrthVPa53VpcV/tAWvhzZU70LEbUvic
BlymiOCtQ+M6VfwmP7t1WkrWx89yFEsxuxBNG9v5xHZT0fga8jO5qoUCW3vxN24+kDg9ZaIhevxr
47p2uul5TN7++w3z3k+XOShDGTKjUn65lgLQJq4GMr+kYdNTD7bcf2GbCfHST+m/glKDjf7Ugbvs
RCdX6LzSo46pXePLrrP/Shn7u4inyhJTXIHORTx/xW8Re04TRB4xAPvRLV1DKhmUfgX3VJ7SucCf
MAQTO19oOgNkiJGrP4Ya5QqzJeuKIFlU6mHR/kwXzJ7RClsz43Gn63DyJ+3FxXiwG2D3DUUviS22
l7a9rFRg2kNL0ynnvYlJ7vDAjKEDS/f145bmTeVZHNk6NaisOGeR1dkBVT4pHbYQILlz/eKNPY73
9+ku6kLsgWyoGS/6QcV6NB9cpzv7ZKP3bbkk2fAW6+D51kZK1allQzCeFcBLX2XzZPudm2RhAaOm
NVLyYgLKoYmohPs6cD4aD6OZ/Zn0nCxlr/00iKqUeNF9T0fqD5nxbWv/yn15OUTMlYLKe6v81MlP
7L/Psddgvsuvwfhq6t8PlI6i0IWHmBm9NvuMqpB+WbXMaJPXO65n77+uOYxyj19Ee8PgXtJu+wpb
PaMCgPYHEMhBipV/iFf/anqJrPUc5c0kPJmi0GdGbfoHdkI1bJ/hOrGGpBsAD0mHBTbAKrxy9MPR
nX0L0mG14Jv+Pv07h9rOG3Hb2SE+2sacSUsv9N1E7OPEuvtyNz+z7Q/j3pEH6WwbLSICsaRub4gp
JXEuURtUESgMFJPHG7ZG3dQVjJEQstpE80LIsTQ3y+UczLScWoCV1tfnMUkZQoHkZaTHKXE6OGd3
mGgqx9Ir8mMdgFnApzefPVedtZX0awDSNiIMtUUXVF39jC8/ACEoco1S5zPz5jIQIrs8vlGoKdqC
7T3m9CZJZPqqLFs0snHBfwbRxKAbQRsmv3PF5x0LTF9FnG3zYNEHDeY0LVlyB4sP3Plu/xs0nKwC
P252IKvou/eX1F7OnmkTOBCO9qr6hwCNOCL63C3aVQfMSOW44E/X10os5HjZcVaVqnWUh+ZRU7tZ
pQbV5XH8PFutsg+vaB6ZKlGih5pXtdVDZtoFGpZA1wwIDlRev/wxQpzOhVrwFu5cKeO0RmdedotS
7PprbQpAjPKKGAMrCfarRGK+I4mK6k4r4yp5y2TPLttZmQzqnKLniOEY1dosE26/MEuSYsN6ChCv
f7+q3fvQ6LigGhe53tvUKg1rkeBNtHo7M66A7nYzIrSfaoJsfdnRc5xlI+7IHoO3UT6FRB4kCmOx
OcSvl28ztsoF+0FKDxZkdPsbtBDwZPv8uOs3J/WWdkaHngTMoGNV9dgl/WbMZOD8YKAQgPYsCsYM
LPw8DB/kNOuqKXFOWStQi9iEaGY8pk6W0vnIUlVDsZcatDpuEMiGVDCY982wOoXsFMxy2ZB/bnB7
JeHEplZivjigfcjNaOevhnvrfoEVlJlLRkD9YirIZPEHiE2kDPMe8RmymCKET2vnefmstAQTT6wU
vkZygIM4V3cNgqYR8xCGli/WTjCwv9nilcrPyf/r74EOgv4Vwy6k9l9ig4N5fInSmF+CNWKN3VEz
b/Vob1ooWNf1I01IKkYr7lh4R0mrPYK9+ajyhISnkp2sIZ+zxGSRdZ7oY9WWAigoxjxo8I09Go6w
hNuHhEmuac2Lo1vNJBUBloO+0fpd3b6q9ksxYtWT9Jpsk/QYLaTq5m33DPXkfU3H8TE7ws6DGQlz
v0Y/eH4iHlK45tRTiePhRiEXOWGQXuAWVkzTOPTfWcCnJjMasMCB994VvSuSM5NGqd8l778uDevR
6pPLKMHAFvBiqH61+gqlO6tmfdqRpz50tCBcQ0UZPNtvaWbNaWv3ccxRgWweszc+VVS4cgvG2eQf
xvu2EPSonZl74RHky45JbdAxuZVzbBrSVO43i+JrzxBS6Nbt4sWP9Q3wLc0LlBiCMGucz1vKbhmU
8I3QiAner7vgPuEqDTNWeX3N7hugw3m4tGvymC0ifFK4GaNP4RJERyLLqvhlIVmQVuF6GgueJRyL
3m07L11Urx0HzL/sEpPZhW932NhWYht9j7ksMLp9eONK8cHFXnx1o+6cxkM95aTQHgsODe4nfE4d
Mz2IsvhADqHrLfjY3E0RS1cRJq4FwhQzPxgIPYNptjX6YCDnGM0ufpiwmVROCQotyHgaJI2tNRhT
y3YI9504g5Gwok7VMt5SN00B0Dk0mkg7soCv3DlRyAdrjqLaKZVuVaZOLWfEtd4AJ9lV2lqVs2Q7
kGORH+++k1qzYOyVG/UaC504OesJk8UeCbQDZ9FPcM0BzFVUK1JyzZlP5ahpPxLhItZzWdQ9wNY6
eyUcVWoPFAvn1WI/XlIBKmS8uG8pxlRlKyFucLqemSfMTC1nl0aWYZ6JVF/sknygyLxoQLFhyg5Y
RoAYynPXiW2tylGWgQgstGYVj0OnQVu1DHTVZjabR4wHXynvOkeYJ4Zt4Kg1nrmMrWckqFhbDEP7
+ehR4NH+x3y6Irm3aWfBuUaWC4ppMuFe4SdZmeVkd4nhNuQK9TT9TrdmFtgdNk8SnBlazD1Udl4/
CczIKbGLDtojMsAAcAKZM+wswDw6tj+8R0dQ++cGCC9pJhOC763rCDkJHTa0Um6ht8YvWceHDLZn
ynaGAJy9wDVcF+qDgX7K9twYPC5/3hukuO57Vd/L8jisEj/VM9Q7kKrPIqZ3aX9VxwDPltKieDMD
VHBUud7FXt0yOkZEYwPFVQ2zOB0/S0EDYz346wT7+DoOaFjdG9jGZEFRjBJHIFp2NIOZa70KGWD7
KcCm7iHLozJrCR0SxMKifjOkasdBeWABtBy7p9Jl0UbE+7JvTU8mkXRlKP1ESeHJ7JoOQRWD40p1
DSKANLu+6QY/TZUXJdB4nWjhoFkd8Og3Ki03/d0Xq2RY/iEF3PklBFzG97/jjhbD/OiGG9I7X23z
xd8G9N0Q7g04tuIk6sRBue+0wuQQf1RU/X80xRj95z+ixF4+DdzgaCa7kO8dfU8x8e6IOlMNLk0N
KmmXBCwtktsNrm9HZ4ADA0vLP0EoDxHVmZ+PBzE216wiY4jUFwABeuc6WZKI3ZBLi09LFpYkXGip
ZjgKUuyJZ1P0OlcHq9YgGfMw72807jPI3actjMbd87Ro/eYlnP8mGNXVlGQ8vEiuXMWrx7NAD6Jm
b7Ac9DQZDRHJq3nVDajf5dj9S1O60pGenqlDLTj8o/D638FGMA0fYiM+RW9jdwxPIfLDYYoooXj0
mfFR8H/3F4cEZeTUTza65yZm8KPHfvYSsF+dS/lafy36HEusiEPl2UvA81ViFRlrdAP1biF8PzrG
SNVbH8PiN0AU0WNevOWe2JINWbZ38mAiVdFpNRnhVkRl0vBaRdy/sHsNeeLBcL6X0q3WuDZCYmqC
r0jD+WLWCrBL0pMzoX9gbr/qb1l51rFq/xfvdo7jwWHuJfYwII6DP280/U371V8uUpPq5ksPNfkC
adqXSLfAhQQgjC1Ty8gE1YiybzxcaYxYA8JJV8yClKT2VaDMDUYNIcYBrqENL2OXUCPWLoqXIuZo
T+txN8CWKcBebnfAKyCZI9sQTHcAvqsboToRBo0FlwvwJfb3kIlQElxCFeL+agnwZWsrDf0gw6Xc
ruf1/kr5kpxwkQIKhlfTbgeEaT8lC6JvGCIvL8nIjrstEBMunZN/md1ICoUPB0BiWbesru2v4BoZ
g64ovtDmsOB3odKQCY2wBmzJngNXfrK9Is862jgFMncWiz6Y0aI/Au3p9RURHJYqDi76nTRzPF4G
TAcz5Vxkk1gnalU8xLE7GHwBkxQDIei7ncXnXLkdsrkobbROoibrDT4MRmkxSL4K39vLkh3lncKY
YBHDvPQRKuNFDZ/jgWtyvnQwPIofpgsV0khPlBMz/T33W4EKDGW+ezkHexRbFzMHGsFplXW5O1oT
tX7GVOSxhlH8/gT2x9lfmd3MBDvgdW2zCqyxyyHFdomi2TST5LY07roKepaHG6RsrB2YKSBnw1Jd
29ZrcE7mkniMGz8CWRiy/6h9kd4Nwe/SvelfwXPyMN0gzAC/a8m/MuwlJT9Nxj2obFltifZjzx2v
RdURb9Vw0Ipd3e8+C53O7MlrxlBWl+ah4YdyH80vJ0n4qUTVtwOlsQb6G46h5Az3H1FBHbt/FLvb
atZ8Y/kYXtyTmnGif4B85kMGA6S/gnKfrTOyuA60OMV7WSXfIULRh1c3BqI8ThU1i2M+AgWVtAwV
UxTk+wxaItmN4KkW205qUEJIGKtSkYOKhUDnom113z+DS5VRc60Lc2rmjlq2/WTo1JimpRiihAog
8Qi2/ILN/sCnGTqIrbWJdaBMpuODpMWGy4yK5Hd/FkXk7lwGwe2e5/+n7ydkB45IUCz3g7tuUXkU
FUwB0TCj835F3P9RrqsucWNw4EXzMGVHvYEDXSqLfVVBgB/3U0IE8ZQjN/ayhCvBjs3iDrMvENv5
EnNHuA0erKYVF26A6zOHt0IUwMsHA/+vbM7lfwzQBuUxgr67AEYl+KPQcR/xjxQkehbgfeQyTU5R
yQVkSJ29VjvP+Jjcm84QyUCbF+UvykPR1AfavwACj+J2MMqOlBJiU8eJvdKu1QDMukdu891SnIyI
NokKi7mG7MnUjl4BzS1llU5Ecf6AX4J5puuPe2H4wtagBwHLjf8BwqiFOyFNpl3RxeA0tqaEIV3T
v3C6GqMAuZzoZ6b/T+re96RtktdWsBmMBsNWOmSWFnuFK/XPKPzGmcAVBXUAI/yotQwpmBA9MQ5z
XtpFXmhRcd2aRIEtDiuCXyn9w/uWlmOEkgyWvGcirIRkKtxBoNv6KggOKLD0UAckGOixHKW9Vj4R
7NXlFGZocrLtDHWu7u8nDMv02iKVJGp3ugLE2Oi+A422vEWd30JkN3Z8qnAG1Y5/x8tjY94FKVwO
MbW3BWtWmEmjUHXIjm5dU47Ffjjva+UhSZnoXb5dUpM6weRjd8zEi6IkgLuD5XIRhPlGjPyD9dm9
TEuG7TVHnkBwTqtsl+BBSYlr+X7uHJQno0KpvDLse+LAPsWK+CarSm3BUAn+tKhdftEDK39vpZ2A
lbBiJBuYsyoJTklhpVS3RcS3ci49SszO2JJXULIaDHS2ZTcipw6DnwgryI2UQKFDHdBEypnAOda0
8LAVKoj0F52SNjZf0ys4ueVQByYhMxZQw3kHnUlBS1wYd1JngGeFHxQ2NZsFr7Tbfa1wboFh3o/E
t8BDdV1Yihr2+H4a+/+n6cYBFhLkbIcUF/SzEUWQEuQgb64cLVkhF90y/k34b5zp5HvslGsaA+Jn
euj+1lVBHn62qyLoilVo60DeavDoyXMsE/53mLQ8akTuNTp50uEpvSu6d0M2ORUzIwcewnCNiODu
Chro7zSA5njYnGB0KHivOPl1IMEy3NBSLF7hdsxfgN4KyztQAuOHiAoHM0HzhRmPtHkm4Utacnyr
1Vnh6c4pV0GsVW6dSz1FYIrrpG2EPlgWX7siiVb17KBfAsrPGx9kejhoX8Zp68n+bhFNAr2ZkOrQ
WsU6k+wniZiDFlhIMRQ4I+xZXfh52Vc9AyzpLK6i2ojfzMSX67Djio8b8sdiD3TkDJG2yKIWoKnx
LVJRv4OZqF8ps5jPbsvg7f7C8w5cX+B8DesaQLKt/Lt8qdNCyinV37oLNawVqKv2N/2/kM9eo/p6
EvXlyWn3Vs1srHq7FYz88e28gZaqKUFZEtmLg027BZ2qXVbi2YcKgWKwM4sw0aA3lxwd/ydKH9+5
Qyp4vzPAsQ5x0JdFZdwPbgIZYYXkyRNrpN20g4ZZWaMKQ+tyXKUF7JNmBCQp4cc6etkOjbXcEoyH
sEW0HYCMZKP3Fw9+xDMllOesw7WsKYFodHrH3w3k9FG1bWbjJxf0xvuSMjhD7tkQ3IYOsKjGUVEN
Gy8LOgQiPPkQt9ovHuxVFG0XuX2d4zuJr83DsTImNQvW1wMtg+eQgC8hFPHS6RJ+RtCoKWhV/5aH
pNmeoa/0Q/S+t4Pcz2cgoPjgfhr5Vd6EFv+6PMtyEEo6L1biwsclHfeP5TdZlPKFF64swss1qbXH
zLd/3NxZA5YCJyLXxCSg73aW3pSFI5L+qR5WQfJxXEVRTT6z1s2iZNqk1zjZoNhHZZW2Hg3nNKEU
nwGj619nKqq+craKIVFoKlMaWxYvJyXFuFLIxJwMOcx7t0DCZJ9+mnnr+y68jclqtCPJjMknvLdi
hIjHh7n2ygaKBP6+SO4o466SbnUKBTaTSggHavMUz3/cb2QiweVUvXhCOtcjoCEpdWXaTsb5TDbc
lhRRwzY/X9J6vKjbZomLmcHB+AoDL6He0KEB9Y3HqCj6xES/gX07s70EkhhG+ARrtsV2VhRF81uL
MQ49x2k/EuIQX2FIQBclpOMtiPz7GoClTwUEaQuq/CSm1e1ZFbA89Q7BOxH5UHTRnhMZ+ml95urC
jFHVPRhACSuwhOdI6gLPXUVx+0XwIB8+zPumKk0l0+Uj3w9t3inXqej63JzTpZ2bizD5msuOEvKZ
0qWeCZXujiU2S/zVGAmw6PaVE+76xUdCn9kvwRTXNbeyIbM3MU8RWSDh/CSWCFuG9oms7YO9ALew
yl8iQ4CGSosm9TSKFqASs+SRrg47iH60d9V08h9xTJm3Du4YK2KplpeN36fDSnZPjI542vzsGNaa
QbXwElE+oon3AKe66ENnvXpxMT0WMc6kvRzk7nD3MBPGmvLidzuPLXa7vX76cuJd7WOI2VNfTYCB
BFSwAEufH8fRbhDtDr1nHsORf30iJwWiGlhG4qVzjv/sczxmF1bnCziDAOKNxlFo0GdYnIB9iE1l
WquIxXP/8xS3a1kSp2O3P9+LGyEDdN1EalZbhQaxuYL0XDFUVoXUvqeVmuF/KNtU5bK3o0aICsI5
hNbx3k7jwcwDJEpHL35W4MKMU6UlcNW2npTL2fjlsNAyDEorMI4UXdOG37ZcKchGFkqINjICttwb
iiZi4T/oidOcIdom7xsfJwFIN7fiVMGjoZds+OLsAJ1wx1udTyEb25ICV71mtMM9WeoBBmF1rrqs
qEnSaI4yR2xK0qoPoXenS0i9oJKcTAsp9nlY0ztc+8ZB1c/m6b/6mPtJasLE2wFSnpks7/+xfFM1
7Uip+fqHy1uzJXeVmqOeVb6CiRx1+kGi5PuWI31hwQX+nSz+1SAPesQfP/mWlw8YStL0SoKWhsYs
rw6N10vstJd+wpVTCIOLcChReiFQXXM0y7lA+0paJmx5Ww16zAQFaVslhIED0wDy1dsWS6HJ06+k
dfIkTPHtaU5lhpjjg1HBT8LD406rWInFkcbZF7jX+dPPvi9kxtVITFm4UqLVQq+a0TmUcXWJMXa9
afphrjyUEBL34mbuHy22Dt5DJccjJd6XtjWCNBP287phWw8koh1o0BNIidOveaDwV8FF/YV6Ycid
sgcrL1k7VWAJ+xSF86v1BfX80VcEZSHOcwl9eL4nmbZYbu7Q5E32DNRN5Q8Ainj8owsnhD0z5P9q
N2+oWPa+v408SGdyiU9QIX2B3zbF96wZ3wAGoj6NO+yaSBrhhZMCryd6zBA+EpHDGBFAJXv2vd8G
s0psI4LvrzJk1DTlDFzrB3Jl/5+ZE3HkgbWiJfmz/KuyuhWA+yNASywPt2pCxNfXIs53CvpsaNBO
XfxebHkGuRyBIjn/bZUfHSKMOJiYLkg2n3nOu5ZJ+thnWApSC7YCUzEK49xwIi1obnCaOsp5FHww
T8bwjkAfxoSmQBJ5VRcjpGeFvhZkv2D6/teLUpLiW3D3ipIZq+Vj2MJW/eSawK5bAZ5jNon6hRzl
I7CZm4TkSQpRULh1LvaIXrj+llT4Mpe4sz7IorsohAstlje2vDb5IwjnyWG4SC6efKdVpZTP326n
gGEB5jMcKGWYFs/J+1GGVuXG6UoUxtL4OsoyD/sk1fdcTpLzJUJyrRQjRjNC/6yrevTj6c+DTffU
GjCxNoecn1jyzQzURx7rpolf+C9io0Uwd7p281/FRXx9hicHITQf+nn1ngBn+j7VZctqKpYsWnL4
wJb4IemNKapjlAlpqdnirKezAW8FauYyybjNMqyBYDvk48nq73R+gUGB2JeqVWOB0Gr9RT7uwQp5
sWFBneuCW4wqlDpiHw6GQnLszEf1GuAG4QyzpYfXOoIOQAFiv0eQDtLqIEWMPZvfSsFx6ZD0h2qU
fQVrHh0q5RzKuTENcTjm2rOZ5IeFfw+AHDY5o7HF1V9FAsONoBf15U4f1C6mCf0stnK2/py2wX/X
EFdmjVXAY4OzPqP3o/+oE+GxsWOBbZqIR+tsGWl/lnWYM9ggIXlRi307iN3OKq7189zYErZKAxEW
zS25QBeHLrd9aYdTGx4TcvbiXw50WxTEe2TOHRUZN298H+M/Ceb/cVXqepAdQZA7yGcR8GIq0vtd
2Aze5pUJ0n9mhkuMmXQeXc8kBCBAMvS5URMkCRi9suAeWI6FQAYUGO215wnWXuN+2u/2glpszqoS
xN5YShzoMvsqO2CP3teAagmlGNzG4eh2SEXJM6sUTMmKVH1kkEVxaXgAm5dYtQ+0YgoYsIl5X79C
ct0Rdm4xohQtcK7g6D6xUGazyUTfQ//gWl8236TIgi2a0qDU5QIuBv/6jkqYyBzFQ/EScHKkK7I7
0M/K1HECD1nn6zuOF1qGgX5b13LPTthL4OmWunSyqeksu5yBtG3ECJxgAuq4ckqIwS0mWWQEpxeZ
dUdaFchGIrb6do9xQmIn6XNptb7hSQauP+4ztStIV1Cz0AW0zevaXgzm5uk9Qg6DdfolPWUShbZi
qX0W6brCukY4YS4aT2igCUGM58q2K9Eml50bFQ41Uo+o48U8WRpKQ72o6P0fPoQ1lRjmfzVej0ES
kT6UOatbPJVhVb/ilVhZOptDbXQId7LHzE+0z3eVtrq/g9bgq+VIWCPv1eI41UsgTwFECl28kLZL
708I9zXn0ZixSSSNZxhcKLjtBbDxNn22Qdqm1UftMCNiZE1U4L7fQpjPMX/M17tov62T8ze5lH1U
f5OkY+E8MAQ5lr0eP+AGLiti7sTvg3ZTwGpKN9+5Rdy1fofbKcuPaJcsdOAPG5yt9jKeD9jVJEtd
lOE8CRte647ZNnXedVam8DHUCbFncZPYV5to4WT85Tv7m6g2JAzeJ1dcxi8oI2WojM7mCBjNCQID
R7RL1tEKmiyQ3erwnmM+swZjSh1qotwbC8bIkaQ4nT/gGsoqaOe5rZpUEpdqAjeuRa2fTUq6N5bj
Z0ydOqCaWne9pKiGLWHPrzit+4SDgBae2O7m0URk08q3xDhFzQoi+ZyVH4WBMxcRQ20erU8x8wpK
1WXJfh7rqJzrCTvwUrOo+/w5bl7MefrZ+hZ2iPEtM2Ld+4goneqauhSRzso3ExxRsnuCHqFSBoaE
YZnZJmAhXh3iQkNa5n118sY+YeEykn0/nrDotnaYTIjhNJ2WiwJNAyb95GmBJ4oSANq1I/XrdbN7
k/jYNeGBdylhx4Ny9dfsXBRxBOPnUAocpCuwxsbu4qCd+fUI4expwMRLUYjWAg2QND9IInBasr5F
xOUkfU+cqQO5IPSR959JE5M2DXJhV7vnIZ5f0D5dfzaAvfpWvPup6fo56BGMo1JHokXTnvd/N8Y3
dukxE+lGH/7IdsHEv0paZp4NUzdxiRmXMROP4V4v9RJePe2g5IeWQvL16O5IIEeiyZBZc1LMWdOo
jPsaT+e/IlM/Hw7XT4p1Am2pcW4brCepENUYURyiJ5P9bt6xsFHZDTu0DDfHiG5ttiO/cTFINcqP
+H92MMo+m0Xe6xzJiOOYdauMQc87f4cZKxzbPeCEaVU7RdpZR6fnRi+XhtCf8gv6r/yrNQEv+vsn
IprX8eYbdAI0WQuxukjaeRQvG/KbZ9mdaVCvWxj921MH8Kb12Egskn76Po7Sqh2wXl+xvyut6kj3
zKu/5XaIjUXOktcWpNBl1pu8I2JG9KAK5NLcTOnM1KgwfD1pdNAwfmMSoblngM7qiPUW2zRdCLni
r1UcMVyNIblEF9n1/0V6bhLlm2rdXpWSycKcbc4bP34HPUlVvRz0ZXTSW6daYHIqRgGli97IZF+b
dx7yJVjNDqPx+71yQDZI6cDSPBhnUNPFkTh9h6hZd+EXchiBkHUESv8Ks52Fqire++l3l6n91yUL
ioYOJPB+hFWi8C13/zYtNqS2QRf2PwpGjb670B3vkePZ2g7QTqO3W7G+3yCFvwKHsVJ3E/vJdOW5
TgK3EEG/pwElKm+Jgkp+TcZBb81RiHx7ZEKrEkYCaIqxtUyRL32QbtADWphFU3MODBC+JQuq1/CK
l9MkvW7I/NWYstubPGSMpKPh1UCjSP1sn2E1p0noHMdLk4MVoJ93UFCtm9MglWG049FxujJEKOMZ
zRiXIvAimQsnQTrMf/UlMOTyjjL4EiAfWjBrl/2J+s63JBr5JRPCWde62cdixfOI6NybEHk4/YPj
t1ux/1QzDOq0ekWCTuwu91QJa7tu9RkjvF1B3boZ8zxzMWIw6gU2juPgdCEQAOdQjtsVthU5eLEZ
sn0/6ziLtdLgN3b8n3RUFMRFRqowbBzcq0537H3lPXBQjPyM3KxKz1CHPHAoc2YtuWLHKeqx5e0t
qbPcU9T7h/9Js9qajX/xyaFQDCEdwg2ZIgrYJ4ZJzHla1AIjz2Lwf0JFzO2qwCRNddJp9FxJ5eMN
QmtAR5v7nyaLPoe/FHkrc10SZIAQCGtCRHN/BQyLES4VLL+A8vhhguC14IZRS3XTGghbotfwtgPl
mK/fzPlu/m+F2qBXCAGhN8VSHTK8Bh5lR4rrJtltUVvVt4HfzZjp5muvapg1g+0b7rzKdmdmf4Vn
ND/CAgdSr1nZVvKbrjauzfcli8U52nc7mnx1jfMAE9tempLcxo1d4tRjx/3ELL4hQ2RxipjLiiVv
u/UZ68F/zhJ2nGYJeABT/fixsHqv9Q7JnxAWrQFkXD37XzyzY792ZRS+mlLaBWNBOpeiJW+6uGIX
dewHaBt6qqWCS/NpNc/1B7M8vF1C6aUDqDFGsjZPHy2aUC3aZYs7mKdIxk/uYtfdqXJFBgC2sP7u
lNM5dk4YG7vzdBp6qcyO26lFmtES1rjzQXQZ9bXM/EeqY7AieHRw+lqyjS2sCw+TZoXaGftyBZLC
6TJGoevC7jGrGRofIbrUCSYV/Yq+CL+tKr9pUDJn50rpAESB5/vxvXkWOukG6n9orsxDYX+CVGoW
ApvhZLn/BhInoqSborznzFY5ZMC9ZF3Y8d1yU9Zd4X587eDKMMZhEN2Gq4wLY8X877ly9APsL3xR
zURHKQy7HW4+owshSpkzemPz91PXvTHZ4TEgqzZgZUnDHQ41hbt/FkH62DV2z1KTSkTfWXnZTi2b
Ki/rWlg8+m0DW9N7TN5zL4r63bbFR3M+qzqEfmSxYFrnzWTnd1clvoehxOxpveqBhOe6hn78t4Xo
blXormmhuG8wraliDhXqtdO73jyfLFFX9UmemUNJCmUMz2gXVovELLcCD8jXnvj2R6ZGayOawMqi
FzE1AV6u1vSYaCLLP/XesQhhA93IW2v7Lx2KYdpMsmCRotd8zL2L6Uc5poqhE7y9lwGhwpFNMJla
sJZSuXxMRmQnRkE0tNyMagGv5j3+obD1wLi+P1WMUqQRuaBmYIqMNQIIiXDyfSlN0Sam27U0/qdo
RjX33LOJjQpZxEynfpHWODUDWEVkCrs94CF6yLWPoT/DafwP83AbHHaRLcTHfWCuUpCXFWkXD0IT
XwGGhCjoQYv1F6fk3jldQvCJLxUcrkZhaqJ6zy/VHBifmzi0Qf4EgEpkFCGZbpLv/1YR41Nyvwcc
96tXbJPF7xJ8jRkFnJpTtzkpL793V8o4VNa5YCMkA91BT13lZgHpmY/YYrb5HWXODlHOA5yDMpU3
n8XU0f29UcrAOtIkgxx/mq9z32AXw807VZ11dHCLERkdW91DJqQBlKN8F3uLFBxXSdyJdfQAPGVM
11tRhJou8fGch+bRDyAgMvtByC3d6fYsg3U5a5QP0aCCEo3C4xG29jHKWe9lhsQ/H4jsuin+BbGi
XYgE3Mh/Gzq2goAsMRcB5cJtr27iFN5hOpRwGIt38zyZ582pru5wHHEeIdyuJ+S1jnjIQ8av81Fb
ojBf4GizoZiWumns2anBIPdliDVmOj+2w/17u6hHlqH/5eFkqp8UwoTGt1U5HaKDD1G4Vug+dmSx
7YYqNsP0sjsGXq9o6vWln5GxemfhjMg0VzJkL3rjg6iYIUzxlM/s/RtoM2LeEF3YtA9z/tL14tt+
FKhgXFf1seR40I39nkasJbaXnpu6YM0rr5AF99/Qw9b1JQK3KW+mFVg5UCexiAs9QzmGarQUa7WE
LJm0xdBV5jZ6kuAHnYCMp4mfhN5L1BFqrGVh/PPMtlKukLidQEHcAHzF3mUtgRLCOZqRotvr9sqy
XtSF7jjp2RTaFBME+sAfvvHprgJBQpigmoq/48nKxyIlQqrR0JJOSiIb+k8zpma9/rD5dVbI/pI5
OQlnRfSxWx7a9QtKGXczHcv7yninYh40zw1FMACjpEXrCq50QCOr6WVQZKqFzq1z93fZLQWWg9ZJ
TxrJ/JmF/ORjY0LxlDAEdPvuW71zz2iNqFj60A8HfmK0ewYvaU636rpiyUkc38OgrMVTpb3WkXeB
kwSySSgd3uPhPPSiOasioX9N2FzHK/vVIhMwn56qmnnyvcwHJUwV/Xx4JnAIsd6O7TPCip+90YKu
p6aAV1PoG9sibylmkdfqQMnAXGIQV6grR9itz4s0Y+0A4kh56VPEkOfzAM7jUpy4PsZwbjna8ONe
R66wwaXubnNBOKX52clTRTUmnVro/wNTaQG0C2i/2r+dxB6eK3qk/xtSqeCyAgOpafAQ/L6A1VMK
2vJsMHwcK3WIk3kwYj9QLWlY5iQh8pwNIBixFmXfALErJPPtsZAGKGh/d3u2TAVOb3F/BT4AoXjv
5xGp9abNq2b843e3QY7VGhU8FOBZRVVitmrAxfL/xj4qJBm2gNyMnGmigw+9HBZoIwvt+JF0yAUn
4nu2lebrpJfc8i4mzjGC558nyqCjuhHncHEeuANseieiiBQR11VFquDBPsLKAsziklJfP76lU75z
1kbvYjMJ+SzG31f450DX/4+2D6Bf1b55r+Dza4U7uB93aF1ALLKAtlvhNr1xp6HeNLb6ZQObZszD
da0nw4/KDt7I4wCUNpDP7zaUXCEGuN29BtHOlDkpELq9ykUa3KNVFUbAS/TUGoNWYqMdq35ZJFpm
vcB8wIll3EHXllE0UTud+7l5AD/iPouLeD3rVxnmR0juASfvQD8r4jZVZvhGTrscF2c6yvXEDQhU
loVxslPYb+SHIsdpZHcNBA359jRA1jCfxSfrRGlMMJPx/zzo9egxMRbcXAM2lweceA8mMc07U14j
/izTH1XDqV77sNBt2shp+AL7VGdIpaezCeq9aZHbgOqvfc4pn5IECRGItTkdp97CiGGeirvNtbL0
v37ZKc8zJjemBGGA+a7G9yJQ1LRchlD98FogSC0jGI3EK37x/qQi8nSnQKH+YKr20en7IRjAJxKJ
JqZC8KMHH9jeiuSvxsyadLMHHBSXXwy9aLh5wQ/h/NUkczgAWlHZekdU4UGM4GFQwOl2KYofh7Jk
cjolfRzi93kGjrhxYp9U/KNiLlZcRhuwLPgjeYcoZxdgRbuejXY1tDGTQtYUFBIoDImaGXMxyhBy
+dvCoBTBWu/bEy8GiZFgLgBF2HB4gZwlC/O5b+KU5UI/k4FLbMIAzdS6Phtnjt6ka/JNlXDy5qr4
/wlhyGsGYpvqjp3UeotJWJ3YwvAMTF8SI/BY6/pqlw5qVExPLZFHpR6FIgv4PWrai3cELbPiBzEQ
uMMWPVwn+0LoxM1yBQIMZrxc0lhR1C8mOlbpS/wCNRyIIpHmshUHON4H/AhHBNJHtOdtAA3IOeaf
QuQHjY5mmU5Bwtbv9XihntCQppnE4GdXab4H2eddtmaTasn1XBdph0zKgsS+qmcqgyRyvY45kc8S
AcW43X5EE9DTQunki3aTkKQ2kWYIE+BIyGdv+qR6jwoyFOn3kpSN1NelueNBDl8vuzsSC+OnC6K8
1dg6GkVuuGDgtYZsx8lTMFgNpqhfev0S+JdT6x8dotgDqAulu87TFRk+NAYz001DlGI7YHEahLyH
KKzOSnACFHGgNUJ9PbKw++7p+F9xoNFxSRKyRNfEo/FJeG5pPxGajKyZxhmQjBVydJZtB2qPAM2d
uRysT67x37LacD5K3+mbLfg675JJRANPq6dOaqz9AuUA2qUemJxbM7fmwSGHm9n4TdbLi7ZcXcJp
ruyJPia6GsMatNAs9GKQ4QDrnOMAT2E5hzorcWuNxOKFqpUHSPMV8k2NjDAK95d8HuOCqx/kAZnk
6/ED7mnX8RbeeTrTgaJdrPqX3EakUS28MuQmt1TTrshK06fzfqxP8zFvY40vlOvgW/6FF0yPsCW+
BLP0AVGh+HF7c641ANMiFhJpR/pNgZWGx97REpxezJtoi2TFplFcwPUXif+FmYqOAfEgC/FSGYDX
gDKQF3RFTUrTMvWRl/mjoy9eNpRmW0weDMxM56zLIsOazvXzW/u5kXxq6/eDmfRN6ObcZ3XVL1gV
DPD9oqCy8wkamb6hDPd/4Et8SQSOUoswFGo9129gaCkwl7vocxHUKb3gOoP4Md+P3uglb+QP08qe
akVyEP8WZ+0Q9KATqAmxkm6I3COXZFIhqXoTWZC2PuTrT6mniXxvAwmPD8w5YlBtmIr9aaNsSf5z
Q/JvWUApMW0/yCKKEFkIPSVZwPHJNXHFpJQTy04VYDIhbFqllgCV3E8LSDi8tjcZOC3p5qAc3D6u
Lo6+ZJHi0kJp8S/LJdHm9mk4HmY9f2/aqu4k/Lb3g1IrrAcurtGjp2+tpBq7vK1hBnqNxs7G5y0o
5qYUxxUSLroTCuM0x74DKWPeHBP+5c6L1IKexSTZzCRBvOE9GB1vqQIwuKYo9EIWjIb926GVYski
Z+MDRgUxtmHVZL7eZqFlAkh7tM4jD6xzpjiBJeMVWgKLoOuw0d2d9qpf5ZIQ4n6GTihPj3Ir48OK
5QQVQCQKMhb/MxL1kmJHUcg7ERjh+KQZw8/imdBt2qqBuW4gwsTiuw9m/WvTWEqTqbCzbjvNVOAp
sPnke3gbFUWIw5Tnzo9Z3W7FKJLC0Pl7+0yn6/u98wnU2MLAeLcnsRgzMbA1HGB4VOxGXwyZDkp2
PnHsV9gwea+wciLHey2YmBsFDNNS0YkOa31q9Zkk7xTo6Wid32VWVBue3UnBxtzW9e4UPoymdw/l
wiSDy9npEyyfjOjd2+U2eJPgB5Quw7zkvwMJVHxxat0vUf+iwpi1i19Nn/YjHCSTU4HW56Ii8cIS
SrQzSNTO91KoCkQod/AkzEVWbEkjV29wRWaK6ohtyWKrLQJcX/bfV11JDRHbBuqszqhyRDsEwexZ
Mxn1z9yqWZfs+2TUswm8sVEJQqME+a9j9TmZEEu3/7/+xt6js4zIcGRoFtu0U9nzBd1+Siq3PkLz
TpTNKT7DbFybwKnMsA4jKtPdTL2Iq2A+Kmj+RYY1V78IeiyN7AzDSUNQ7mPIBjQ/mJngJdXP0zXD
TOLkNI1GEPtN7/qNWKMeZZS9aUsZmC4iG1uAR82lHrKGDkwrxY8UnAioxOGD8Xs/HCLAB1EKw/GV
NNFWmttLrpMoWY4HDeJOm0ZLeOf4bsc6eOEredMV0BVQJ7Rvfqmve3nDXE+wlAqxuWT/W1UfyfBr
0tgYHPN/q5yWy357M24adPBrTUjdPh5cRx8nU/mulfvzmDqu9HDpYFKXcAUezwGBoioAAP3rlWIg
Khy3AMOiHy5UEmBU0CGDCjIy46gKOPnzVnfrUDl1VFJwARNc1aHm5kDTlvba0LiSBKCDaOKMQ2bA
pAUomB4lmzj9mBNUxpEHRd+VWHaYxunbYz06B3ndV3ZziD1cNhZXipRhaufIiRBVNjIvtOlAPdrD
MvOjNd9FF7rL+j/3QoqK7fIp1jWU/NrZD4HQx8n17I5eGWHqk65SOGm/qF0GAN/0DvMchmelK2S9
byLXLROZIBER2HURZYFoqs9itX6yjrRRyZYcZWt75oaGt2+zwCGQuYFbPbMzfYu5n6H0MygaU+Mz
heIWQNpfBSiobz2Gd34Rx9F0awWJkgJA6xAcY+Jvl4ONbg6vOCpC5zEkWhs1fy9SrbZSfHTSClwF
Ac0yVExrIcxoJ4wNPJLjIFnE2fx7PECV+8DXMhf6tKoVTlimk/54pEU6ZF8mBqBxdw0qLA8PHZG3
dYie4eiItGEWH5Fgmy2O7KI1B5evoIIecZtOUJ5HGJZLm/6tP9BpJwatNmjIE62/dJK6CqwsdRjq
N4RQ5hoZrTeNSYIDseGZnu6dx6f0lCSWe125KLZOCktlnbXdEElWVyWZk2/Ak6m5yTfZ6DYEL+qE
dENCDBLTUVyXh0nBlObBT1WYFJmZili1fK2xUqifnrY23Kf/4VQY3QjJll1pSltbkMYJmhtBOR+J
p39Zi44U9PypABQGF4HHPrKzZSwOcIU3Nq2sSkycIEuUUJwIB9GXiKzTnjKAWw8a7V1p4i1R4mPT
aiB6pttF+KSt/af+ShFqX/M7tglf7ihkk5nXNQEzEDegOaXX2Fr9S7Ni810QMG1nSWgtZ71yJo2J
dyZQQIYR1EcuknPP9OgayuWPOqwoh4LnJIHkq/QF0W+/QBK1dg3lqY4W7FV/XVCp8a4wgVLckQXU
eEdbijD5ChsLnOzebGvV1X7fqYd8deq/Aq5ZQqaf+7ilblKk8qAdqJCK+rv02gNtp0DeEYMrxfAL
o1z2kxTpSbPkHOHuJIZ72kOtkDgANB0kgomTI1o1al9jAO4R8B0hkkA9DWNJI9qzgae10LpUpekP
b5o5RyepD/A0xFWEiSiGQ4Eczz6TZlxKmCylL3xptnNOXP003cO2Rsv56PZJBcLqgMzUQLYpDNAL
qkbWpqxR4gISVImXp82Yio9/nyOHiYeS2qgaN5Xuw5C85d/CbGtdF1CRFPxqKJELc+iwKfKZb8pS
pPB0/Wvp3Er+wLe/n+3TPM0pAA+Xt0/G4hNZ5sePlwg27GgfsvTsr5a0/MKzFnPcyXWaw0wbNT6n
4mYS92Bvqt7FL4LBVE6For3nE1dXL4eRkt/vixAXjDG3JG0R5Vkpk7fLTvUGDp+VpuvkQ2BoG6OP
pmtlPLAkYwxmSjfuesfnNcTXT5/6LJE+f+yHQdg1kHxDJHU7Ezk15+gJOlT6klo7oXAF8FNMnQj2
ueHfYZCHim9du8zNaxzrbIyggLYBmHGFFMbCCNqQds6HfayZIYjHAVZJfGSdSfO6OGgIdL9kC3fI
wW4YtiMgfIsu2cMND+H/m9VwyjxOE4giQDOaDdtr6wY+SVs8y9VONIOSfTMzBu6GTEF9rZCg/mcA
TLW8G1fyoGF2nQWTIugbLXdgZbwwVe2kxaNne8y11dG+ajyt+53BR9wnyDcbvG6FybSli0ptnWFy
WshlryVRpF2fnGKayoWA36dUV+gVQNUCGqkrh8FdcI9l8CpScZY6d7mkFAgyYpbqY7+HpHUHcvlu
PFEzaUAiz2klc+AVWDEN4WA9ZdHLFuTe85DcSpmCLhIbm/h/5hRlRRJJFu69th1l7KPweTrVBDMx
MGFFwV27UF+rlxRC23Kny2ib1O9udNyPIRRcPPJXtWA9uQUPhzpW8NO9U8cqwhzeZ5dk7etrj+hv
vDy7wZkpsW0z4qSouD00+pytNNmdHa4l4BBHIQTaA5ly1fbXeitDlqhjHKMiwxXfV/bDOoxFdRdh
WZkdcyaB94g+6WgMagNzayPJ9UYGWUUEavoIl/qK4XG+8wfa6GBXReEpUsWH1BoWgWdStsrFPZHd
IC/f8AhZFNRT/eeq7+em4IFJebzzeeOJxwav/ETRWUmYf/Mf592wKmdwYsb3pT/oOMbw4Bao3ZdO
/UAmCe6s+K7+uN2lFqxISHi2lXWgJG0gewWmpKBjO1IGTjrtyllQhJCZuL69MdGJoy7UG1cRXkUa
xbCEFP46g1o32SBUyKJD4UiF5i3wl+9kvUMGUNaAlHDVn72j8SQ60gRsDZeiBmP1XrRPj0gyt9Az
3KSk9HM6tHRBb3gY6lEJa7rxCoZzM/8m0sFhJNpAwLv1leWNtAIpDmCFBJZh4rxiu9oUjn3IAyz8
K2n6S8JL1v9wIlmzFa4dQsirFy3biugn2sft+WkGKiASCyrsB4XS5DB82GG+8oODPPt81Doa5KSW
rrH7sbAqlIp0DMiXBQSVcjW8kRLu/gvYF4GcsbjhQDfk/98f2TTSnDMHvG4El9uR7Ia5VeHgFzt1
oQ35N9c7knWKOfqrj/B1AwMxi8kvSStD2QcYZy8ZPEcQQKQQArxIWs+ogoS2eDxYiV+nUngzvgPe
817jW0th+Jr31anFpsCkl1Bo+IHBuZCGB6aNkN60p/YO9oClt3pgUDieZdM0NAju3hTDPvzdA78n
ml6WBzT9Fy5bYo+r/WpralxdI8OooCSQudyi3PQ9TpMicIADBDN8jyfg/ospeTzJzwDGccsoknUZ
gKOmBsNkAwQqL36RJqUqe6NU5yIHuVb53WykmihL/Zu4c3ikjl5G1t194A5EwAN858I27Mc1ZklI
hb/ik8A22Rr6WBW5X2wlPvGeAf/OnSxdA8Fa0DoAfj0WfxscvB60e8Q2eNiJIu+viS5CkXKpzOdM
MtBOQRZNnndqpbUvcwHk2J2OKqcJtV4PkI14dq2rC/5V4ziNmGkx/RmR/51Wb4Jb6s6poR5mjwet
N6aYaKQ22Iw7V5YBMolZcRleZvssUR4B2b8Dhewo2dvoaT72r4uGHeFreksJc8YH+g5gxX/cLHtG
GDz6lu5tNsUX80A5pAcU1/lmQQe9+Uzqme6u+R4qEopCT+8sE0Nl8sM+IDPi2nJJPmv2kvwXg4pB
/MhqaPyvn4iC0MHMNbtt5QaZo+OpGLWnBAlGLjknmtEvNYgNz6yPsT1Pg/DehURyqZ6/w4/qkDaN
QROtLh01fNJLRaY7H9KPjcLZZtjf2LNHaqeSL/r8UdI22+ST7qgi/n5lB6/RkekwODvkzt1qlbP0
b40lWvBQSgkliX+c6x26NSrWP8toRLqOSqB5EH3QYtKjWX7c57j6M2ggG8pmUgbn/6U6svNGmTP9
seTOioct63EYmys5hmpBwKMuVLGNckG9quGaMK7Ro7ilatNyHhlTkn49m6LyadFbxLuLTPqFaHVB
86fW9kotnbI7ZmMjpVLpCWzwFeTELRnp/cFHU8YFx4CVtgbOWp1OnqcfLwaSWh3KN7GB+LAGBbXB
KjwcW1rSKXmv6F2PgxrjgA91uR54ndVHJ3D37zGTwfH5XwcPyOOxBxJ8hlM0XCinkq9ajNcGusUL
emuGNICXxXJDbAPb8E3Jd/AtpIjVAZQtXGO2s80YTGup1Vi6IxIrbZiYdWwnZ8XxvzQCSZFuFuhU
1PgT19YLrx6CmGg6CbrvqgezOQtvb3A5/FYhJzemrX0bpd//FADV9YY7uXwGmLYWtQw+g3PxPQLu
QkVGQfmAeHa2u9OBxNd1CABSfdIBZAytvzwhMsVGryPvGXqbi4oGXjIsbwC/4EfqQNS5yuS4o/nu
i7lxtf+6/34+ZV++O8FAVlSmJAsZ0gEsn/3AG1rNllQE2BwGrhMBaxeomUtvCgw6pMVt6hYcrV+3
OMBlGa+QLqKLWjeUL6rV7g5+gKEs3CYKi3cQVSulVFP+roSt+glPbqwe6Yvz9vHwfmhz2Sx51o5g
NwefIPFAL/k6xSk8nr2LmHjFD072eR1bokvGsOHvU1Luq6C/a8m+jD/dBa45Vjoe47jj/Ohr4d33
ahMbw20XMYX/CwIJxbKwtIpvtK8djbfA0bH6rAD2Xjv/Pdv1eeaxZntCA0SN20Tnn1rmzVy7/ZTt
/O5/rKzNCdP3W4gikI8lAMsXcSWxmqCobrYkv/ei1zpO9r8f5FTjF51pIg8M6PrbPrKlf0BNsbmc
xeJa/QM7Sa/zCdLT6tonv44KPPuBx+S/ssXCOLNinG33bQ7QfJFOhuqtSOgVO5583YXbgcGWsWTp
NHQmQQEoIjdtqgFT7hF4SkcaDSxvRVU4GJ/wwMUD+MU+Rlhr7vIWQTATAiApBlXG9liM3Md5YAZC
Q/ix73SWW/CM4GoATmIHAwwSsF3tonQSnkAwxb9hNszMgGrceme4jp2U/9c1AZ+i+tXxaL9BXPWr
zKTdbDjyhttpGvbuoxBaTGpC59uVnII3q48bw6SMMklfesm2KMU5XL0zAPnVh9mYxbhd0DGl5bMj
zru+139xbA3X1/OwVCjuMQ7DhFkjMocyXBx+8DX3oS61WG0Ttdct41tA8xrG8191tJA/2+29Z1t7
RnxzQut6JHXZ2rgXQRyW32qnmp3cszyoZu0g4TGnhskEySn2/ExJrXTV0nL0UXsACaZs41h+6n5P
HKihNZHHwYIKc/NQMB39Lvp1H8EnvkMnoooxi+PM7gybB6/Zfs5dsSYHtfuLRXgGG4U7zkTjZBoE
9f3bAc3koAgPFdBl6dWPpeCJPru7sIr51EPCOmxQzgo4rRexW0h8LMQ/3JIvfDupvDneDT35+GiZ
jhwfSnuXMf7pKC49xhwcgQNY/neP4F5RScMk7itF8d4uZQ7dJD7ylCfS/6oGYOee9DA3pGGihy8A
k8BXVVYQHo0oeb48DBRUyTDjKTwuEJenB6LlxPm/2MLm0avp5vQMtQ0VYRBbnchLTam7MV5GHL7s
52Fz3cIzJJKasm5ZM/UpZjh03DnTKZDyEHeZ5g24aTf+nKIavUlqG3xyjLFHZEbygn/VmYUT3lyM
70uGn9+eMa7d63IGPVA5hTEqbWKZ98s64TloiFRMMLP2BFBb0Bi4JOdVhoP8Z7FmnrViRKTpqWo/
US1McJmd+RE9Fe0gmW723uLuRBOWeFPH2FECsgieQcezkDxr62EsBXPKVbZuh03tXXy60c4lLx/K
aU/hr7IF5BnIuNc7KHftSXQNSQ3SCepGBzkO73ahVzxivD+iso9LAqyXC5aozFdyVPzWyPvx4v5v
MpvwJgKkp9tSw3aY/Ouw0j2IyoHLGBPppqriZwBLUltowstZvgnA4xaU7A9BqDdYZHzL08ecqskt
CzvKeFdauh1uAHUBHf5zcvDIZmVDzv+aU8wrSZKdZHYmQh1p5My+lJ8gwrvLLYndMm9I+/WelQ4S
SlzwXypNmwsJOWBu2GqSxS1iKhATG7NzaSeqG8TMYDhRKEYkT89Ph1f3hPC2bT0HGoiKtdztcsIM
KtOw6ebhwc+ch/wp+9Yzsj+ZCNqH52tZLxQiTk9XJAP58PQ/38NH4y5/w7fEgoeO6rRFH8+dMVOC
3bRtoX4YXV627jZxzXRvCU9ojS9IwgrVMbX+lHMuQrwFBf2Bjy25qCkYh84RcMoSXxtfPPYMo25o
Pk7LmFQKq2YY05WcYbv21l41TjQoFsAXK7bMWlRLL/2z4NS+ZenxmRFHoHW3SutnpIhnOOn32Q6T
8CwoI6a0FrwOWQSjb+Aer5JH5WjFYYYJPKkgIgMBGels8U4TfwSOdWHWlm4VTpsubtvd89AtKO4R
13JamcN83n9NkM5wek1vSd7Tcyf2NcO+xqI1TEbnOU2c7oyRGJ4eJE6dNgIlwP1bMgPtY5xMtM/E
K66+vfGeQqAz/CZCUoy4JCZlq7rg5m+1MRD7yitryD2sByiDeNtlu2H6Zosduon4OVX/707TKksp
+l/5ur+9WKjhC6vocfQ50PTXuWDYcN0Ad36QtWPTTNSfHLvtlkkM+O9YghjJZrXMzBTvWlkLt8/e
efcsTHET8MYZYAODCbZIGQk7oBNSA9z1LcgUYJUd47cQaMTFus+dDNNuKLUwDH3ifiHutTKBAsPg
b/fghzTHAO/7n8gxaM7nY4KgbLeI/xAHMfhBbSVyjx1AH6nDilW8SKI3xuBilfGbJ3KNlQTE/ive
pn9Jgg/OWdXSsSDGKbKsDoA2DMLFT1HdjI29pwqIFUqOho1hpaTvMMzxq5YFhirhkaKybnMJaYWU
LSuFB1Gc2f7O3QKZGAZxkEsiG3eULfCV/0kz2JX9vLxqSvXEDSfnZPFFV/Lw5ZcY5c9rvff5SDk5
oN0QFQNFdFGi98l+0uCnCTSj+mXu1tXUovWHVuy0I98DcwHh5t3Sfg+fSjNqgi9yKXkzB/3/OFSa
qhjuyTqXmDsqRWay45MDhMrc9bzxbyyURm1eXejfE5DjJohBluf7V1u0YutgSnJgXq9CbfZfascv
DhX9e1+nQf5vciKlVDE3MYrTcep/NsKBeyMdIPJmA1DcZ3w1sbfFjsaqR/WeIWTD2P2JmaJlynnw
QSoJt5cgmKkW9QHS93/qSU45yRJjrS6oxp9QeqrLhTGeeOj86D6gudLBmajc6VPZS9oWINl8+GyK
5sazcauSOMsAomDr8htbPsTAJNUEAnUQbChEtj63vptL8pj1ZuXpAcUbe9JdXSr9tUfTYmEXs0u+
iOQ5DIR9zS3/gsEX9XtCZKouXXuu64c8TX6MCxrDsFc1TDOMZJMSoRhpBy8GeMDyZd+T3ebYI99a
l2Of0wSeyPipIuSqFjQHAL6Y37h8U6cqmtF2r9oxVjwzlnkpXlrSNCQHTcC4lGTZcWzCumG2aqSU
B+lg7WbNgd/i2DeoNOTg6LTp3Db7fpvYFnGM0eq9uN9PMAIowbPgSkwyHzjoN+4hHxYytv/6TYKS
wikR+p3O81ffzFJiJW6rke8kkMNvihtiGA3N5no38yX72yfjrCXlfW0u398y5YOM/QnFL5r60/cW
G/LNhj+YWaGMVqQUyIQjHehyTzEO6Wg2BVSPFJqEtImYRwpne11F1f3hMblq2QWdRYYgHeO3p+w/
/G2d1iFuMSd2HftwoZVxGQxLetWZ17F/SQjiX8duy/qaJSmS4UKsFGpMC+82FRCrlppT6BYAPRwk
YQRE9CkJJPSO4MLZ5SLM9t/svJRVHQjP92zKk4XQ/bTHaEQlFxHj+sWwNqgNhG/u8pffIsiftlHw
srquhmxMKqIaMjgOWt2IZ8wdYSU0zlOmD68BpPkTPwxnN3ihFkqS6n91i0lDVcVYOUSEPg5doqV4
lFHPFdn3mbelkgWy/iCnEB2vr1S5Cfqe5BV8P19lmViXjjYzuRpt+HS8VuaPFc0AZAqYBWGkcu/q
io4u1tXU3oPPtzy7Rl7rTi9d3hQ/qfgFcRD8gtYjhxvubUmGPIWHJygHBjnPQu1u1z1oAqBMCIqV
kf8oH8opdYXdKX+PocLefgZq4yS2Eqti636uJ1rlUXmbdoij6WtcO0qS28xmO5jucgSvcWzr5qVg
wWSkcnmJ36Z8bcWuwiO6r57euH5T2QQscgw4xujjQqdrNzQCh16wao7iiIWZUYnQbrfBX3kkhV1w
rkgQit74iy9cBB8kq2iPwLd6Lpb+zo1vY0nNgM0dRGdswVop8vPJGWW2L1PMdVgdjw0NUZCdt4yv
Bv3AV71+f3RaO2bO9j+1ePq9sHPliLXfCqoTbTpoFK3IHZ1eniJ2HRK5pzEa/S4XFi/panM1wYQi
RahAEVXSPLOglUzd+ljIX7Daw/IxMwhXCt1d6VxNaq/uvcH6o0nMtfgeiR01F6DbtXYN4S4Oq6h9
e1dYhDrL4byV+os0gMSI2GQt1qfF1Wc+MKUhJRO3+Al8+TsZD0j+p3TD1Hv/k2Z6wdR18i+8q+RG
6uU/29HRWeILKvP6eYIBY2RREFUgBgBndCLHyzCG6BPGMnr6g209o69369Q9Ih0ks+Jd/bBVoU5g
NPbVOa1UV6H8otOooGtaPNc4zYRR40L/skttv+U5wafwlAunSO7Iin64nPwEkFJ5wl8QsuIvwc0I
hRdGQdbN3BvPNyOWZ3Gl9DLg6ihePT38ltVWNH5Gkb2a2ZNQHxkRoXFUUZbK6mOx10bZGMr5W587
0FJj6yblSEPh8NcKH4qr4FOpm5TgrWV9ZeNmTdpMIDKd+4spes0ZWcAVU+5jw9SvtHUZuzBY0N9T
WAFSz5fpsiKTwG8xlknfSvPD2T3h4RyJZfK8tyruCward5r7aJWlm6KBHpJzmxOczIUXBjVpTzHd
5EaDqls8mBLTRrFVFRFEakdaVdXeA+kQXPXqLHcUi5goQJcml4hD/DbyRKB/nA1lFx8nh1bebXeH
puwuqSXMvC9mw64KnL1/P1qpNEEytt7IGJO6qGmNDttn49OOUDlanqoOsY+rWYseiqCRniAcrnsz
lYioOcEqNmJgB188g2nTMlVLFZmkqxDn7TcPGs0WZj8o5JNxr/a+/+SHl4ujh0o7siwtQeMioN9s
gXqqnUO8m6l79rliSfX/VHCGuIcz0IDTHuoczqtKDYzgnXNQWY8Bzez8dINJVpiz33Cz9hVz2z/Q
/iM4DthCDcWfexu4vewhzMLT97sjzWuskh5yO3TjPvCYtcdJxvYZFjUFC6II22AXpv0IkXDR2GXz
US27PIwq97jTmt48de7QNYJ8x4hT4GoIKZ3nj9VQFZyXNkDoReASSi27Il1l8A/ESJb1ijXRwKg9
424zbCScqI7xVaH5+gQksCpdOCASI7cVtmpRUB9DbJYpeJgmiImjGnaS/fc+jFN8ho2fXEDMmgdC
u3UyHRyddN7R4OYlm7bu77EFHFS9clUmds71+ArcP1jMZKOVx4XkDfd2gdNIaMtFyJ6X/x27EYrL
zbU2lWTmA72get6GOnRMnx1lxtJm0bu4C/44voJ6jJJn8JfXxjJhHrHW7biu3nOhEFyCJDmI80EU
is74+z0kqFaaTFEuQFMJKkBtuP3yGnFOIgv+crnpV/KMTE6Fjxyj2vL2BQsHs+oGvL3BDrZpht6L
x0VcLJjSl7gKKg4h/QgoojZOwBCQV0l5zvKb6z1dPlr/tRYkwb7qswYBlKq+eVQIb4zdxRfFIdC1
PlFiABGFHvWxKJqiN1SFjtnRufymmXIJBMxRQmUo8ZprBakCZCXjzFI+3lppS3YBUH6i1/8LO3VE
Ah+cSYhdC2FFuHl/qDPzA/XjlGv4FeceveJ13MJ3rzJqxNQkVZaCznRu0TuRfRGzqHN/gZH1QLZP
OdKuMpvY05dCQt0ucc4q09X0P/pOrpk6B3JLbdVkz7efmTWFRMBkqcgVdUsqtXd25uj35d0oaYmT
aUUBR7exEsGIDTtlXt5jij6Xc5IC2KekL6RmcVSTz5W0+d/oYK0PEAE6ruktp63jR4AubGQSJBS4
x1Cj0wEFcH6ZzVflbs/XEknmgHnoW2xotPcE6C8JXx75SMZJ+tEcUAGA8XSVzzeyppkObw4oVnf4
tFMexdLeuLrBz5qgV0v+39cWZXWGP6xLvO1rLTfl8AddQHt1cc1i4HcH2xizKpS5fTHEccRT19X2
0YpSEO2ju2a44g30/prE1XsqynI3GCEGbAEhpgATnAq6pkum5/ridbGtLq4XOPYhw4mFLtn66CJB
trx0HAH5dnNmtzkhcOuMYw98R3pD3nzcMmzDjAs2IieETOMXx0JhJrnmzPY3Mrgr6H7+3POHWguy
TKedriu8RjoJWUK9HtBbAD7Aem61clBdOmNov7ultS2IHlcH50jwXOxUUU7or9Pt5sDFVKUr7qBO
aT7u2tejJvp3+CDVytAx7lu4eN+Znnp+h9CZ/Y/3b03VYsxFnUuyExM0d7GdILVvCJQHASkEOKlo
2Ohu4YxN066XoF0IOOQZJKQhUwZDP7Itz9IJQje9uMweplY07Txow+Dh3azgKuVWpFt5RwmVWMHk
ivsB8imv1/uB660iffFb5eHupTX/5LZseEkZf7zvKn9kCRgaQXnOJzp5hbf0nYLRzJcozOS4Lk9s
Yllt1q1MHH7Z3qGmtLEjB0DQTNMB65p7qyIw2+fS+ctJRh3+iVAG3KzVxRTjQWUQRga9WZD+Kc7C
pM+BBamZluBx8f2Q0fmV4o4djui2hY1w1niRidORLGbwbcfMwyZu1rVH598hUb7upuEvfp+nmrC5
z0sh8XsaER6zcKOidbNXjSsYVQc3+TgSFluvCTpwLa7HZqPnEgd3id8C6C2yNBafVKDeZcEizdMu
GwFQWpjV5bVMYbtsccBHRmhMwAWff8yY40w+aMAadiRVx4TgvbQ+JbEsFIcj7fs94hLoKNo9L1tZ
PXs+LnlSaCCm++uT+jPSeZgsiRVTkqI/ON2JeSDy5ni7dP7eUh4VovdhlOCAz9y14HdpO9Cqvrnd
cxK9aoN4pGKCgiV/35bSMQePZ0hvP9sdp0LZY21hYde/aUPN+3AhdGQwkRrUwH5qg3iiDH3qxjKO
1LCKx3DYrrTT63tdAmBcsMAf+zEaZdCajR42NN2Vjfu1t8ewVqQZludMRAj9tJM2ROUtVjMKagmr
sGTLiLhzEjSKBq2JJRgN8ds39UcEDmG2xtNrZIUd5dnIhveDvJLNDtPdCc+EHWIV3uzYaQdxXtH3
dtk9JFwD4RLLUdGHnjbkMjUJeUX8mq7TeiF1ng5+1yOqV+OKKUV3cWufg/nkVoN4u3N8s79S6czY
IllB/RBsvxl0tEWDwA0sEWhKceMSdQvwyo0d8onwHqQlpcCH3o3EcK/VlSWlgnbTXbG1/g3hda/u
y4d2zd/sjMLzr6mTDImE91O/Bxw1MlKXbeKw8/y1jnYWvGfMzNuhsTpOM34jYIQ5Z/dWftBpOVD6
Y/veya0wmdyCxoeVJjcKPPbsPfQGmXqi9F6D6W317BcdShdeePWmiJgIBNhpYlW8qUgqQRcjVknI
q9HtEMR/Udnmc5Or54gVyh3iMIl4hxY6PvrDDF+o/0uBBgyY7JhR4FVwKKRnF4t5G08e5HpzBcyb
HxR+Lt5vJD1twM2Usxss3moanqcDBeHc04GQuL3cgczQAVjoZjLRa1WqBnui45nN+y89TygDoiM2
Uxp2f0+ApjlMhhByHUTJMpF2xPaqYJnMOCv+pYeOrBPb6+MmMOFsFNxW0+y33C8Qift6DT97ym+/
xEHvBvH1TFadthN8TeOWeUUgd23UF+GrlXk54w3J33JaWHmAqZ730wNXlbMn7wnFeY8kfmt6qb8j
2nhyQJnYXYDTnDdKHGH8N5CvNaScH5zBk51YXrUT0jyo/4cqvkMJsw1SVftif3CXg9kuTBuW/fvg
J4FtQjoMMfxXHoJR0xexy8zUTT4jvy02EgPJalb/RmQTh7fYP09COmTKlqTagdiW8GCuaI1XSCg7
Vmyq06bu0D1MGWKHZsrSGR9oTICaMIlaf8ZE14B8pMxshg+Rds6j16bLv9Hwx3O6OMb8FD9st718
sj2XY6cMbS7LPkxC6ukfmz/mmC8BGaWKALD/YMkB14h5jfTTnAxgxJZK2pxfaQbO4XxRpdCR5qf9
UcWCoQDk4q6HNnlOl3owX0rQFNImYBjqswOiLdsSp0kOZQpZVolm1DJISU9cY9i+2vu18XXN1tuw
7LfhjKpWbQxtkX2EWuzLunhgHUC8rIdGelVT1pgXnp40yl3van4itfZ9b+rHI7zDtj71sl8dJ3Wf
MPBQtXIJJPmdhPwJwnCtzHyvwvZnoY39kPHSktT3HGpv+R74xxrfuMDrnblsZpg7jbSwHFwnh031
qeEdb6gBBgPf1C54eMRkJDorquLGiT7X3bz/K+rVUA0ubpYb/gz5UafN1fDjOtf7wUx3aDVsWcyH
RayR+Y5umxjCDfqWnzoZUPx8Wl6g45hskLSLZmk1jHDlzbMKQRuLaFBCj1UEAWbFUwafCQSHryC7
Cu4ZZcXfNvN6GpkZeCR2Qe3peNsoZU0rAxsAHL61dJZWNScO3GLoQoZv31Fl/wbF0SpvYLFrkT+x
GrHaP4LLwESejC09ohGvj/mIBjTgvYWIgg3hOtkCLnCfll97skeFH1x4KJnJpk3DYFPFcDWe86xi
u5XcOMhHj7+P7dkLNQdPLfDPV+2HvvYYw7Hm9pISWcq+aV4P2tbKVV1NnSYBO0YB0nsb1vAB4LKq
PfchaBvJvM0eW9AbF3U6bEnrzlTQ3YAfrr5pTbVM7f8ql4Iu8kt8stNEQwvLM1UgW8PR+2KTa++2
o9aGhd2w5dDs9BiSj3OZH38EnHLyh0e83sRKuJfDbRoUn5cHuZw5yQjY4AxtuiDlxU0hhN/UrjdI
Sx7zKIgoabLJdyizIVsONBwY63OE6LGFSHP9/Z2zFmv+S1I6PnuhuJ4G60e60fb7slT0Rk8c2dnj
BS5Jgnz34wMHT0LW3vIa/3voQ5Tzyiuyj999TKUyO05TL3T2V7nBx7JZk/65wUNpAX1/4FpCOO5C
SJN7qlNma1TqieAa7+sYNdhdyzAFbLFzdvIKGGKmldsjyzVBcHug5maU0R+/FDlvFJVKvuQdErki
MDBdXnuedzpm6s9tay8k1VvicEBO1QgXhd42VzDgdItXDKpWWs3osz3HBmi5825UbZ0oMfPQEsni
QSQQQ2guHIES4GTlfOQmrDa0lWjZaLDvPfYK1hxOi3+RNSNs/jw2kw5XP19F6f52lLgBHgk3f8cD
DHqffXS+VcLGvf8GltgCKfnqYKua+XuNVZ5udkAzik39c3pwy3SZ8r+K7fMRRWLLxEigbjSVrL0f
ERQOUb29LaLh8R7J8Q7DK02TVzjkLFOAp6LmYejIMcB3gyJdvWWLb0p20G3Ge1UHvn4cs28K643p
/R/A0BO9NuEl+8eAFBWi2NZ/zXcYMfOx92uspOrTWBHqfKE3IceuGgViMLnS3fipSVq/G2MciHwT
38cBlM4xZgJRBHl6ke4gto+uYneaweEQj/D1mz0GN475EYc/KIaNSN4IDg8pKpYOM8AI0X5ji/oK
hj/SDk61QwYvOzkBROImvyHOvSSP76nPEwtY7He6P16lpRPs06NisY7QW95OQeIpyo9lkbXS3Sz2
fBJBVAWZMd1VTb0tWcTN13dCy0ZZM68QGBSa5gzIz95vqO+xoLf9KgmGbpUo9DUZfBgo/gwG6euG
WW9zjyC0UowOBmX/eabeoRUHPGcV9IXoeakLzgozo8rRw/AhBOQ84fvsxqVkVTAqoog0JD6OsaSL
NiFeYWI0eA8sYQbVYjsMfjG2M3Yo/YBCRNez4/VttVCUR2jrRF1bSGv9cJUktjoCW5PCDiOQYVP4
J28/f/rRMJjnY0PYegflpvuTBZlPgSOoLaBaz+uYA/DbA/psPAKC2/i4SmOc5mYONTxzznrqcrC3
8AkIXXpphid3IxKmpbt1oftPOfFbHVVDGI+k7Q/6UpoI2j3QijxfeP6O/mtYIaJ2/ctaPlPx+6K+
uUo0Zb4QiMetPKoZqMIiGw0+a10a+J35112kHr6O5WxjISv1CSpxszO2C6U8XtBOTa5BHkkJbuj2
TXJN1MeKHAOlUr1soICsTh9kpMC+1rjkymmBKWIj/Ek8KkIiGRro4nHXOxjaIDemlEDvhwtzJhvg
ZG9eiNOJaHUcfUGZYA9UZjURF8g60lfTh25ADX0dVRzDjrBKk6f1tiqpWsV6jVyn74jNyEXURWX7
Q7W6HbQi5TZ0PsrO9f6eRpQBKjkW2hWbAR+5cekvG1Cg8Cacm3seg2tKx3n5j7XHEXn/Mq/1tDAG
7B+IouOAPP7hX8fAtXBD8jJi4MZM3Mp1QeCHl9J04T1/Tpq3Hmp5XR43+owGm1a0Nud19kxX8LG3
yZEcoC8obU99+chP12Yi6DqZ+cfTYGbrNr4YUlvD52/wgMpekCCwgK4SmXVWKJF5kHJWcPDmAA4R
Xt0SNbDAh8E+z79XWhe5Th6teWqFU1SxRYehBJcWpMe4QXjoIKv2joXGU88pOW79P6HMcrSQir7K
xfkID9X7T1OyGWeyFNA5KgulUFM1+DM5X7za3Rm2XVFAU31Ou3aGaafU9H/O/N05VZ3I2wS3Y3Rd
Vw9V7R0nkhbU9ledbTDZ3bCIM+30FmLFFTKdeayJyYugy99APvBOtHm5AmO1M/0KTEoIGLn8zH2G
j8XYACoNMBSLij+NAvocNzYDe6/z5Jn2AvrGtCENlq92EJbFaUWG4OkiTp0/Eobaw6wHivhObuoU
P4lbwW+WHYr7cSLohWwD1Y10Sqmr28tnYoHk2Ra69l8+LrywJMUDpZHI65u242cavvUqSdV7oais
mJSEsqUhu/5fcnZk8Oah2LLBtwpwGOzur27wglvXZwHFONb4ZTh+/S+bWseI6zZ+coLrcGhLlHFg
rvohHF60xgSbH1blW3UT44zBdF0A1eVQ/gnUNTRSPEe+kzMkXOzo+jZyIRQAe2Pw9ya1xBhKvJKG
WJOAkgbMVh5zurrnSxQmQuOKHB5zkA7lgMSbPmiXFAua/WbhRa2cM+NHngWvqjKoum7zp5zGP0sx
s4PXjlJfiqzwQngibMvImPA03Hie59h9KGvDGTG/dvi/tOXV8tMsmtEJrEBj2Ow0Ttay/7vb8L9+
LGGwVcEPb2M0MWF4JB8WH0BRMMMkHMrAmoZ8kfO9slltHiQN3EZcZUWDqyq1k+BaQBqCu6C2Z1u9
xpjD6cvea0ZkQ/k8lUh532CBiL8JNlgJI1V5Plpb9gnlqex8gRVXlua/3wP/tVBcHCRYqpEZEGyz
vj9Ox5cBTDEzbJyLaDC5XtsetTYdZa3NQ+5SFH5Wu2ItvDR1XuKY+zFSju177GcAjQFOxxTFPzku
u3b3ckQXn3WwZtlUPzlWlqfXfv3SjG2lQW5/k4JksHJFNWHsCoLdGGT1XR3dRzdeKoOu1TJGXiGi
fCEXVT1auHCDiIVMSlsU+oGPGaiELn3e6bpObVEtmauWOmqXa0OXK81e+PtvqyI9HMsnJX7uKWHG
OLrS37/t0+68/JqexmbypVO3eQC8+xKWEMdQHLCbu4e8BwplQHRzXq1VHKTQtMcBBaGWNguRYmwC
A+qdBPvWDuDMeIhNwOD5zpbIaYIEntC0U9yucYhzKxHYWDw649s2M+olKO1QYjtTUXJpIfSXPUY1
W2x4IPyEMJ22ZS+qNqVFpr/xeaRXhQemvPUsGYnBukvLPBvmrjNBGoxa/jN7Cbm2De+QFfi5mbO5
PK5XrimQd/y1RBGCs5um2lL11bJSc2eFJfQkiyGzjme7vb2XFOcNtEgHu9Kj3oCaFnJ8NjCAzurs
YnYiVCx9lyWn3KzHeQeOIRAJjpQqt+sd6OLzp6io3GwTDeAPFQU7sXBnKDvHp4eZOCp/sjEivlEg
26NYXnbobC2fxjms9tV9/579F+v6b9be4ysGptlpl9ASTFGdmktlAN/joubS6//qwGdw2CVkaWhj
mydl3/LSgkab+dr1Ed421odh6Jg/sIwylBk5LVdtZuvqVenaqmXXfneW2NGLgltPMxGCcYpkoyg4
kMygY8nLGAGNBRdMUgv/x6qyUg7fOeuP+5t4Wb/0FBuwGEuCmaZIkX+HR0Kzn7boec6elJwf0Vns
F7YULN5Viq7J9rWNJl2NJ4WJB4kFhG1kWigoGYna+V8txHC8WRWUqdVG3ABIyVQNl1rjPZ6tlzmS
A6NCwPlAmYcbtQKcZTODchctNH+j29Zvu4LDB/Q+5hd3ImX1+khNL0IaxzmY1h7ktjDnN3SscbAS
imvomrbqp9sIyWXEDOE9O72/oO/We7a70QXELPNSzLZzcIRXcM63eDktVwLRk6yTfhlamS0qxoCp
QSMEHfjvNWD8/ltbSscNnN3SOf7af+2J4pLMiL5wNzeNwk4w7FRIFgSTpvIr/jjKGdA07P1qmeU9
pSYvKuDH9S4TuHjZ+Z7pBfzuTdebBadcvj07palA3Yrep00sz0kePZxONzGfltY/xgUmZtXmV9mG
P96IHiICeMXHJgdIHkmAya8Ioq4858MUko3kaq/ZBeNqIwt/s4Z1cvGrWW1MvlmfD1eqjij80iyA
9icrJXwlSaqyEyAaFW251NwYpbYTzlp1ENz/LEvUq0c+RLemQCbZ+mOm8/HK8moHuA6uma0kTQ0J
tSvuvz80RVeHTTi0HXDWMqGHt3w/XJW8rH37ENyXRvOA9k0TTJo5FObXUaeFupHPpBwYsn0LQ/H5
gybZVkfzd5fQn+XkXnX8MRjCWVqMFB+GrLmSSjTUiyikZ7g9r1/LlwMNF/bJGzVhpCPA0/HP/nSl
7rhB/O5rfQDVSE2Q4M+U2ab3qmLtQtPxnaWRIZhUu8jquuhT0uruPyZ+slmyAAQ+CywmfRKXzH9K
QXHy/Sf/O+YWYalPVR4rdEZKKj4ccAkInC/0YWa3cBJrAXNxmSUVkX4URVlgBSBx0leppBwQj1qU
yf20xfOW1RAxRyjqoGk0n9ZAvuko6VXjHBdToDV4Zq6X9ua/HxnQAINzSEf7SJozA5uz97qC+IUH
ZozoURA3g7gBy5k0dD/6thkEOr1Vm4HnQ6U4ZDVkhHnroXvNeMGiBhg7Dark4lPdjCplQYMW/ZEw
NAuT6UNHMe7MlZ63RncfF4BGr8JENP7uRaS98HLhPflcmXbGHMUORU/jgCH5VPAwsh8mroJXDDbB
XQ51RDm82XAJalu1oodhKfdRlf0N+N1UEDsXjzCxm9Mxl15+WrPgjE77L4tcwOAhNRkeoDPfj6Jt
B2Ri2B3khCHdXPdGbnsVWFOFLFskKoZAu/dsAZmVTYrWsiCdawt8vXrF+OYaZ2GzIRg2YeJNvrH0
41yY9z4GCDQaAXtN87bnFi72pUBG8yDNDkgNnOvFOxEcY2bicNbmCnQo039v52OIRx+/U8nPiKmR
Luk5G3gbW0TTps679QWJ73Ps1CTZWMc6bAKK441uVrJDAzWGjc7eqVXWJLcAUTsK64Q42ZZUWupf
H5ArZWhV6NHaxFlhpMKQu16e+DAYC12f661p2dgRmroA4+f2kgUSXaHY2B8y7FOwpcG73pofDOPs
WOLGxy2g3CN+4j7mTsOZKjJ8F1FCvS6IsDrBF7e3kz7TzfBo/+qnLz8ydUEJKnEV3Ou/dGivhMXd
VlnteQfZstXYpZ74S3V/J9hRhR7ko6d2ayn9BP7ekll2cXOFPn4I21VX+Nq49tQ8ib456vtRtgMa
n1V7sDZdJlVJ5rmyeE5hnyZhALpfen9HwkyWNsvWUlRmI2Uc+1KydzOvZK5BkKqTNsa8VJ53pYyF
POHKnfriJZVsHeuCnMVWun3w7EGwNRDcIQBTmdvBElo/dpa70X2S2GBCaGSiFtq2aZ9AJBglkSuh
65aN69XQBZqs9gLb9NOJgr1A9E/TTNLegRbPK7p1bJfEc4m/8PNFpuGUBAoGogoQWRRSCflrKLjW
w0wmXxCcj26E1RfKgNXX6tTJF/3mGP0WlEr7x8+qT4QkmIo6TdRNMjMhkoIMCiB1QvhlN/7ReBqq
RORzZj/OHV7ke7HoY80qlWCADPhzeYelJdQWMZDbHtTd2+g7L0oujE95HvUQJI6qWXcN6ZhptP/u
rqBf3d/TGjM3wudqfTTKN6c7vRDOHPewnMHHIhLTjhs/lWH7YzyCo5TYc3xEEqc/mNKIGty8uJV+
9yW51p0yaJyC72cqLlJZNwfvRI1sXPKixXlrZbe9WGTK6QoSjwmfzXnBi/t88j03XqwjS0nu/vaO
0pvyjwbk08jvGzu7zAx2PAjzWS4lkZZVb+bHbAsNW6/G91Yuygf0buStmTLMA86y3RGI/LLc6OB5
Wyi4OK/LOTZPGeQwj/2Ud6Pc8mUjQN1YcGgioU8S/loun0g9t5U8EAi2PlpPCoiPDUWwDzkO120i
pWsm240QNR3plFLQxkjmeYGy0PfVQQ5YqTp6mv7pI8tHCxzyx15QXUrHF2/tpcMqeGFVPyGZjqqg
jSSx2NaBRk8tsL7mr+2kC9B4QlEC96HNK/jIZopv2TBrS7Vvs5sJxmfRbRDURD7nL3CX0S/1cvJR
gL0lKTHA0BBLM2VjuC/CHNrvhpk3sP+UTCfyZZURF1RBruTKbKmcL+avKH1wMf4tk0AwiXfepKre
OEb2IR5NX46pIYYrDa5RFW2TzY91s0tSSymNdkUorqk/Ep61eTQybCvx/ZXHNHC4gglos0pDRusc
DJAAZbF8xTbm4i/URwUDWKo1P3YnsDkO7XkZiDcRLo981IyQH/33eDHATA7IrB3Y1/D2p/etMITQ
xyrx7WqnzaGWtctKK5lSX0f0C+MtCGLVOj7oykirczm3uRcYRHcJqFqqsYywV4fV/j3Ydie76q1s
MUSXlAsRIzhekoFe6gghWhVJWNWmLBlN364Hi+sxw803BnTiMzkTe/GX5xOXO77ONplQxapuKGgt
3dPnO4jnyvjWm6QDhxqBbYSfMlfjbSf8UbA3kC/bafN05KX0PoC+rpJtyuNe5UHhXT1H6P9r5AVQ
ob9Tb2v6teG+2OPAa0epGLU8y7RoxDUMPgo+NhqLEBdWeiabcmGDcAcuWvRvnxKKFZc8K5tAYxJA
SDXrMxLpP8IAmlYUYHEXEOtu1L8me3/sJtb7k8aNYjv3SQ+nc1OK3coLudo03RdSsEU5Vtk5ptuc
jhSVsJ4ci4mnulgepuCTkhj6hblMfVPzUL3CU88AJYThyoeH+G0HoK9nn2yjC7TsJ3rrVEyGV/AB
agNUJrXcX+3Mt7EO5Of86lIEVmEHlIvMwpLzuZa6KNGPVLmIPEMQuO86Lfz8hGTir1ZCqr4vYoXG
1nie5QUndNPWnl9s+h/VQIjX3P3JQXbfZmDQfGjZIFRQBndkEhT20XWtdW/ApDvLwFmfzCgQ2JqU
FaL7A1AvMNZ+FGaTaATh+zvOsM98k5c2LnuTPFjZ9jTBWW86q+aRxtdwfTq7m5QlwGqyZtIdCUgh
kXy/qpT+FNcIqhpOmprGN0RPmm9/sX7nYJS4MhrIIZMVzgLOfkBIlIZer6Vd9hE4nRR9kUneg1yZ
i43//z1eBg5owEY9jTmKYk4QCgcZ7wMlmdN25YK3O3j2AaQQ/hBezHcdMHGqUP51ZgznDUNIg1yp
K4EMyMz4vhkflWI+TPGKXL2LlFf8NewYCFjNLAA9PG+25p7v3iP2qlv/Ql2ZggGe9q/NhagDPWOM
QM6NiRJ9sLJUNWRcmEXIsaTHD3NVsey77lTk27kHB+P5Hk2dxeXmFnjbk92BQKEJpJnjFMKY4KdR
MUh+AsmwQwkg/ADctjXtXq9mt0WEPgrKXlfaQsihydvMq127spnr9GWz48+hb/2RzXL82tndxqJC
fI967DhO1D1HBRWctAJD2iJ6Le1LS6855rZUiLapzQTzn1M+Eu3vSTuXmDTFMmKZoUDHjB7BHGxa
0y22eYvn/QZFuBYvNMeYbZV77iIyksJk3mp39N1NBncQDh8nIi6qnnP+zLnl3DzNwYxYqM0peNpR
ycOueW2reHpgcs6mkDaRUXg4kEx/bAb2AeIaBbEabYHa5Os76fP9Bfmwu4hbGlFL4ey8HgiNmCsU
0BQmFNob8TN91VW5hx6/WoV00vIzXl35WGpXLh4+5xKxc7oqXlFdcNE/s6UxevUcdt4X7mK5RoQt
T9QojlrZvWzlo5ayczvJEG7WZe24VdawFEnVvf9ZbgGBSmZsOOi64sPcW4FTd4QrzRvpHbjNUQas
E1nlc43yWEwqvl+1x/u4Py8jeVBuwKfbyUYOu5sxFkXYTfiwLsXC6VGiWiTk4wLBe+K0Qo/LdN7a
sp+dYvZYeJazHk2+eFiEV59wEZifNmyvj7KT0t86PPo4fG7gBvwKCYMG1IxDz+Ez53BB3Mqkd3pb
Dw9TEyc6f5EQc2fa62VPVivVMPGlO9cAmWb13KLCV3/sGzgk1rPPPuuu54UYVQObRD+eYnHyWKyD
LU1dHHYhlUeT09a7RfV/06b6kVmaVKH0UjIYNx1jPIolIOC2aeMhN1K/LKzxn4zmeTSDE1djq/uP
P6MotZJQ77pYmC9ERIHMgIQQDKc7u+XDcEmRyB5koLHZt3rnc1qJj2Z2VfYqEI8KmJHflcjwHWv7
KnwpCEM1WRKqWSbB7aXynQj55CVT2+BEAQBpJpqSL1kxPiY/wQQ4Vgr7nZjyxnymMw+NBK1O35Os
mMfsNdrgNgK6K81n7+/X9fdGNdqALb7GWkf2GcAzFrzS3wI70IyDamzKCbOHYBPKTakmkBjNtIVa
Du97taTrLHgVMJWWqhf/Kd9vYdq4IuLG3RjvwYsWe2dzNCV0m1QrPLX3Gpnf0HqRTYGjxjqCIJ23
agkNiJsvgkD2lshuzjY0yFESi8Fs/6tDeK6jgnHcuHC8fIzeLT39Nj2619sTwiwbSWK/WU8o+QUx
kimbujBjPDfpTu0k49qS7+mwhZfx4c3w9KsWkt4U5wPmxKT5V2FMKBXomVuH6f2S5DcYdTG4gRJ5
3Fe1vkAI4mnSYiazeW2ldCkZrIVpTVsNCu3v4UhBcGgy+AEO9u/7ovbQCzPDcwCrHMZgs0aKRH7Y
jGcY2PUeuRazLHhXeu3xVv41hktS+kRMzuPQez2ZfD/9oJIqcM2ug44e/k18rQSe7R6nHpSaQ+Md
eKD8BouDc6u8l5wzHMh/LEpq1WnWmdnZQxnRai5GE/cJqwV6ycJwffXkebtdNIumuqvu218YlrCc
DIV4PsTB1c4xGwABJH8Ytgi4XM1ysOMR+Ou66th7UCEF71aQ/IjKrIOTJJuteZgbPPdAj5k7MCfX
1ljcB028TjjcZOFH2dUBZTCLxGd6hvGzrbhCBa5+MIRCw1/B2U3Rw/GA9vXT56j6kV/hkjhYfNQg
jpdEFiavOIpYZB3KADreSTeyNKUZ2jadVBHZvLD5U9Ctk7QmO/onJvOvoCoKtcvtPyvT27GOtLw3
f+KqAyI7NTf9A+mgSo+wH3opgiXENk0S+P0AKG0bRmFQ9oLKS+xlWcX+6XjQimF9HmBuVaiOd5Yv
doPbsWs7+ZAAlK3uq1dPRpHA4n8WanFO58c/7HvEbYU5PhSbY2M+eKakr47SmajrKCLtEAD4z+zK
1XGCoYgkBnBLSTcFsxIuhlw/7ZiwCeib1hjYnP1rn9kzIq6QgHXlx55EYUWSCjWp7rXOIZCJjf4C
I0q6AQsKCNCRdZU50IwdeG/YOIIaugPMKAhBgQNqQy/ePNzeZ41VXb19jfHwQaHzbj18ugW20CXn
jv2D+TzrMeI9o+NUhv8t6T4qbzgKyZLs7qh2cSFEf/fcXvcI94KopQCUT0j7SYTEUmSm/vL4VN0O
1HcWAuhplB4W/RV1YwcX6f5BlVuwdRWw/ubA395Yys+waFx6Q02pHJ7SJHcpxqj8fGuEp2jcvoqL
u/DTDU/v+59Qd4kMy2jhQbJrQpErSJJkUOVhFH8WQdBbBh1MdmVqaKZ+P59Tx+q8bCG7U+xNizkJ
1iLEly3aSHRnnIJXrfM6kunxumL34z7t1/xhKd2ppiBVvKICSx+VJNU8mrumWdASPqXW6n019vtL
OtESgiuEHtKTTMExywf6B1tr+1k7Y0YXFSTqciBMosp1M0yyZGTqlXEbMEGW02KvorEZ69fhaENE
Zz22cV/PRxEMj8wy0xXIuHuGeivw3h4WuS6g9KmhJ0Nfh0Z9JQ7iAFSxUhAP2hiUjXVJfZ0I2SSo
a3S62o40Wr3uEBq0RNZp0loGC52bbYNJic6kR06WOG7PDw/9DqHlp02YSSGzRDcGMfn3LjjXxovZ
NY9PHRcW7IZWDbCXg2F9K4GP7jNqATeBAbOFVpwBgoxmJkaXxQm8Ewoe0kBvGy6rYsIV65gckp5p
z3E8LMyXtWhYscHODyxfjvQbfqh7MuK2PYVbdHMT/Woz1fOzKsI4Q/cSC3avMaufDOmiAy11GeoR
mVB8YC1fVQXZj9Gabe6xbcjc8Q/GBeg8TvYEwP5GOlt489M3iLxFhWsKtqzk934JFEr/6+HAzrM5
fF/YXTqjuw73XPfK2vKqj+CLjoqHU5MD5u2KAm/Uh79hQgcPmtEuUJC5OxYd+IF5LV3L0RGyPhvZ
pf0ajvkcO7k4mT4RG9+zxax8UV/ct4wKRMxSve6YQ5oYDyV7Lym5q5JTMvYfdUNH4CbQHlxwJC/B
Nb0ADOjAtJjLoEQTBKyJPwe9Zxo+bYG/zgkoScdbxwjeXn0UPvNxXNsdyu3LgZSHSEGjtBn/vo8i
c9VTKXG67TCjj1Bq++VP0g8hf7eTq/v/vj1KLZkfodCoHUZAquvMWE3o2uFCE4ydOT4LfcGfLk8a
TVGeBUAX567DU3jyKEwp9JTFqb1sGO0Kerm9JeO6Xz8JwCTXw5VY9tdyNdKOwI0jEv+5zlHPxESe
5m05NUjPmtlxT0GTLQFiNQxA+ORJyqT8pZaHBMk3MAGhhtZVEq8aLhMGwWIxR/i+NIyzHI5+YzZy
X0DYSMUKEhRWXnlBs/IPZoDWUqChplCDyoi9fWXofchDG9l6IYYKPvzIUlCuNeqlzfLftpQsLTIu
oCzWG78ZXpVmjl6G5dw30WbNm8vntrAxuUu7YJxkcbamPQM+F2D98gZR5qS9A1Pjup1oQuHWnOL8
DWhIwGyl5V2X538QjdLsr2YAIqFf0SEGbSggNGYCuAk/FhlBLxbto/dcJytOfQkUDwA2o14zn37X
jqK6oFABBEXW1oCFvcEV67MLLwhnibbuebxoYQi4u+gEA53YcO+4MYWfxtfwUp9iNnppTGnRxKzh
90mDgdKAw6XnIIY/mf6l0ayvNhSrJJQgmyXat2P2GvXxLVMu17yTYMiCB+pgs7Yea6VJmMCz6SHT
6BkDgKuVYAjMliT/nfUJw5IDqBzOmqp8wuqLqOenOm5gC6jdKZvgs6EyhCccrL3JIrpWtFbzuVOD
j1EYMosLqm9LSubZBBilm9yxCXbcqmnuN1HeesptSOKPyLC7lYDZS4r/AKdXrXDM3eLwpHP6qdgi
d+ltJA1GsayNIXmaWFR9kA4ROChefMZZRhFgkMtNh7tXsTBcc2MiMf2cDM3TQXI+VKszuxHRi9XN
YIZfb5bRIhuykpiq8QsV7l+SY14+WW/q9aIfbfksxseJDBidfmpM7J0qm8QSywTTS72mi2phjAq8
3wrXJvHSclE7U6Al+6mB31t5OhHIMNfSPNACj9wto8foNZH80+lFJsl/3xnruaU4LvTadG6NLq9v
AFbZpA3UmrW0aUhcOmNwiLdclP3tkq0illgQ1HKg3NPUQA9Df0Y3nEyuKqkLmL7QUUA2Gk12HD6N
mOi3AgHoKXj3tdiyrQiIHkhv2l+kYCkmPxx1E3DyADLyMWbq+J92QHkVqRYIbKmoyo7hPTEI+MUJ
pvyrdJNChsosHV+8Xb59WBsFjnmrZDM9BVk8Q6Zjvb7TYTb/NujIn2ZaAUXjdrwptEdcq8uIMOCs
U9rrE7uJ1EuWh8P3olK5EhSXGxxjEulP0RPb3Sn4OxQYsZ77HQhWdBhvMWBQvGARQN0eyctfY0PF
wPHOaCg0lq1VG0WSJ0YJ32BkLLyFqJPYRnlHe2nHCUGT5M0nWsiU26w9AmviL/usORLxdTkdI8Mj
tN6OKvcgyLcfsNlWuWKNxI3xhyVwV3X9Gr3cNH2fts7qZ7wFPRB++nDhh53W2cU99WUFRwY5hIr8
sjuF9Fk2zYIhspy8k+xc0ANnm8RuSvDDKnUHfOUKNwBQqryd1BqCe1GpahprvIGlKli2S/NhGFgI
+3MATE17hHim6+APSrlhrrK0Ie26w6I/FSYcnEC4zilSTsWHQkOGXx0t55nNr9ajCHAf00B81BCX
3ai02u+JK8rp7AbXip4O1wt3ZNSz2QlcG8LFQJQte1A0FCIcoj/PxXoYdHbUSykmY4ijmtDPdGBf
8ArHQiUFTsXeYSPi0V5Z7UYLhO5ag0GbBS0XykaEbfiNC+H2AAllLGYduDrpZNUTiif/lC2YGLwc
kL6fK2z6Tzq29US1Xy8X+y1Vury96w8fKQWXlGL3y9AI6+EhHEwrvkijlOo1/hCQtjv7P3gE0+rt
mIcFKAycWwlpFQpfQG3PrDT2I6w5ml/WCaGGQSzRNVNEoLtUy42mgF6WhJ2ByrI2lEke/H/pKaZ8
359H3t8KF+TlmxPmFFMU7tw+p/0WobZPo+olyGxs06rEcyYmcTvIMkAibnN1B0l7O37w7Uawrm/J
ioR82376hokVLTOqW1rwgXIMGzdknpcqgyTRhk/JgUA7SMgdkbQ+7hiCU+8ZTV3PLTGfkaj7uoI1
tTHtoMFOl8BzfQzsVIPPeln85HdLR4xUrqnDxxIGFApqPRoTzLiCOccFmZKIGInqdV+nuhaWshNp
GyU/gMlvZ3OapR2mDWcUIIth+g7Hee3g6Ln1p5k4OLoO6jCrn2oRT6XHQex0BMBx+uS0Fig8QPBJ
465mf100LEa89XfP1il33oR4Mg7Y4l0+T80vcWSVjhYmeWJzOq6VmVBYicu+hTXoLDkvSQYgOALG
h26pw6EXa9W2lfPV9T9kAIDS+kLHLPJmY2GgJpXrSOFH8PUkurW8jjTtnnBeOoLw+oHKrqBPccTI
xubsqQHt7AOTa5swbrCuKS81ErckB+f7ZIjn8UbOzhW79LZTti+yJDrTHwbE9ovolwdIKnq0Nhff
AFxKfclbQcEq+RKG+zzUpcKrCXmkD1/1b3iPSvItOG+3ghH5GHTTauoHcL548I1a9fdyQbhS8m3G
t1CQEoyRV4ZbWWAtzwJ0d6iTeWJgD51YboX9rBhEyDrjm493zYcUqe61ZN9LWqgqbzoXOHTFJv3v
9ANvSfpj++dUoUMBnv5yzJYg5JKnsWf30wi0rywY5l4j8tpDAfMbzwO21GeDIoVSGcrcRYz2ET1f
RaHiveHz2VuEbPltS+ZtvyK/ySKGvVoERp27MvMOjx31lExK6ycuHVuZ7yZOL3+dphd0p08HsLlT
UwtSTgvRyz0HRfax23MVa6NdQp6cW5pbc+u7J8ZybzgAFT/8i+zkYtSMeeUcGeGTyOJWiEbs0i7Z
+6DL9OOBJEaI8ptsGtabB5eEkci5i+8WhlZYxH7TU7seA83d3/bZMG2iS2ZMizVP6Qg+Qt6wWCwx
dciAfeDKOaSijSgTz4+C6h031ka52AtDvItIjfFB9U6rBFNQwjiC6HaQ9nDvSvyN64d763Fk+aa1
ZTFZLCWoLc/j3GRsNNWmlUBSXkuQAvDqxurfABK75jjNCyOeFZG6YlzDk0B3TgbCExUQowG8A4Oh
jRzz80CnL6djUVWmOYgyvfncmZwMk/Xih/JyHalwRYrBtIjyLfPhj+6BnOZJFCkYMZ7EjUCVqGrk
e8V+vFCRQVXcDNHbzMsYtwKZox+hSX8nNmLsg1Ql0P3+aLYZ+Db+9gdQgO7GJlThJcwpOwUQlNJO
O67ePaPM5x9DL45Qgal/GyhM/Bb6YvwOPr95dCkOy3y0zFu6oF1r7uj7p0mgMNxp/lTBOEa+ocHc
VLiHG1lk2M9fKys+URqKe5Fi9rTLcnPi4P+NC8uKbXJFx9yDaNpE0jCPM+B86QdtHtlg8QXQFaZq
Y/W6dYcFf71sTPGJkKrMUd4go118iNQKymXXplQnJ7hYpzp1rrRdZdw4KfNutsrr85LesgMmBcmO
qb8odr0FGhUOhmqLGHIxytBJDiDXH7Ujz3SBvrp7V8gwKNGrAAkN9iz5ma5n+54B7m+tvA5KcFGB
LBAyelMhvwMFj7Umc22zBN7gf/aH+4R6LX9P8lmg5RrSMhRMgUOGGg1lCxZgJwlbqHoR9x345N1B
SC+sjH6YYwhfPP0onoyZgQvHnFSyxEo9tUeVgX7bB0pk95neuDoqBA3Xr3rCWTpqIi4yrSguVylu
YksYmnMLCWME8dXaAfFNoTUfdY0OFmWQI8rsvjDLAkJdSO2mpRC+7xKkv6QhuL9O6pAcDksKjTvQ
+3FeasmdLwYsVhqZzEJRKv/D2PgWc+OKIqnUMmZ76rzUPuCWtkcwufcLlQGCOYI/I7Xabk5ttvAR
RvLMm+DnxAb+HhNDHWmgRuWD2F7zi/33fkMClEwhdH7twFlZhCH+YpboIOWiR3o7ZlfHP9DJ3hKh
snZXkGj1qO+4bCoBFBuj25zH9qMo2Wt/cg3phUQQHlaiXrvV1zXYXlL7izmfYejVu40LkDzbpMIb
wc5xh2LTc5EI8hhISeeWN5qvA7fSoTZMJbWHWn7+T/UxwsdOmg9wxb0RaSGC0eQr5lCAPNhDafDI
uJcyN6RP3IhFUtdgxHrd/Akf3QC40ovjWxsZ49oN4ZSJbHeAmUMPJEFyPogHjJG+g4FL6egtOG9Z
9gBNctUHH93XSBSpDj6CAOyH5lWJvn9TREPM9VxPmS/Mut0hYSHDPoqlYTedfsRIFm7R1gwErVZb
bYNBrKILUWmODqZM7bor5NGxhv2bsM/SVfq9y+oBjhdawlmJ47SBhAIPjVkTmSvTDRC4/vAH69oI
E0Q4qMYcwA25zcncKSd1pghtqGCC0WTQuZyokb0FvES4kxhGSsqAR23/DKJrgjXnxKTX+yf18nSJ
mZLtZW2cR9i+nIWitvhHwoqE04w0sq9x4/as7911LogJd/fNh4xCf+mxdIlDP55FvIYn9eNaSDOq
59iQiLH/vo1b+eApqGMNiz2Y3jYVBZoZ4xjO3nrxXVRmxRaNcbz/1zm2TF915TCr9vJe85aKYTSe
qePxvYWXqdrx9QUf1Ke0v3YgwMr6GLyel3Ex6c0xEK3g+YectlJXJoZI5lm3Tq0LmzgpDCTHt91V
gaixMmPU8qtaDmFlAUoBG+B/JZPsZEZlrbnpMjhYVPF2BNuY5oM6E9EuCzZKq8zgkgKGh+l0JoUq
Pmb/Ut6aYpmWhy14oylQWOWgpjR3jItoQxCSR8LKhSbdc8YqE7hElOt6iEYYfsP1AQ6+ICOb2ncE
0zPcBOFxv0PvfZbW2l4PEIHYCqOI3tLf8KuAi1h1hw6gj/RTwFmjmClFqa4U/036UsL8//23q9aL
hiFkZXATWUtmh5TDjBA/RIB0QRJqhsRcWjoXWQ7/xCM2+UFeaVHgaRSCt4D7JOQkcJND/tyesDPx
gQgFTCJ0mefd1TGnSNF5LiEln9p0RI1wysEt7BnrsCKSawA/7RVeiQmbvno89uC+f2k0g83Vchqi
ow+FV05uwvD2Ex3wq+RI+fflCiQbvg6ga9qvvL0+puWhrxVPkuILn1N9qTzEolxvhro6+T4mBof/
XnrnjF+kip5kbt5eRjrLGKSu+aEXbNvv4xR7QYYktu6JR01sfvG9rTlD075d+j6TuWUKDTvdLO88
3d86GzVd+PmK9wlOr+DmGDu7di534A+cMRlsrKrGc0SiXD1IT+KbYrzXJpZ3h2I+CbkLABGg+Y+5
nZrfm6CRnG11M/B0rreoXFEyntU3o7HLB/pYIfVvr9PpmRp8ffj+lmFq7sIbK6G+BcbTqFRaDhWi
QxrKvHFad8bs21wkPsR7oHBlFi3u4RMhBgDRL6Hl4Uieh9p06SESLIqkgg+UfngU16N73xfwSFGo
gkFKRCqeqJM5anTs7bBxS02TwTXOhOgZrA9TJcFnv4Qr8/0ufN8QOMw/WUGmljRJYmdMktYm/eA/
Uy/XTiZYeOagR6nEVq2j3R/oZdJmjFg1642snaLx4ri8bPbjSrjVogEwTlKvY8OFd5s7u77LOLVJ
XNhNCddKnhenSaWN9kvZ4iZYQSfMIUwU+5b18Px4tJORz9MtEKUXNVKY/75oe5D5bvrUcS4EJ4qc
6bLovCH3FId48h1cIa2rV5O98mY7Nm26djlExCq+WR9htyK5f3F+QfQNiImXBcN4zS1hFMYhNkWE
DINk0DggfVFp4dPvlLbPZDf8w2Sue3lJ0pnJKMf8MxPXr38+yi7TcWw/aqLm3hDc/v10fTUx98Vp
BxCzewhMYqh8VLqSeRdjVPDz24wXXpVUDrqBu4oAZ53OBhyovE1cxXGtfCItbj5syh9utFSuoABx
Gu+A/YE2A58v0Ew1FPQNb1/jQGTm1J62T2hDEYWoJ/snhJ9oqIlW/jrjErHZ2S1SRk/4tT5h10Ju
XNwQMDdsnmvr2oCDWO8KyXu6dvQEqrVnkKtw9Az1Fh92dfvsN/4M6JzCjKmhx4USthWXmjBCMcOe
ABhIbA0mavM4TMP6XFTLBCJYb6hZ8vs/8e3CD5caVFSy/IkzIMaAefo9tQVAgA9z/VXt4oU6TN/5
PWo108VlBIk4sKcqvgkfsmACzrs62KfnTN6+ZrQkPQnne87L8VG+ivYncXrfVb2JWKybLl0b19dM
O9ov+VziCNVwkFxeAzgDnD5wv/h/pWSfQsx/PGviF+QviqAKYCarln52wTg+8h5ghJB6xcELegwo
s7zAS2yeHehSMmVr8QXiE06VUBaMd/abordTZPS+4mqHMPUkEShWOPos9EcWO/ldnFD6Xe2yjPW5
WRB0EOxENZUnjdnE7taErVJ24hwK11T9cbuKKnZc/6tqAqC5ypyF+vExHxMpO7+a3NMxLLrphEJO
atYTt4ZdFo00Eo0pUO9rID96KyHRlVbBMf8VlBNQPsAPIwi15ynxaGVqjMM/cEO1vtd+WOAubaVn
6ydJdsiwg2UJjyD9ATNWjp4Cv9jqPFz87C8BKhh3In14fu615V4NBYQqiU+aT1SKGXYr7EjC5qZ4
51ThefA2pxsaT7/ip6PRrxq/q+w/KsDzbsK7tEaPNGa+G/0YF6ovKStMByehYMpmobLfddZp6KhC
8/tEGpE9t86hj+05oZHFwaKkJBCOXPbyYL1Aa2zIueYo1DD+tp/X0fe2kLSCBBsRjm+k9hdu48Qj
1h2eUaDx0XjcKi0PXM/Om46Xp8l38ibk6IDLuT4I/Aa3uAVVFTzirmoyu4l4a29C7qtDXx0aL9pS
67PjpNNqzSf2gpdmV+249YpxZakRt3ci9KeqarqqtrqyYEihpiBnIkzTt5n2A2qJBXYMe6HJ0xw2
Bv4NVIORlA7Y9PjUf8DBtAhjBFBUYRfS2T1DKTsBJ7IX0ljYgB9Y0LUNMrMA3xlBaSMN4t44azIN
BSXkAPxbvrgfGwvNbygll04ATpImiDDtqfIRa8oG+tJTkFFt4MWWjNaVT94f+bsiQqs0wzSIH7KB
ZixDXjxnXed9YywWSo0bmZ1Nir9TuptEeWyWZ4sSicqvNDcD3xe6zZjzgWJplVQ53eCRZY1xnzp7
F7Hhim6dxcrJjwG7CTqS+pkSoZqDjSUIRsPMWQHtRM1KtWlMr/TykUexkh511i+nvmuibRzxr/M2
ANaIByj+KBrw67q+BQrrv84PP3PPCeZu91mXl2/WnaihVutiIu/L4/FeIQn+I6FETHGLcJUfCmpH
+Ap0V4hqLEJSQ4mT1E/I/UHbC9++ayOnbIUI3uestY2gMWXEhsf8Zt8y/5xciqXxfm/gm2CQTrcy
x9bB6KUA3XcB59/ghy3x9LIPC87dQKLGFp+g4MqHIu2sPh82yiGGDVoDXVLA1O2dfcg/twqhO4w1
XRHBe4TXCGIT7a82qeYopdCs55tMFpmtiUzlce3k58SwkWMP1/RA4envEPkMr6iYW3x22JG4GbHU
NU0L/XfOTZMw8o/FWHTG7YN6wFTNlt9Q/YVx4zikIRYGvM1tIJmvu11KbF4jQBzxVFquMOOSZWfs
l6JFXzOZ5g32j+EEvqwkseaTzCz4q6SKUWZHzrmaysTeaBxtGKJnx19EoOya7IkVrysXdSfzRLoA
kSoRDFYYXJvh/vzvIaW42aBFlGdTDzxbKfNBq5Jxk4h+Q5kJFlnXt4vDwCXumuLr4vY5TEDAyM1n
HHxUf+ecCiJB+SgURo++siwFmrzhSJhHU9o1HKZEKn75R0tUZh1JhWZ7e4pu2jnjz1ZCk5AQ4bOQ
9MaLA+ihVkIy457UGV/B5YrUX2LHCczvdwk3+631pUocGMa5Cmyx8hW8BkHobKcLNATkXg2TjM/L
Icrh+hQalE01vjsFSYY65xmtdz42UKXE8MXPIP6kyUYVfsKLFRFSJQDke9SPB+yZnAsqKEJlQorc
h4FzxemAJeXc190dQw7mOZD+ZMMixov1XF3IdNgY5Ube8/XVd021nXcFjqfL8k+yLEupwnA/slyw
gqw2XaZ8wUuZqX+zHYvPxY4NFX1DfVWQaqJai//ayj7vhzTC4Fjjk2gdI/1oVme02WdgTDufyurS
suXhocmzXMfPF/yCWaFdZ9Rho5vDAQpiC90/GcwqZAJHSw7xxWa2+/ibty0q6TlpMiXeV8XSkP64
JWPmb/bocu+cdkQzbeXFKxR+Y+LwlgbRWzf33UTc2PqabtuMZJVgf4dZwLbRE1+LBIKAWBNgCzhv
4QI67OUDS6CGV3DuhbX2PDfqPYse0eXs0UmRwwIvjxy/V828XLzfnGIgdh5b/O/HfuxeC+H/rP1u
XUtMBAvsH9s2YTuAJt8isecIoxOTZAT1jT+DEbos2k6vmJxzXxeVcYTMe7qi+0S2i3ykqOJxdtHZ
Z+oOLSEfUgzqMlc0zu/XHKDCuXfI2CGWSgCBcwybkARznFS7uSdFUCHscjgaaZYheiq8CBe7KT0d
uj0usRTcs6Lw6NbS405qxIMfvZI6iKIqCww2jbr8Ud9+A5CgyYC/gLCOcg1KYJIY6I3npeZS+rJj
oZMv0YfZYgAsh7XGpVEHWZgBuScWQIs5sk2KN5IJ12JlQM1o8ThB36Q589hSWaqdikZGvw2OYKaE
L189jQ0+6HRpnx6b/TJfJWLy1DPGS2HTjolONaAqy8XBjb2F7TKwodWA+ovVbRrs4MXPqrpZTOzk
88c848ruchsDTQ0O03SJxo7OcNdCOGyaNvoxkviyIrayUSTHiiY5M2AsSxAaHK+Q6N7GR/KDA0rS
b6yNgU+OM6GXbzOPo0ocdOJn3Q8OMdI0f/cx6gU4+y7dJDNsEM0coihwe29pB4bI/5m3VtGusDrK
tdi1yj41qrjAjLf89hF25GnPHNFVzqzUqIYihm+sAcilQOfQhK4Ey1e6MQww2GagYw0dAdielvvt
50//c9O9LiZPIMVsF4OsmyIYlYHRruN3Pi2f7RKiKsPlUeL0wqxvxmNRyIhij9ot0eX/lZI8T/yw
ecaGOBqNwfIQ5+efkAwqrQv/Ja2MnYzp9ZiJenSfe0nWo5P094h1wGG12BSxcfKiJgbKbLSYCC5C
tel/jee++9mZGntJj2reTZ0IvgoKnFm8ucezwM//cw/jHTWEvVNEomVYAaSQkXV71Oxb6QNC8vjV
1DE/uDGAcZ02C2Hh7RneVNOqBICsGB67/WfV+Bax9o7FJNPPtIQpuVYpgaH8JH/OJ/pigasy7JKx
9oSYMQtlkwd6MyYisPhtwxv6QExSupJjj3Yl7qnWBTW6VfuBRPxWsiJKPkPGHU0XbPWkzmq4msWB
8gtEi+YkFcpxZOnWjavsJvtknA1MX/kFM7FL4cOWW23VOpoZa/6r9dg8qlmCKr9kYxc1djeZRFyd
WMAp7y71gjfr6yuQ19sNhkDhC5RgeVNzXX5EWMHTDePg8B3czmdVNta6qIcgIsJwVMqinuKwuN6T
f111s84SqbxjO/wfuQZQm0heVQXRsWFmGexmXIaxJ+doKKiWLAKJo+l5opYUts0ujhG0n3Wodxk2
We+XO3Uk0rvE+hZJnyQN7gTK7FI6j3/3PzUCsFftkn9AGI50MIX4XYceeezc4JcgMdXsjrIu/XLJ
KdN2+MXR+15OXBpXND3QJqDfg4NisijDXPs2g32c9R+NcH0WYmru72WoMBpkPbGn3rnPoi8OhBdu
djhDi5sIwQ2g2NCvARPPCQXf+1uLsdfA58iintT5HFJPtbUxHgeJcsydpP/008VBYy1rkw6y/d/S
ndR8dwARgpAZzpF8IIRZBBrwBCgqjqR0BrYQvqyPLsEtB9gjBLZ/XcLd+y6JZTdCilETWsDCA/pI
cMImxpDwJTvPKS7SrW+RTHPDYphmKSm0S7OpR+glz6qFpwtqq85vlvOI0toEAGPlwWU1YOgRjlaF
y8p8+MPUx0nx+RhBYsaT9CdlSnRc0hvdCXxVHLJWK/VhnlJhxBfG9YwCfNAyZ45jQAgCLo82kvle
yYf+ITgZXu9W5EbDrANVGoSWrn7I11JZb1KoHNYBT8UPpS0DE4H9MhLXDKXp0f4K8cJjRsqGLqTs
mAVZt94sCn/f84VSMH7dWZ6lhLghTW3RS0PZUoE+ncyRoUmvXNmwJBrtM+v4kJUEpdOT6ugE8xyx
XFtHrI3Yasv/8BZ96/HpDCG7PpY18g3yLQ1xtp6j9tztW4p4OKtQN8Me9mQQGZdwkxP45+fpIJgI
T4PqD8juWDPtdUKijpUNwUBopQBJcVgOY6xZJ2K8BhjBqad3X39G/YqK1Kn+ulrm9KBwxhF58Ur0
vt7aeKK6Pmi+xbwAHys7L8QvI8zjpCLUIq4FB+wEIlYUCpdPPJNrfJm72D51SSDFloR+Ao712Jky
rM9JicO/umpYTnN8/M+AKOBbaoREN2uHuuzVklGCCnq6sogS6Yo2wNSodrnj/KFQPOvRKvoYQMke
1cDwFf5v7o8ti0SyblpuDAQ/W6B0vnEAj0rQpTwF9p/3GfeUzLxKEDcKvC8StEQEjkKjr18Fb/5v
wCtTWj9blXdJkfrw/A5dy56GRrtMx+BKlSPTs7l3unbRmHap3fKNOE9v8SUybn2iRc9EU6q67xYA
sPcHypxwGeYO80fWq8NIQBTmo3i4GT8mdDZTWWk7+J3++43hqZpRVAUuAOtULSyf6vsFUSd5j8PN
I80Y3JtPNDMDTZxZvcHAQDU8aiN2zuaPS/eEOc1ZqxsLoRj9AZlzj9ZEMbzToa7eKqdk6LWLrLL6
XFfA8dHH0rDO2DEConCc4uJpK53xOkLYSuft3nPN2O+7MaclqBycmEKHzSEO9zpTknamyi1IDQtD
ZkXFQF/fGYtqkDm/u/zQohTMmTnnor7Ea+TJT7g5sxr0MuD84Kx/3p5gIta/M6Wsl1OVSictvV4f
N7HimmoJkLg7BGRcpM/OfR8cen7xKDUUy0WAFv+Fnj8pM0auimd9tVJvW+MXZ2ZGAFP2lyvfIhIz
ZR6cqmgv6yBuyulh3MGGla/p+ksPhKHm5ndxwOTLwAbUcGbKTr1NK/xS7Nw4lR5wX/Ub8ZvqarG2
Es1nHySj/iApiEMUae6R9OlPjrRc/otyPwwyPbDL5nKUYzPWiymlC8JYSV37dI6ctByhbBzemPcc
0vEWlSOW3wnOuXD1fP4FuEn4GC5gROPMzMM2JaRcpX1lHTrUR1wJoeh4VviAy6cDjEJn3tl2WXuq
HXxg//k7I+l7AoZjOQgx3QXxyXY8Ez0kxBaL5DJ9vBvnSrWtJFmf8usvna+Q5mAPyzRF2oW1ULNw
QDKPCxdrKVjJbdAccIfElUavhI8UwRDkXYieJrOR4cLIdi2R/V3IINkj3cCf6CEmoqnQvK2Fk1Dk
fVQ/8VP0YxK82XQjOR4sFC2CyDJz147FBa8KPfIvP8F/cYE1IF8Vt+MV2K5TDTYfrxIFQLVHEHk9
QM72EK90yrjPImHIbjf3M86j6F0vtnFSF4WyaISh5Rqg+yZm7pUpgK70ZDMWeQ69WqDj5ftnC0T+
iXMjBL0drhWZI2LTnO3aF5xmEPlmzRjY7cmOULPniUXC6bzExkytqdyhcwwTCAbopVanz9BJBoW+
y0iQ2bqvj7N3cZEtKDTHbG5qSTzT6vpO7L9mPJbVbiOV7YfuF/QOLIgP5ppt55Es0GvjsjujqR1d
H2Oq1XOxXqUXNDZHLYZz/UrlXYO3jTiy4AIOvu5mINuCb5tLAe6YASRv2e8LfhXeAdM+28cDDyYL
6FMgbRSJn4Q+OHaNfT9n3deuo6YIyqXbMBcbm1GzZd/WzSIlfsB+DsE+zQRdj5iuPw1D7gkJUA6t
HXRwACDt5HBSQCJZ27joMOe5QF5k/WxefF+T4BZhFJ17D6g5TsrCWOWD8UhH8UVf+WFK18ReqNKe
C6uZe3P2eLRx8DXO1xFqzpl3xu/K5FPUGZGvpSDo2VnO2vEkUpNQ8G8IXpJFYdSchxlAvZd5r1nx
oYBZ3J6yIkMgxeQb+NfBfE8Jt3JYk/O3mP9dG/2qmXE4ZtLwgGfWCRIrc+YTIFHOKAcegU2fgbFu
UVFa5kep3YRUSEbsJFirpyuyOa6QcnW+eTMwAa7MlGRDt/GQ3hG9spumAAm5cm2aOMxThLb/MGok
fUr3/z7BjQN8NE0AEN255s+KwS0ykQrNZxvl/ASbTxxkX6Oi5jfa1LHdOsYybutMOu0HDconmRDo
pac/KrrH8ZK3rTxSlHvRd/5zXm2V99Hysa5dvnht54whSuF8TKmkv+S2qz6Y9bGGCCaXnWqiNgeF
r3FjfbiyOYM7f2hEEUeY+jkyFaw2zp+cy1VVBRcs4ykSBuiovD9kjClxuyDlGRsWu+i/Cw33isUr
fYervOojNJTNu0YCJFjb3iAxsQPHVA9ognjp56E4j1u2ap1Smb5K7uApml1ht5RlvZ86zct+PKOo
SwJfh5ma72uSg2/7OZNwUYBE0v9Q+IqgtXBN183ip7z7Q3WHyRf9LHITY5ly5klK5JVqS0w/2jru
MdaYVSgG88yUer1ztJXPDIJs7T+9RBd7n5WOLrm/GmAIHRPJ8vSIbkfoeVZ3jpNlIhtBLLzSCjBR
48JdXSX6XAON5D6gPAYTtfJDFz4L5CZQ0Wuty3S3QdvnEs2JoBPQKsK9zAxvCrxeB2UJ4V0FsAt7
sANe9w+D8zTlIGZFDxTKIh83s+6wot0ZaMDIJm3YYM5kY3EhbmNMfyrUqD66nSPqkgrIkNlSFc7W
ZpK/RbKivVWXvhy14XQ0XE4QpZ9wLC8eOugTOw6KVu30GS6tJKRPJksYQ2ItTn+Ub1hO2+QGs45x
/ZvQ1EO+QxEmoN9s5CrlETHtIpE1/sWZINtFRXmqs8tWhE+K6Qi6nv9TJ8+9ShcoYI0ASvSDJ0CE
k/EjwIR3veRD+AH0TCb5+1h8qQzM2CvlIu6CxDs+YTB4xH5aDSlGiw6t9XDkYhxaDQjHtCionVOL
Y+eNyNn51fTw/VcT6o0pWCqf6e52R99g6XMEMn4Lh9tWLsSGnj5T3sKK56qO0eeHdVY6XSxcxJrd
nma+J9GUKMNtcQ7VvaoSjb3E8aDd0Yc/v2rHwdY4WEdMdqjglu4VJfOG+rp9QLi432bMx57MIhVA
qTsu+VjU/ETdW+b9UKxUxooUgFrAhxXD6kc3mXqFZHjxnrOzboChtZLmBnVc6eOMUKqoR4rsffYo
uSkHOpKsjeSxMQl8uI7rZ7WRGPoNwi2s/t6aRqgBl7OWzLzI39J4l7uzdqnkNEokmQxehtEnizF8
F38daGN8zGWLQNgXEhfx5nlxdu4I/1zrZpml1t8osRLi7qUC+XlPv+vHcCy2Ybj2ijsXlDhUqWU4
FlkWDdhutHX1xgH8+bdEWh18gJH3+bNL14nz7KSJilgnwpCR5CKMRgtAkwcpLvJa/Aiu5otHCcsq
pETXJgdxVaB0ZGuOB7Ucr1TgChVep0ndNlMZMtzVGO9hVHp/+cb18hbkduGaEhrOewNZFhZmCdE5
t8XkmMrMwaSVsZgMkI84DGXctx8CnYnSH4/PrzzqO+0+guPQ85sdN+KMpSoVAoa4OB9BltXSKlmh
PZS3/Pz3HZtWVz9EjJiHLtt7fAxjLHChzHAu9zCk6grT2fFEji3xG3ChjcGFl8Hny9NouMdEmbGk
XrvFNQsKkMewQQs/a7EyB8jIB2A6lmT9K4+4jRWt4jUIUFuXHIb1dDZ8Sgb0np49l5N6SPSxjgBj
fSwg3XYm2hag4JCm3/675qwKoyxUTeqNE7GMWRftQM3IIZTU83khgejwmj3W/v0s7/MQL/Vid6pE
CL6BiMKU73Pbvi2bxFtOP7YKMmNJ9mA9gVarYSsJHufu4+LayX0mEKro18/+O9hjkC3T80bSSty2
N7mR0/vhMepaYWTEP7x5IYT8InL7ZLmXSd/2jBoLDq7khBtxjo2JpAfY7XKvmxC8dFJmjaj57JW5
JDoNyM8XA0hW53CH0wB93FiX0EYcSKZCESA/PCPM3/1Fw71tutUZRsu6LO4QHjz5x6dYTjo5VMTa
wFm5wb9sRDX4Gw9dTi3xeRnxjQ9WL1k0mNIztbCF3yCVrBEoWisk6hGBuhkg30lMhEXKO+xqVsQc
3nad8RyMAq13uxH2Hwfkqgy66KNFF29hvIIBTix2zhAdT2qms39v/Uv5fZt7AEKekaZ6AsMa8LyT
RYNq9lipbv2e878OLWb9E/qvONH7dTnhRqNk4T46xyRXtGlMGHuIMZBUftWuJOz+M8yKi1y3MJZV
aE2eQhTT2gL8gYJg3eAAr4ymvWV7iixiF3R7rpjXybOly0cwi9k3RbrLOwk2Ink+C/v5pTm/iYke
t9nkyco34wfMq7U3OzHl/kix2QvsaascpuGJ24Fhds94NKljeoe/SNtbv+g1eCCJ64CBzeasXNYX
ATvbKrqHi9JnLXJnfk9loz64cCRkd0qa2un7F0Jk9KnhAEC1oUtkOhUK7nEkeIskTfdARghS72nm
tz+8K/N2atWWEMbB1/9h/kM2LDGNq61DLOidh+ZIJKOiURlpDMb3Tg8sWywVSjYtkQE0o/NqsE/P
yqgmhdEdol08JRT/iiOuz/sJn2rYy/1GIUdhNwdO+Q2D0r3n0AcizKbQhNRSDyHwsopqG+OgFY1l
z/uWTBG/b+eF4yulo03cLkZN8p6jecwCBrwQuf1wpt6mIGC4aqYbY8KZjwN+7Bhze3oxlWdUo+EU
xlJJWAZgwCVpn0fZOWFPZmaDwg67+DexPtRC2rl1parzselAbO1aLPMSjIhqKmdcFkbumRMG203H
eJcMgsR+u7eEOkTaVX2WYf4C0TkUpVUNN39U5AXQhj2RnpisDI8+hr34LC5cw0daUWUquFRtynM/
bG3f3itE3/aRJcago01VLe+i8rw6DZ85qGRoZKI0eZYSunzESuplLmq/eJbx7rLGy0jY920GDL04
FSavwhiF3MkUzozsnzzVAIAlJyzZUlby2QP7YoqN8FFepN4hKd46g5nMVjdJ2edNn1Qk/Ok7FaNS
RyL7V8A9R+tlSRlNuazSkoTCUqshJ3bCTJe2w8d6ptdxPCsCOYX9Buy4vokL8NnCUp82UEJQsKnY
dLLt8D5gXvg598vMuR0BAGtF6qE0aamiyWsDFI+NbhwA4RaMBUBNEaNDKMqy8ORdc5qnjGi9TpuD
rwc9wjdROVaqPFPhCu/22VZ/pMOpRQ/McrZQCoOZI0P+n/9HR1UBRLJtytnrM+bKhYKuMajgQnPE
nf+5iPqjUYO8ppWFngwiT0p0mRcA9MGS5WgfSypUdq4nz8QeEdWMSj2+BH+xslsVqj9NrO0Vgrs2
i52llsRzrxBSSA2thF0+JuQzT01FfAymoPhMZO/VhvtqYpELeJyJvDoY2rMKZnAiNtahwljJsNGO
DLD3SZbRMQ9q2e4gqSGUtcKQiuAL5wI85kBHsl/VhvAPXDk99CQhDOhLlhDsfl2IeJXdhp43CdS4
g1waYhzCegVNiPO5quUR3EVaPS1pMZXDJs2EwAqZc7LVD35e6QQhePIK1PP/dfZce8Xti+vVjAqK
XNs9scvxRB4Bw/17HxcW4n6vLs0Z7sGVgswcOwnma2i9dmXMJ92mC4wLzE5v13HIA1lArzxkhz9n
a0+xZnW/4Op7QKSESZjc5gsjHFT72lRjLKNJ/F2dxv8mttDH0/qbnIsufIKgaxfeKFOQX6bWe0HR
YuDxYvzTH4jZOxDE0Vn/SxpcyfKEDrYaYfZs0hWDJEwwi1vDbIm64ZDQbmEORHdVvEn9F9QVZPPV
kVbGui0cFC/hF+1MNt4/y8Oxrkj50Y1TpFSqXT6biclpuNmhNB0q+X+8wp4hIiAy1EFMP7r9qlnh
y6C6gSBFupKorXbuE78DikHagIDq9vYmRiz0y5r0b6ZAjTkxPshKI6X1lnvGewVnD32iB9UuoB2m
QWoNRPTEtB0yNnYYf5Qj2p9HrZ8pHUsPsGbM6KOHfCxiiVQwWHFlAm98luqG8bgG4PpSjfWZ84Tq
/SG0Xvkk+HG8qd128Kze1K2q911tMgRxQc2dbxtHQPib6zlHoeBj903cVMFLUqMHOgZ1ZqOPFZfV
ztMAZK4mOyGDzI8BwKLIx0nvCx6MSk4PJLXv1fd036AzyZOTFsXAfM0epSrmjKdr3txyAkRVzT3h
WcfTjLRk4JVc/9SnzIQ+FBxylFvl6wAfR1XsG7thKbpZld+I2xkPH1p5rH3YbZ79y8RLqv+m3xNK
jRp5ovRZEBWz5lYoF+asGJTOSmftZuKc7MRyhc1Bgi2Hu3taDsq5Rh0N6gNk0vkATo6qRCJm/LFX
exf2mbWg7J+GOo5t6d/YhlfZpxb+QXeKxu21b/xfHTgTTT+zqt3G/9FJaJKlNLUHOg8Yx1jWlpFE
MRGnZ8sTX0oUTKTenlOhmkOFyhYTpevegvbPlSi5htX+ZNk2Eamgddu8khIKwsefYghGRXz0v3TS
pO417P+8wZZKoNQqwggVXFMhcKdbSO7NhpoToRYqak0ZHuA9VgJ3wIfpuk5N/bJOsBX91oRyFNDG
e0FY4Tztcl3BTSYhJ+kET4dTq3gJkI4yMPKV+T4hN81dIB/OwUE4nzWjOFZYS3XLXlyCqnySESA7
741i9SjMY69Frz2cxWfoSVKW8Vshju17qNMvg16nXCF9e+j04I8pKSod6f6fU087w8KzOZWfeOKM
TSpFl/AF6SusraM/DZ/Lg98MfPWI+ZKvDlpQBt6cGP1nCzhIThxwfDw23714VBIGCjJu4xK0M75o
8/L1PfANSQuqNbsXpjtLSaPqCezr4yAhPFoC9HuM2iIgmU8Xr+E9RcGuw7c6PIxrQrIaUrYiFd9A
E3YN2fBXCmF4JR4BIM8fbfmBwDUlH7YdP8Rg0tkdrOFeOGZdw+Wx8hez9MVTlqADjFtdVZsPL4NP
QMruQ1/Jcsr13geeaDEULayW7FlIAeNpqCySZVRwv2IubercTEB8vp6Eq+6rR9k0184cpkBIG8LV
k3ja6q4fDe6ICRID5VV6XPGzpbm+ExRT5OcTSxMEQxa0U59Wpt/vgCFMNF+JA4Gu/y2OjVCW26yI
yfc/ww5OKY/0Mng0L8c1NPZD+EboN3i0NddsZEgtCYtsjH6C44vB1iMPMdbGROMRYt44JG95T3+W
K+eS2jAHzBUt5/xSEBzLM956L3mSBcGuISXpqkW/Lw2qlysrbntgduC44VpeJY7JyIc43mJnetuS
hDnNnmJ6M+igv44ju9ThJfeO8fLrtBBKgEhZY4Gi3ZhKux5gF81nOGOf5rmjUPUHIuQytftYxWp2
LtbtQp12VrLP7+2Hn7V8rHAAqjm1YVHKAmoiXl4P5twWmPXjSFGpNrq5PLvYGcCsgozY4jgwzLhW
5cwtTj+GI7SK8EdAynmBhZ+8E4e4JNbxip3f7k9NZmhACQkuVIxFQ0q32F50qRWQQ4+djPQBNgOK
m8EO8z6KoAO02i3fP3p2mZLNh4jxN/0D6xnvUg6/mSum1hY0Gz1T+s42gf5UDeAXvYrr0KZPADxZ
RRdEB9IzlK2C1IRDaeW9nnRU8tbPlLD8NR4cqgv+ZpYRHp3mmQu7Jfhw8Y8BqCldAjKZBkaf4GbW
vdOI6y86EqRDuoD8WTqgj8ueHqMPsjy0rbLpdfkG4aPENcr+veoLuFllaAAPSbUmeEtDiXXqV3B+
VLIQIxop8a8S9vOA/TMFG6P5QHrH4311F74WljXUaGUtPTYqNYEurogWahYQGnYSBfSR5HjvmpAN
PZIRgezQ5yV6exFJax7cavsgZ39pXZtfOXMDlx1LTfMPA3Hh6H7xD1OpEJCXUgXjJ+hy9QP1XDNd
hDEsGaKmQEevJmVNKyTTP/mhS76VXVAEecEs2KanjjiURGmShoaqCHvfzGWxM60dNiYXRLAAiDwO
PDtqB7rYFYshI+LS9UGzQNnSKKMU4JRbiSpCqhNMNTDgplxhFK2z/sw2VNNzI1A/pY/IbGe9Xb6d
IEJOGxOsTJZziB2fmy9o19aAePE9gVd3PYNAZXxXt92mulbyEcyThSMooUxxkVK0lS5iw3o8qmlF
KkeIr7NRdVj7BhCpMwC4O6fTNYkwwDBReeCnlKWX7B7DmJFoee4/6nTPc9DDc7EGkZAdiNwsfh38
yCi6S6nrjgdsw1LDrS+lBWkp0DhqzPh3RWgFh+BvXFtZL+88C21+/+1hkeAc4xltHDYjYJtFDGg2
OpyGDwDkHZy45eOqYMPBg4zilbc8niU/VkSYT3NQeKHh8UcnD7ypwevNAeQ4lQfnmlBMDxEXhOq6
7ws93gE2XApOyhvPcsd+bHkuRaDNt79bWDMxmfk+WbkCUXqwqkYrueJFlHRj8XVoUEQUZ8JwUAqs
WsWxh9d0ZRNyiOuB0q0XMjKLK7Ap/qv0srHUkry0QKW77h5XsiJm/Hh48fhOd1ZODBj0jJaVoivs
TSP9OkvYZdiBBz0jRlJKvZGeh8O8S0yzq0fyIl33wlx8cbtHVltN+YGv+MjwicqfcMIEeou9ZImG
Ld6f5yMxdcUhbBE5QFSMs1rQRs6YDt4GJPEqVq6k6eRj93Ng5cH30oqt+4XgoGzgXdPKjKqFo6T7
zaGY0ap3LxMojbdeRXDDC2oUYxsOUu4XqciHFoA7HfMXGZiVyrt9XmwMLGUEzdF+xL+KwsL5k3OD
yl0E5ebYPsG1mSmujaNYZ+Az/8w4Qy05rxCHj8kpshT3bwL9G/gcO13sKcTd66cBmluVEQY74Pfd
VPiZgZRbKA/gW6/6BA0jmzGQ9qJ889DKC3/EddmJKlb1szbC+K9XFru5lWzB+UPoOaXfyCTNOKwX
wNP688QAgLoV70sSHeh7crEiqHlOCnl5NIpqhJ6LLHTVDP4vy0wXLgX1DRCBoCBbkoR/Jn0olGbh
RNAsBg2Ul67dF707wBdXBaC1I5xU39nUHjB4mUUlAdmhrbSM9+jWrBziwTuGJytTJHOMerBHnjxV
v5DhE5UOiQqxr0rMoqpJkaa3Ug/GCaWwmt9b5XEBy/tS+jNw0BRwSSuWHYjoU4QmthBmVSkdTGX5
mEwcuw7nl7j1HUTmakzRG7dCouTg8EU4suGzyP+LNQS2JMw918RharW53kTOjEFZ/FUYmcqk81sU
i5X8TXdSnL/O4msH2Ioynw2sT6JKFqBbPT7XBz0uJUcUxKtFwaMwOsiR1FqRIwNCkRoRrLXhdEeD
yZVmHwCc+IUNihKb+WP2TKCYNjJcEhVAPnEqoY1qz5nQuredONBH3pkyv3eogCVDVMu2hxcUb20o
2VEbm3WyFJfpaQ8lySz6YmSUS79LIhk58IpOR2kqGryXNjLiaSuvpyz6l41ptojtv4TQi4eslTXo
wZaeVxLbc3xGWV2tQZZzKz8Z1LHFFsLYg9Bj11fF1B27WB73zDYpd5IVGZ9OMY0ZWzFEA0s+AhNg
clzfcB3Fbw6vfwv/ZAMlZttIMAlywZoDMNJdRJmjMqGxVoeWOIAb+nvK7rtOmJYd2HJVMSjhLyTo
SlbJdYxdgjTU7+axHXoJy+x9r/ukAt4qOWlBfcAvn42ZM0gR0GVWZjaJgIOUjZPphH4ZnMDESynJ
Q456N4TrSxSAMVxS0A2lueYfXs9w1SiWgUx0UoHgs4ClsM04aSPW/deoLjxV3l6kDMXVkbVocmAq
QollvFlAE6FbVeopxngJtE4nXObDhzXpofU4Kq2yx+sfGa0iKk63K9gexAL5+Hor52/MEw4OLVcD
WIk8WW5eHFlUpePKfioEyEVIN9olxSb6E30jvC8c80DrE/ZChZglYNO7eiNM3JBNHXYCHstRVGd8
ip+2jX8osNMHw8XzchDpK08jMFvld8Lk3vmggo7tXhEhmohMKoAXcUiR3WkwCo/8SpJh92DUOTxL
dFW7Dvdbr6a071kPmAf2SxjHo1lEUbGXWJkCrXDAM63CB8+EGn9SvhoksDL8TC9eyuaqfmhUn3d+
ACZwGdh8U3+MRzqbFofmhGPTV1iRooVOytpYCPSHipGGsG5o0zTsnR+BnN+g+pJOE6R5his048tM
A8XiXsUVRAmiZJq5DUcoCPXiARam1jPfX6FVX6810h6aYosKbH/MLhthmRVGqcPebAF+nIsjo/Rs
EQxUalq8QccNCQT4+tpxDTdBJlb6YwCrCJWcqrPKp53RDLsjyjQGIVC68fY/OMeVx4Y75dtZE2Ya
zSBFZjamZibWcMM00AQ6gd3qMsKdBuXgcYsbWoGWnRK/HrOMDlfzjFQLAAaG/eeXUnRl1zR62EFX
R5hVBgcP01TCEg8/WM/ZFScY7b2JEKSKVSph93saRYa9fCwBArIOMAJoRE0UtG3ai1k9wbnocrj9
T2oDbEREfzmzFeiOJe8qEon5kbzI3+WMeGJ4OFNNiIVAfebRUQvrqeTeh2fAUSeDGFVcDY6ILjyS
5ujE4Fwofd0cQrn5E7pS2QzNO+M4sFnP+09BvJ93RNhE4cEEW/WqQwcSNCeE0EAGbfrvdJoVm7/c
pZN9gbZQP8EoQe+RZAGVWecfX1Hlrgc3PHJmnL4Z0iGLVZV8dzbuOSI26o566y7Y8BqoN0s4QcSy
wFncxT2rTtWgDXFW6Iohf4h2A693WOXwyeANevkvTMJC/OvFGRF+sKJMxukKzJm619BhmjA7sr1K
ZeJasWXjFrG+N5vCpA+PL2qOsAIkbur6XiUfUYEsonosmjxoJO5TqTqAsLq9Ru1ayUHsxs49lzLG
aBrld7570MZc+SbMdW87c2X1a1yldDKrH2vXO2qjtmJWu2hALyKa4qYhGL3ExRkN5K5FvftSsrbo
OfXt2FtxHxuKqrNTyr86jL9quOOtKicCS6qSb9yHTkmd7Y/Nxwp4KiiSaKoYbSQQNVSMmiD/Re9p
xeqWf+WPRayKIdR/BsT4VTYIuC3WCsCRHfnccJpSWiyNk7iuW3/c312FRiEoA4p9XTirZA5V0i+y
nepAR69uJooU+7kMrNlTu04VYTKaTJQZHZOyFwnonZwehq1TY8/USTKIr9hAKqx/6HApSAcZU63B
r9EjzrzZmupAHJH3cFfw/5B68R2xUaTb5OZiIMguq1vqYI+OxzotMDpCbQ4RZFHubqlpwmC3U0lF
PapE9ARQV8yXoCFh4jbDks9rnjBFhvcx2kNTMKNrMV6Ym1NXX7iSqrXNpspUAuZa41eXy8lFguSe
hKjYbU7tsvTrsVaNO2vYHgFr/8Etv8I7kfzHXslQo3ZQU0WzIMjAAThF/s8y/nj0B5lKUcxHtkZ9
XNHdsUZGi8tvzGkgDp8GvidVKukiJWC4J3Q/491QMbirCPK+FXPeRx7gbri4Wtb9goGWIKoHMMX1
9soaWTi/fVyj8aytIPjoEPIt02u5gYBPKcJvKKLL7dt8XzfNKV9SQ5DviCxZr3IoXZLNXvvQHA4j
B+wzDBZ/zP8IMGKqcSPJ/jsDrQQJF0YNLJbRluitW/FtZEGKkJXRwYsLpPYs2ixUGe8PJae9p5wN
AMVEDu8fUhwfG9hQlY2vxYou4hfwEeSXCjedWZpTe+qtV9KxSEFwINP7SdTEP8sIwRtXEi+eRIAG
7Z9Q9fECUxW17TSXG8nOZ9IeWZUMUmu2cSBnTvwWCcqY/3DHDF/KlITS/k7hYeQ/VokZ4TUdgtYQ
sO1tXb4bSPZdVHgd8D9Akv4MipJo8ffyJFh+3ZqLmRI/P9zBQWi0pI6fHg8xucaI/XFq4sn7iTfc
CK0VzTO0LhwFbd3lO/xEHpv9MEphNR22nDihpxxf36VLyoTx/gdp0A4vBwJNjVAllyIPlFTDg5z7
gAnItJ5Ri3fQAotJ0dmRnovSUcUoiUC2CdZJoZ58QlsVknDws9Fjxf04lijgu4/SOr8EckU8CoSQ
gUbJxoGbGOYSNFb39l42w5r7y9Hao1HNTJF/mcpVyUxkac0RucZhJjd19Z5ZYYSxSxqDzZRmXwut
2P/cYx1wseBWCUK6TthjBzEZqK0rln+N6IPHSirFCdbzEm6z8SBK/P2IP3yx0x7dRaMJHkRlVtUO
sgGG630ozolXJ5a9dcSdd7dUOfFssbmvrOyj1XHVg9HTWkHQfNfoImMyFuDbfitKByNCu5p5AmTn
x2uINLbWmqO1iNoOq6EWYOj/qr0qVOTew/DsY6AWElYaZxv2bbiovlLQRp4pFs4mDwfSdYVaD2hg
HL4plJBNE7G+3bPxeaEoTNkKr41t2D8x1D8VBS1Hd/53leXJhQQtsBBfYp1J3mfiW+Da/T4gu+H1
Soc5ig6qATGAeCYqZx3S9vvArzgKhaPI/hDqJjsA8JOPhPv+XZIX1XxMh0LLqs0atf+POOrinYDU
kx1zA93swp/qdNCUUEN2iSTc/RvW0h8ynch1rYrmrpaqO0ScbYHqrTlpDr4C4cRyf7Z+eeOr94+U
sS2fzf89YkSMs0ANVmuAgbBYhagrveDLavuG/mpU7MxsjksyeaOBsvR4DPYG/NThLhsbYiWEqWkE
CFw3GCz/Zk5VGUlxWAvBvjBaG5UOiaNPYXfHYadBzlbwBIUzDGMh8fMZQyO8eSRkChIQkce8/gQb
hVtOqj16oAncydcqJB3v5w89ShUPoJ4eO5Vrz6wYXPtyMKsIHK90PiurqzMhpjBN2EwbblrRVOsb
CESv0LO9LGVL9E5WRw+w9Nu/woARsJEzGH5+cTm35WfbvpFKxi7jkv8Dfr5uTD8ZNgto5Jhr6i+2
m8ivQWD571XEIwX8qLcxnXTKseG+Wob7N2FrbNMZBug5LVzBcjTW4YVcm10WSYdPve6JvlFi3ifq
I2OZY/mHqlhEzhx2IMhqv755gtqRrnnPIfY4d06Ga0UdD2YhgRYCykdbnz+2v8i0kdoBj9iEUZIm
8MsQtKZsfxD/aReb5bcYNMvOJfSOxVdVjI5BuEcYOb6tt3EPXnj+KmV2utnOYBbzEZThdWbCTNHm
Gos/5vd6iOnwghP+5E1j/imliCIbihceKtihmBIr2dA7IgwS1o1W/Eu4Hf70b2QQd3EaUXVRfg8X
IvGFsKrx7WiX2zIxlM6tb7UU0jdu9oVTOo9OqtopPxsrLzTyyM6yMcc/Ftk643/B1Jx4St8lbFCH
UkJKW1/QXwIx6qfIY6NK7OR0JfYtMckbWlp2+Fxv8nEIheaawXEU22tJJTvSSlQkv98kI5x1BfNq
ty4ZatU/kIQWhJGna6kFJ48mFp/sHlAR3zd9yJ7CKEqYj1PIrzx0vfjqUV49zuZ4oDCYcmbI+qBX
VChbxlqziw5uvy9RLzKBK+j1wg2hyJv82TRUZCv2ZhCMfWv2gpzjUmKkR/55NxfiQ/xBqhjqdNWO
VXIWREnEf78asn67CwOUGf+Rv/fhu29p+t1YiSdR+vB3EvxlPc06QDpzvb66nhIhFL/5q6tx1sJd
OOlW+F4CxfDLwwxdYZ/JkZdhQl6Y/Vfo9Jp4YDu4QgpzVgCZHNuc80hi42xneLvhi5PJFWxUyRZF
xjGstUOTiLxFecEyYyI9XMokWK4hQyiL5qVysgYl5c2oYN/tAOSm2xrbBOdv65RzBXYA/zZa+kzl
bQcHiizBIRz4nwTrjMjfpSnGJsvzNfmZRNVcSF3pjd9GH5u9G/Entvu+1IIVAVeVOZCxmCgWcVpa
4IGk77Tu2/IZ0um+fsVdaUlXJrYvVQ8YgZIgYO2RHPJLD7UBIX5dXK7d5wso2tJsMd4rgdvyON3x
4w1SyUbKkUM28aJwylXRlKxasDHcPyjvqP4NnnK0i0dENnHH3AHW+okEYBnKfOOQju7mIZFrqBhK
Ho0XZAHnILOAtz0OjX9QqDVm58to2tOguhOHrKaQWsF3rowNw3Pb4QYlI4li/ix+xu/NA3FIxW3n
VmnTvlUCcLPTtmDpRcLCpcjSZWJiuUyQ+S25GpJaDempyTiIrMuur4SwhLXqMz56slaJvvwl0dOT
rzbDYVqdYvBxtp7csP11X8ACCgHGE+CoYNz4Gw297zJlWtMh/9ODBjmxHXr4Oyeeg2gAM1a7YVC2
7riVifa/Q8ZtPAj6gSvvmg/coHSIwPQABpAtVca2dRHIeSb9MCf5ITLr78R2V6KihWAziKIZ9b54
m60WmHvdt0GRb8Dydb68mXSHcv/SkE1GbweWgTks31CQx6QvzrtTcG9EkAelcYgHZFD/FzMRN01x
9V/YYVS+Zg98sLI1/F9KqyrSyRB9ra+UXPKudJUe0X2wAWjubYbVbJE0XDSrDfp1TqggTmekOO15
BTAvOk5aIMvtsDDNeND0cm58qcGOZsDRC6BJrhK9yDfPAphW5VOqeYq68CerYq+11BLC4n7RcSLh
V9tPx8DyxbIC/ne7neM+ZOkkFdCNTbJVNzxsig3qjaJvpHRnB0mbKNF6G+XZhlWJnZ9UFoB8LgsP
Q8xx8+D82OPIpTs89PJiQadSRvBdqW8y/J7jGNjncDGQ5kpawtaFCHFan3bD55iBLPIXzoL+Bz2B
gNkEMu/+3Sk+B9np7gnEmyJY/o978G9vZ8zuyESzhMOAWPYCbg+CR/A6HT1oddo8lXka8lpME0MH
xvlPz8L4pm9X0Z09x0/O3CKWXh4N6cPQOPHapGlwXuzAA5Prov6YfrziO4ATMzwxQNtk8/Wpg9Cu
qElG1gOnYGXFM3hXlwfv6WUJuujhkMml3QtrdddzRGaqoWUx5SNC31RaUMeU3BD7kBPtwCicPcrq
TfL2VWF1oQs1+5bxK7njRmtyA+nz+/QBZx5XdegtFHOBmbD2xQfmsw7yaKPqRYUkCLNQ+up2zSAn
mRl1a7huvWC2eHg9IlBwWUy5C8IILpIHcI9Nm1BU8cHRrV1oT+GOQ9T5IglF06Zih3kbMb/LqsXr
805Urc6hUYvmcVaRzlXD/LnsMiaXNkhmq55WIWPAT+fWplISBylVBDFu170wMaePOKXgzCySb8FO
EUjdLlgu0X5iYOF0GyNwUvc7lM5J1P6qM/pwL2jmIB7MOlh5qApvV8isag8ygdOYZdqzD3Eb81lk
ajcBek8ThNnApzU4FY85cl1oYOKa+MJCM5reNaQH6JS+h59b9eckUF52/ZUZ285lh3Ne4jGahawc
0oFUi1zPRBiAazsUmE3DQz2B/9Rba0KgumGMyIJetfOQWw6hF9dppKtLFWnlZWvxV68temWsG0PI
qlHYScnBRO6wqgzmBqdjSNLXAPKp/QG+zfSG440Ljkn46ewyiwMHT+usuHRjQBt+7C7u0QfUDrnn
ElNY2Tex2yrSLM8geC8rtUVeyXe1cGcEPbwyonwj2sjbyDkOMsMJOXppMFGK856evTImiWJCPiUH
nGQNuqxx3j7cjr47Z4mJgRNisZTsOontRsNaxkmgmM2seKNfTVXncrGbwJr1N5qZg2fGdjm/9F43
wDT740XsvCjgOeCBTqv0y7XzF2r5XFo/+RSjddg+rZ+K2KNgQRglUiYgTAvHnHQQaVmUzMWVkKTJ
FE/ZRTow1XU1UQH6GQ7BVjpHCpPdr5qx7HhYJEnT3cx42WCTkRFDylduN1fU/FYMrpT6E6dGxZEM
dM5ckHLFtm1p0oxYKsHAbpDsmKDLeE4BdR8lDsqH5QfM7RLRsaoZOK/hXjho4deZcxP4f8YSFJiY
sSAwZf9ZvGllafrendssWB/+tputmTafa0XKpxvxu/120hnp024HRTRFdV647LYBI1lBQX21ckjI
qdycc1Yxa5afa5f4XT71/wEmdCiXJpi2FvLeLf3THTtGFQcn+XGtxKB+Q3rlYOUrR1EM2MLYlr9N
RLyeXaGeKgJ0T4SoAL/HtF6S62GMfrqJpn7vZz7pHQ2j7fmh4SJAoqGmaVrEHpU7RLcDU5j8P2qh
xrHtFpkT/AfFq0ZgJeaJTcUaqx91HOpPRGxDtZRiRKjgKiWIJNxGcGTmFaqnbvdd628tIFD4Zu3h
qOfIlqkUgXDqb01+LLxAgruQE/wZRqEHJxrVoQV+u9ornXHLLNFSndqfl/m+YQoKPs0J5mTcvCkX
HTpCz0ZVHPhyq7tMXRw8dOHBcp8VtPYMrZ9/OD13p5srfIOFCGfpkdu6ndzlJKASKnNPG7Rxu7wm
tMfRsGvKAcNrROTj7w4zwiWhl5nF1HZKsVGizKZ3FuVkRwOI+TlrdTU8Es7M/vlt+uYnxivXAh9S
u9csr6E9i4pM1ObHMfDskyRClf6o/+F1R/mZjQJKiRkeVHF6YKkuDAZYxn62O6IPSK46mx8wrEDG
42G2dCWPn0tqoiclgTjXz35i7XaMH1Udtt4qY1UB4sg0qB9xudEZa9mJkA66RCal+4zTEl8xDC2g
JVf06MvrKYahHgYD7L8lbHU+Ntvhvpd8iQB8lotL+dYPtTpYefgUJfYnqHifhWQZkWYKx/BcohlU
dDYmKiS6TajJ2/dsM4t9jjzBn0p593bUp0HIBbu/8uw0satL0IePi4cToMBHNCO7g7Wf2htkTSPS
+JdNWAnYCKGbV7BkXEsuboK3VLcUrb6OmIbYi3nv4XiP0vo02bvCL2JMxkrQCjivqiiS7FeKf5Th
HSqU4RqrYaIOnAq0IkkRd2yT/1yig7JADI+gQEcJbKZwrpmj2WBrSqWGokuoHl1WLKW1JvEEiw0i
fBsB07l/RKMmgbDQkSw511RvY77KXd4cdKJxEZz/tJZvrxlTLfJ9ERb892Ww6OhfGtCqgJsPpSih
U9ew5QR1Ji8181EYF1V4qu9tNyLdcg0AYlW133QWx5cztNE4K8eoBzyY9LROE2drvP7FxLOXEFFL
QGdnBk3ju/YVXC55tE+iPMqgR4rhCS8UbbVyN7otkaY2DrNZRrKhiDecNM+10faiXpO1Fd42+tjX
W5rXLlW/Mt2/otoFbl03H4BiX8RCnPlWUJqRw+iIsgkKxVMgG+MYphhX6LLGNJm9MTyc2Rk83XOe
m1a5UKfYaH1bpypOfsfnQVa1rEyg7yD8Yc1lab5EZS97+8WBUlGBt2GeC3heD7L+p4fhi6TqXkHu
nNre3eCWbjahvvN6f/FaR2Tb/MDWMKbCuOZQAO+lV/+Q2kXLA5PCotzGFFHb/TW0sf4WxsLfI5Is
oADVnaBLazKwxgkbo5dkYo+LAQjT26yDaxLvc6C9aH5fTIHy48UWmayrGOJt1I/7nBcofVYjyB70
xcQp2VME97s+FUsO2j6PUiky3vJcQtJrrKpgwsziAneJMe7iYFiUlJhLiIrXbNB14yi25cXiH0o/
xasdPvfT4QO9kTgvg9FYoJknNtGJUgyiW30FmyRnkJ/Qgsa6KgChfUFYsxSL0Mp8DGA2XvcnfghE
t4pnWihemvJN88PhcHISfhfBFX4qcTxsmKxy40UUwC7+4ueVcI9qWbsLdtqBqPv1/iYagZ0wo55y
BZeLVpocMTsJWCkXDvMVvDWq2rDNumOqD3EdMfHa9Kv75rZukqMm/+FYBPX66eUFuZLymOiK5iwv
EKaAxIxZXcQTRtoh+ZZfkTcECV2MrNn9oz6ZIVfBFboATIW/Edp/XDdIFR2H8+OIAH5ejSdeNEY7
SQ4R7BwXxidu/TjZBfNeuxReDLoTLoWkvx7PGtrYt6jSVgY6drboVl5jloS5SZyKOt+4dA0BwQ3w
mW8SovgMs7Yo1TPuTmL6KmALmGXvUyNHtl8t4r8O7kdmsEeQv23+YUNjFhKjtDENPFRDzIbltdZS
vtqkf4/ATLYEptW5PaG4xiz7qfa82wRjUzRzUcu4aqZ/rqCetQGgFQqLduv/Urtb8rC3Qg+MAB+k
uCQRll2EUiSwU0z0g9MhItwV/55m3lNFmMfPGKrlpXaQoiVL6B3r/+UWRDUhdrh1wYKA7JqvL+dB
kfCFr7vAjc+FvifHpBF838QNc+tVAkvAF8rtSn+o2rm/u4Puq474oui9ysdSsnu/Nq/Jj7Ai9a1z
MM4yKK2AvP83GIdK1e6fo/m64PdcVb1Bk4L+X4IhizcVQlgDqQ92HsPwJViry/D6ClXiH/je9bTm
05FYGLAsFbaPTOG7j6ODC8jpUiDEniTn34jEM/bSmg1I9kNgZ39YE9U85JDi9jn0BsnIYVwC4NtN
Wpey6KiCtcT++87nsap9YVAnEiSsurtNPxsT4BWqJAmn1wftdW2c9bJqm+Y6tbmQI9LrzodZPjPM
lOTGnclepDI5USZzQwNvWa3dy14RAUeSlbUo7kqxawxuqQO/FBAyxy7LoGIGEySsSA5G3G5jGEJ4
TiajgIo+6o+3bWVlEeH21abQi4tcW9a77BnrcOANf5mxwd9qye3Tr6JQFpujAk/7TYnoMwEJ7wFo
KUPPcpWJwBwzpSTpVS5qE1G8BcBdwphV4i5azuAY8F0crMUmZr6stDnCf5JgaXl2prfGvrEr5Aq7
pV3ILMSU+weVlJpjpJ4u6aFNVI8m1M9aPYgZwZryZ8HAyeVKzh12yksgVVsto8H3xBUh56g+fWQV
ygGNlw+zrUklk5Qiyr+Z1ZccAbMqt+sU2YbLs6E6Dcii3kqHXff0aKxUaqY5apC3HvaVhzZux1Z8
3NI3iOzywxu3aF0KhN5CKcVzTqDiygf74k6CQZUQp1avQIiRW2GoY+3L2GPZKLWN8rlhAFx/WtcF
k6e871JJjmToAsx1CW0sHT6kicSvkqVgX9was7cD8s8PwPnRwpRuIHVuoI7j7uenQvxApDduskGf
M08V8RghVpb7dSdYueUQmjd5fY41cWKFXnZA1K5dsCMw+wf4EqcgeCN4o701jDChz7XMzneB6oN+
lLp3xYGXnyJfis7+dE2j3RPBYGfXldADhHaG9mYHNdOw+rLIiZWfdBcudTMjQTE772KbISPfggxa
KmB463FfdmiLUmGG6VCP2Teih3OZkC3DGu2BOw4c5hmt1FFmyTu2tg2bFGCMR5rBNaImz0XzP9QH
zTSglCm0l5jFh2CZh9YezbqAlKEOVjl3JAvVZp6hK1XatExSEqEykv/49ukZh5pDIwJPO1kz1g05
f6y48cNsqWXa8CfLSlGoCdu8jv6+nSI5z3HKk7bq5MJEND3aelpEybTerHiY3V/zOBqCtEWaef/v
K01/KAskot7uddeKyUAj46dFsIZN7iahpgeDBnTR1lAbTV6Et67YMI17so2CVPM1yGGProuconxJ
fRhcinBGklrmrJNtyo+wzpUJGXyx1z6pvZxeglAgXo0ZmTeb0hc1DGFu/phfPpMNsE1TSLilw7am
980PWeJaje+8IxbsX2QnShUGSbPxtW9rreuwPGNzzMcKE5NRMvgbfwnGI0Vu0j8Z5W80X4qqyzb+
r2gwwOC1pVH3HXx6fkVx7+Kwl6v3m6JP1n3l3o+TaXeHtUlvwpdCW8qOZT6o9bY3eRmfzk5NE/f5
GlE9yG+94sVq+8+JYLnMGkJfV9ZM3vO5ggBU6ggV2h/7+O2CRO9JnnKwirKgo2BnSgKW9z+10Wjf
CZz4JA1DJGO0kCA2292zpqlRUzcCY+sF6C93L3xd1TTsVWPhV0GEcMI5TfDkGmakovG7vISG4GtM
vMxExdg6IITcq128fkaBNBwnbzMZA4tPzIlwMWsHzl/CcnguEV2cs1aZPwm9cpJBlIBGI/nxXq8p
PpVZr4+pX8GkNHvupMyih3IdD13vF3khjf5ae/FP/9+YNJ6y1Zy8UFuOgvKRSrJGBKcvZgW57SoH
QmVJw+ZGejXOFpFcdqEtDRXDHxoQwd6I/i1P7kw2LWLhfgJ8RycHq1Osez0HsFwN3e/7ruXq8781
W5qjnBsYUwkV+xCZFfxCMgHpfRSTCgQh8trJnJHrh+lEz2UuA1SbsdLJ3jPpaPjbGjG8/oGF8y0X
3UM4ApKeFCLFRhqVVLLrJ4E9pskl0l4jj1mIoDaKbKlYiOYsx/M4NwodRmDezb7gKs9v/7Lr4hsZ
JKayv+pfNuLM3jMTfLY/7+0FX8vj99qmCFVLRTLjilMJ40jZl9LasEqzzBCg4UdQRQmBAiJ5aKhc
smIMKK72Hc8NRHhUeJbXChhmo0XuKt3700FX6uxMtfMyCIOdYkfMBBbyrsFJJjNG8PjcJSP3jcZv
BnHjKH5t6LO07drERBTdOEJHzaz4fMDAbfkqqJxoXTgBPkWDrw8JiKHXm+B4qTp/52NSDx1zt6Ag
BiJWwJgB9fDE9jVc8Hl+w5NrUmxLQqLAIeH1WIhBdnCFxiTHzKQ55HH4s4/vnB0JKgxL+UUc8VEb
5tgNAd1Ptg8KtmSZkQ==
`protect end_protected

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OBkwz/2CmGAMb8FOrdhNo0G5iwoR9khBLcDpQfws32v2qMQbN4SZdQbSMwcm2q/C+9Sv2uwuRPSy
RUv9l0tlcg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wUktTDaxRz+gY25F5JayMC9+JtH6VwIC/yvvIcfrLO76EQ19a3MUZjTGOLhL+v2DwypC0R74b/sK
he7PDk1moxbsJgXYeC9GFD/EeaS/4XtqLsnlidpfHnqL+tIp4Q/X4qDiweCY09ivzQ1gdIVg+Tfa
LEdw7WOQHVR+CPDpbnI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aTW3TXFemqcKFqov5TV/vaBSAkJwjfTKZkkxEt9ll4EejxgbIRPSs9Fbd4BD9PjK1VaL1oyd2g0n
4NowocS3Z3d/43d+z7cw9ADKNI3z0hry3pMDSLsO+hs4afRotJ2VA6UgOJDjeb948BcWu4GPhvo9
b3wnibJxFgANvqkm4I/rzMWh/sU7yVn/IqdSDSKZ5ZNBgbXoNjImLoRN/7mLZKMhRCkPKLnJVJGU
EmIWDSEpPqrwXvDoGXFfs2vTTYY5qGAG5qL3Qp13xwcGIawF3XU2L11ZKQ0cuix2R3hq7NhSSDV9
4ZhuCW341rILQwyVL5OUHUQdeqxTbkzCisofMQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mJMZzB69IbSHZ8mSi4XLgtVEk+xk29EZmnxjmAcraR6c+GmgeDlIPJK9b8LuFlbr3QM0Rna4eupK
+ImuhrQZEoDkhh35twt/CrlYjdbOxBb1Q3FFxLNNlqUOlbOlOn1CpUH/nT0RNTz5+Nau9KNK6YnF
/oVCyndnESWBauPql7K3bFuQBo1+lgjc8mLp2IP7WWbTwMC6CF+Pggejm74uh58xKfqCQdZhbfEv
agGgt0D+ktUtWcPvyst4MPgAPUVq7QiAMFcwFVWF0oQfuFAcyQ8vNV3b14wiWfn9qldZ3Q2xeoSC
T0WDwCmB3WtQf4RLCZ7/FfeiffrAJML7c/y7hQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PmJNQjWSUoreiIh/3oafiJAT/DhKbJfdgfBAYO6sctS1YIUztgnXnmw4AX/4Evk5pfDPGz/CPkQa
OBqRaLqabq4Nw42gCVARcTwpV5Wpm5uPUPPWcuvMhavVOxQ0f0aNm408+Si/dWZm/5po6pUyHZBH
Faa4t1wRzdeUfSRUHtfOZqI7QL+g4mBL9Gwj/6jNKLfkb7uNslIj5SGjWslGq34xr9HAu8PymK0J
zuV0Zl+T6CLHJGg/YWuIhqb6THgksnTJrHQ1qKxczGtqtBQDkp4rw/XXMso5vywc6UbrP3kNhFdO
JG6tTSYOHBua4Ef7/zW5m1TjVAI/J6YjLXbIhg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LpdU9xd0LWFvNRJKPgsbOGSGvlv74xMrEkvyUDsaYMAassaGjaCdykNlhI24kihNGW2GHmgHNxDW
QnTGXjxNaCfrmwZSlBNBfrWkqC0gY8H/sXPRdqpuTvkElGoM1q0FUh9fhtOfr4S2DYPRVmC6BkPf
ALqAw3HKH0hi++bXO9U=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kdvreOD3VuHCLspQcu/ofgv5FPL4OFaXLRfNC22e2xDVuDg6t/AA1UtA8o9+javKE+gwAxBnCiGR
RXhsmZDpWOjmSSGFVNE5il1EmINl3QbFCf2um+9w6MUatJVQDUUEfrSeC7841MyEKFc1pF3D/wCT
le/6n1wDtU1BBchHn13u9IRkiCCGwuHk7vgoE0yK03RolCxoWb/Mwv0Cobn0JMTyq2L9N5z7n3Jj
T1/IYvpC39r/tH/vpwM1JmbctpGRY8gm/qGgbeIYpiVLbPDd/8O6F2Mf5zTHqOMNlqNxsjfqk9PI
Ujjjhb0RnO3alxzrF497EvKoKFoIX/7mkxEXIQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
9I1pFIA2+ocxw2qHcbK7WK1pBGGERmkLtBWWyzpz3Cu4Ez0lWHRV+jb9DQPCIgMs9olyatsC4iFD
3CTlRkGyTirITooYWZcTpaQcfqsqIwu22upMrIXObhtSRuk68+6NYCdznFaSP+onjRlS0X0ATRVA
IWU/FPttkBNUJchkRFPMU9MpmeH7fqxWBl/MBMbvSzHXd2xRcMASGUgri00W9q+E7QjDfZWqtYW+
QC/okJHf7Zdjcq96lYXxMrx+CF3TTzykosrMILKpVCTjlq5LCYdfF2/ZBpBFiL+741fQCxFEJs/i
f2eCvXx0CIvpLLdE3wdi57maBSKprxoTsKth2dnlauzJV8jxEcEQ6L7jvePRtM2v2Hmr4Qca4Vi9
ofTZTe6gOY5X01INZFdllgBPHD0KRjua8Xg00rVqJVxkmQgYGsuEXsdC3pZex8j4xj/lPBgRKI/Q
cP1jbxioXiFAeKCRlIrufQzXuyYDHDVPYBSxq0mQQr61K6IaB6AmJPanbTZpkG4AwbIvO+mC49E2
JX3RmvJR3pXAZ8vzXdCOLo0SX5h0Esks8HjJa8SBRd5M/6V60J+w6t/KvM4UKx6vfhNjtooagT82
hahM+pv+o20BX/vlr75iQ7IO39d3l6ykgHfDQtwVV7eQGOpV1l/UsdA9r/oYn8qtfNXguB2o97mu
ZK8NQjzt1UwVgZCInvw/BsfQlDF7hqcfaJ5926veOz0OmhvBwNP4fMFWL+owtnex6O3f6bmslMs9
4legjjZI8Kn0ccFHBaB/ot1Y+WhYf9ycAA460rtH10xEnfEC3VE6Vw36fK5yP5NxLt7wTV0Z41nt
7PxZcL4ttyZjTQyo1IsOZJ1+q1LDHcF/7dzmOryC8AjS5iEY+PsGesfprdFkgOxY6nh4Rw9ki7M6
6ILihlilXV+rXJ9CzvRQLuu/Z/tURTOkg6e0/8h5zf9npZHttbERRnP0M5tGWXWyRwID5iG/M3te
WPwxqy3CrNWwS7Ygf92SIQvnUm2lFQmXwBLfCmDy8nASOi0Fq44V+d/j18j57UufvSi0n0Nsahp2
ZJQ3HWzMEgkL0vdcehOFhSG0QJFZ2zIrbWdXeTq/JfBKJqQTC/Ngbh1aUvJ96Mju/m49Rul8MuE/
UhFA9prHxNQmW/uwDub6+ep1lQ1BTLhwre4700ftSZA+yPpU6TB1qNU8HOftlv+x8jX2KDvtWbn6
TJo+h4hZcf4IFbtK2PcUDKA+GiiAPUYV37eOzt03+jE8TI+f7R0vdnaJba7Ih3Q7I2wMHkxPoBbT
Va6dgYUiGAa7H3xSzi4LccF+aW0LdrzBDpBU8vHBQL8RxmWaYJRUlGKj+4JFKPQC2x6w6ytr8cvI
ktfAcAScDMIDhOySTj/2UKjn2D1+jdROoDpZeaEUxt0mpGcNWKgPohp6C73zpqV54OhBVhbiTsJe
mxGSH9JQTJ1O7zzp/P6EP/YVxqVp3vMpoPLVMsvXu3YMpM4vY2WF67YZDFczKjeN4+LRtbtKEJum
8PgQZrlLRayy+MmTSA6GjBp/uLGuOQCi5qyyPK5jRLWOy2e58JtvWuYAy/oJVbnfL/O1VcfBuAkB
tI+UfaY2F53aMn9PMiMI8qeGqjafTn0EAkL1nJO7QtInEx9/98psmsliDdIjf1CWTAlFoq6TOiG0
/au4T49rw78ycNcgzOZmn1EM9UK6neCPy7y0RpxiIVXYi7TQio1QxUwQu3PsOl7C6k3JoLlbz7ea
DAJIrGp25egxz7SNUj3SpOrpPj4ApLfj8SrSQFeLAMjoFcmBXyEgalWetOudEASILb4rkN7jrsCQ
tYV8u52m+2bO2Frx53tWU155A+syzV8CfiaWg5omhmYgEZe6xA0S5qS4orUZZUgl2IAgkEVNc/An
tsqhEndT/QOm8kzGwM5dV9sDjSZKlhCpxahuyYe45yrvlTlF0DsC4oP294Lw7OqIN5UvwIDL+DeO
EkD31sfR25eG/IEgV7cn5WRLk0t4VS2sdU4Tpc7KjqKemwJHBzuEuSGgeqKkqyNgkfmhclICYowM
mAGfIPVsbpni5o7nIbIq08k+xmEI0co3OR8UYgvjSnR2c1ce4+55pzng3R16cc6TvY04JYd9wWay
DyRhw57hkEu6rfB34RaksC2fUpmh//U1eOnztM2ViTm6enOMweoHPzTLnCXyAhbcJMuLeQicqFjC
+h/j4MSqnM7MSoxLyyzYllrN4iiVyhWImMGBOenvFGqQF9dcj6ZlvcpMFp9pbVGpWzvc9e9rh9Sk
9nm2Gx/383c32MxxvXtEFj7HPSVWp3SiSkqKPR+y7LeQpPeUaK0D9FX/iDEeasl/3JRouWZCk+dm
cEoQVJmhnuCxyC9NjIuIFcbwu5r9aJzgW6vdF9shgaytG+MTwLxXhISS75hiWMJGzS5REOhGc1iL
w0fOFsP3sqW1dXDJIKiuSoSRjgqtKH6JJwhaK5cyKcz5YvqxnYV+SEqVDyJJxxFafw8PNtUKF4y9
yVEittcZnCD89bE/8kfph8PGG1WerIfIoey4kKDh3tPA4a7p2hPEgBvFdlEEovHCH83JlHTLyCwm
Im8v1KnZt/Q8wOjWugjJLXjQa60FX0+NDmHnZcMx0b4XXLs+TdONftg/Z9SmUo3TG5zYRj9LjdPb
paXrY2XbKgiDVkMLOgaXdhtB9mddjOjMXYMxb3gTWdoRYmSWAiJlMK+pV30nZ78pvKlTxgA22+bG
HkHVQeh7MdO0gerRGVG68UFjqSkFWa8ot3aCLrl7DYdf26buGJCdSEgzYhIOk9+2qoArgINw3jNY
2v6laTPgfgCLvAi8wrbIvkkrljdZicz084lqf8se3UnTJsnAzzGpYJjzVgpn15yBNaPKh3FVH6g2
KA6ifiGsGqiH2g91qvRgrpIE/EnHP6fjaftozyn+thkHkDPbHOddb/SgGkkmbHv2MY6zilUVAbTh
YQo85hVmJbWM+xjFT7VYrgZoJR/GDBF+yDg/AO/14+4BLqecSiY3hb/hW3SgFqqELTCbVf/Hy5dv
qXlYdogdQYoxC+LWAYhx3kuRe2CO7omnUkTJ8K3pg5Nf9IxvUP98FDGaUxKbAlzXNY3xhzKjpFxg
5ZuBNddWmaCj9X0KsQ8dnaldjkaNPyoUrwZsdoh4ON53HTDmyJqKAbCMjelVmO+QLsZW3RYCAwHB
UD7xMyz/du5WqnnUzcwlSIqcAhbGkyOfUeH6hwGBe3Ds8tCUrdia28dWIRqIM4MySk3qdf4aXcOd
kp8VUatxepG9/kE/12pGDdFa1KdJ6Kv4AgjY9eMz9oJZfyMeoJa6u7geV6WykGHbLniMH7ZE+jc4
kmXJry0sGpK/kjnR2pQ0KWxDCb788DrVfp69RNlTWE0ViXagtI/lggsuDFwyi2CJTCBRz1Rm8BM1
sFtB3JJhkeatNDALB29g9hiN/8Vh8FYJAXa45nwXhQAqWuYKiFLGIrf6DLugwHMErPH0eYCCiq/c
EuexVHo/A7WQEM7xFfkkpyvPv7LfyVSq2RbBXjkClN+1gHaFXN2vT7Rs0BwyE1pVXksChQTIYwWS
ZsmkS/gxXgokZvSpInLykj4/08QYWJPqJzOgpuCQIdv+bxYjQNPV7oLMh2pz+VyaaQw/hl1cmTGK
tB9GDcaUbhwa/PBh//mKx1SxA0fp6Z2Mw4ox1zxsvwfb7hT47D2jjzDffJkMTNw8kgVuHkslBPQs
JryzbxK/lV0ThthsG7XzIcgpcKV8mxaeAAvoK6iECkzwvPXmIIiJMCTm7JFs4wewvixmNrY4FoBa
Zk1HXFyfggqxtK9w1wiKRX4sJmWFmHJe6Vf91k3obyJae5zd/AcyLqGKCy70eF/nbzgeeb3nVOmD
E4yNAIU76KXaEiPKtlhUsDhPCnSllaWKBx3Tbcqpwfgj7dye+WQR/gWJFAk1orQLwijPx/Bz8fGb
YKiaf9OZMMiz33CsLJOC7K4kE5dmvDQprV8AsrIC3JcFneuWMvDVPvQn72NPqrHfgf5eRApBiX6R
ahNywF2u7CJbALmaS933dj+M1FcsAgqM4tqtp7cQe1hmM+q5rTHUz+Nm2MQG+VZglvKli7MRQaIf
4Z43dq9xwMwAYD8JISM1RiBXeGP9Nwg7UdD8gEZao5z7q7Wx5S4W6CcaQlFFh3C8eUxGsV4TJySN
vbeY47BkcVaspo6Zbke+sbMiIlRcMCrzbs24i+PHVt2RJdJRaiUcdpb0Iu5D+/pJUCOR/fEcf2dI
u9/oWSDjArgksCgHJvEVbb+QX0NFQn2wmFw2cTkn2zbdhusw6AzBZDyMkfs4496Fgy8S/MLe44Fi
ppxPCOoWFmT3nUFb0qqZYP+CLNOIy0AkUJdtUpth0U0dBxqNEEtKrXk6MEUJNCk9w0onhwez7wlF
klgaqxqecdb70Fvte6Q7eeIKtppRM1JXU8BjM5BXimfycH4V6gQz2zm3q8KiwNNyL27A+791klRX
ZZOC1jjUrcInNjRuwBELuHyr4h58a47YpkTzFDlNI0TUud1F9xa5aqG1LHz55e/Q9so5bDvZ40Ab
Ni3ZH0Q1iSfZJ3rgoXDSerdFecMqDcBsuew+Cl5PPpYcLjZ5aBBTmam60jCGbvfcx7zjyQ2z45gV
G5h7oGZHiWuYYvvPo3yRzNoxHihY+yH7b96/rjlzzfaHocwwt/+iPWnOkst/mHIF5msFlNalDRkL
BFkGIWWiuFC1q/NhtfYsR7RrvulsaFa4UfT9lafwGH2c9P5vHq2u1oqC+z50COhgniguKT8Hkptc
bYRAkTXLG7Qb2NbdeQ7YcSpRYHiM25NK6grhg7WJWL/7Jhq/EJH8YDMjMwlc/7c81F5wgU1XZmaw
sQAM9CADy6+HS3ANtu77KPaYAnsnyCxYkQ6EolzngSzjaadNrDsYpqp/J0i9CTn5PpMomWhIJW3N
5qr819hG0onL10jcmP/pkkzl5vw7OWGQCbTdG1r4/y/ZS97sFuOwFhWXfdjNyE4Em9MKxr7a2IFE
sTErHoHQLxq6Qn+SMGSukWppZg/mq10uJN1txUKqSJSUA8O5Fn9vd33SVWcDPZSOr92p84ff2y62
OqyuX01BJ1dtoGWRAwr/NrpEqOQJrVyjld/OvRxq274SDD2QZpbN34h+lH+ALYK31E7AuN6kk67N
2tnPkasBvXXlVwnruq0vPpYx1qGU6901QIpOeRe9II8dWVTrAvWyDKd/A+FnhbYpeUPgBh02xikd
yJFPKTrG8Jh+AdfxKyOBmAV6EhRVRWz4ZvX3cQzW1z0gu7n4t5Z+dvv+FpVK9alERgiIjpvgGYjk
0bqOV1ru7o43Wv7SELcbek31v9VNRdUspBP0BsN35XfhIEev3ShwMTdcDrdeCXqAFJlg15QaOUI7
MaiuSEi4EuZVyklGur2n7Ybe8dLMsntRNr/jvXGvmEEj9vB3fgiDjOd1umYA3Bkm3mX8yqPQD5Kr
ajdnxthMSuSC96e7//LWOOo295vtYmz0Dax3KzG5MwYuySXvlPudf8Fo6pcZMUc3wzD4E6XBkP+U
4WNn6+FxIzbZqp40N07ZI2szMkGyLF6rIK1e43cBlVNtUQRY7Fbgkq9OeFt3z35TdIo7yMbDaKm3
fOCGqe3ML0RoD34Ik52Mqj5FpGvWxWz4Cp2UqFva8Ul/rO38JE+cf7nnG7tApci1XzmvSJp9nXh2
/zqDL3WMiKGB4QI29mHT6QyXEqrTUdR9loFAp5yaQRa+oKjcpQ8aJUTo67UWHp5X9Mx4Im4KQwjU
dsMW6+NNtKx1eE1MwV6DrAQm18Z5Coxitn9Fu+86c7SW7zRbzBRPIqtyDP4YATxm+PpEBkmWR2Bw
RZJf9aIt8TDZwjCUwuMVNktUkctQGHGS8zK+N8WYktCaQNcrZkc+CEZxmzhl1MCKkQkuEqEhFaV4
Z3oNoupFofEYFoM3oqOpoUr0zC8abiBfgSeQSmaaaX0ugN2nyYpggnx4jGlx7YRLFQsTZFowdmLM
J9fn+26hfJ29wHr36pNOJ790+3APu7/4VwHVmJ39fYiB9xAS6+esRu3JYYsY82Z+blVaoUk4923u
z2W4lHNDGF2HJKohrGtjr8u/FNp7I/lvjtYS/lj0mPhxe5PbQBn+OroeW0nW2AhC6O6qUdEpRIzY
1jrMnuhrNLq2Uv/AuVJ6NUN3OoAWxMy0Zse1KlVtTo7TnYTPoQGfSg9O6ihQ3CxcOe7OdS7uGjj1
Wm5dVkG2+cuHMdETCaMKj05yG7SUS3SI8nwGRkOpbKXeeXG/gU718G30FN1+HsaQnoLlbepCCQZj
G7VzQgLm5J+cLrOyyst2Q5MniAq/4mDulZdU84Chkex45HpwhhSmbDIK2V0CKz56B0xOmJL2ZHRV
RvGTZKDT8xN2gtImTJJhq0D6av8rsQ+oM7Ka+xflTIjx6VOQf1Nvhkbh2GDWiK3/gQelC9rDU+jv
CtiI8zW5vS/LldWpuvqW/Zaum+j8OsKf9GtXObMB1BiQuUJuKaNbSdbDJuaLtiawXR+CrSqzaDgL
6tSTAL0TcXRGvjn8dkW5jfyMhDIK8v3j4pspDkyyawHDKZgO6gOTLWvaoKBoBje1CYfnZYFHA9E0
Ls4GN3v0g6loKnFRlLd09DGhGVbv9Samd4PDxaMe/gd+JQhHeed4Kfesu7KMJGNJRUQFISlCGvtl
RGTDG2rTI+u5h7aS8jQkQ5DvdBxfM1d4N4tbw09j/rsfgp2tNslkFyMJFGL94SvPqBZHPtmNJKu+
8/MEp0JaC1IP9qM/eMCIJpVa1aMklay5R454d6jfJm10FuK62viJv/RVmIBfqvYWPrxNvJoQT1zr
09QIzCIKTxxU4cI8MEc8LlhKHqqIhiPmoiCSNqd/u1heKQ3BD7RngvVw9tG/0gEobnsUh5dSzK/A
aRQs4rB99O00mAIxZTpmS+Pz8l4tBj3DSwMiCpZW2/jGy1baQW9PohBBzZ6vQ3NhUTu9gbINbbti
rPBnNAbnUSlIlF1UREFIKnxkhIp/11t+uOHiCNA3DOiJOq2+ABO9Etn+VfQ3QXoTmTFnO6isf9xj
Mkyrhk39KjQHEI/cs2btKuIrrXU5q0e7wkJgQ5IzO9VbTOsAtgOkHEJrAQGRm3tHEsvhwGOuIcP6
VrlGlZD5ERBv32iCoIGt1HnOZvlMfmnJZSG9SarSGtF//gxb5zHSfqz/NEinqI37KSOMORsj0lEE
arBbwaJK7mriClFJ0hkHThx7vP4DouNwcgD0H47TL4y6TsLpr6Y8fR8ku8Msuinhb+rS85wnjgt8
BDWr1Ld50UOiC5oBy6koYrv9v2sM2ni2krkli9kEHv6M/IjSZe+G5YUNDdfnh701MlRFjn7U7Cdi
aJCvKpRpd6dlqQGcZHXmzXSH3yGiZhUjTRjEUC5dOZ7uEXPxjXFfJctdT3/TBwRu//MS/32oUDlz
dWr4YmEfBJJVP0u19+i49+4ZbEpr8DmJ8+Kr1EBcHk951vvwoO6J75eWMPdgN5R6M/azBrgo2TPt
eZqBqrriImfdRrwW7K6bv9AFxRv0i5nmZqSulTvQRMUxZmxBs3+vyAo8uXffh2Kdf5JVq+l14SCM
7q+o/RjDOdH0FDB7y/UIo+YhGO0EQmUJZBVq0EEJoOfGx/YHVNZowJ59heOjpS+lnUdk2ryZJ1cs
ruWKsOpkm92KWZ9zAH68GZDDW2D441hDm1Zns1RSeAz6asOg3F+aCZ9Yu2xtA6tDAfrx9lP/Sylx
sEe8V1xzjURUOkKgzppwpPtYTenCkiVUi1qgvn4rh/g0RU/BPuKFOAnQYzI7Dee3P+rWc1XfYuvX
cdOaIbNwqGCoYzshxhcwreeyldXcDxpQ8nixZ870iSn/qs1qcVOtP0F+VGM36gAt3rAaQYTIaKem
yZ2OCHsWehVw4iSfL5bvXp2EzeSUIRZu29Iy3S6ZUn7mdNQtKLKFjmrhoAiZEU13PjQcU4OSFbgg
R52c+2zazCQe5BfFkZakAj1nm1c/CiH2GZriX6jB3/63Dk0eyhF98qYFFD2/JQjTRlaKGltpKOOO
SmtYK3wycHYW61AvQASeFV8zRv/846fOrITdT0u2/gtT1bhK9QssqO/QTaSp0ptQMD4RYKSDh3ND
tVR9bjn5zRqslGoSoXJSn8FL2PTyw3kW5Lqa4dsT95wyNJTbXwFMJITv1Y3KOp+VuvODWz1ttR51
bPG4+MdG34fH6Xh71VORRjYHO/ApjOmP2103qmtjcRSq7Z+CFB89rarXUyEFSODBsVWv/DWlYQ41
InxsSEiXbrrg32qqPqE4VQRR9ZJh/wByo9U11prGqSfedWLGP/kysmo35ZukteXwu7rrHyMJ78pv
MjJfyknDs91E0bpacg5hBjI+Xn/5cgX7zLnTTh8ZrBVHlu+KekILeanzIQGBTexJ9xHjWAAcR+2K
+twtXIjNEKVsOBsYqiT5TvPF/s1wNRr1J4Bj7XIAVqpndDh8wMF9WbNGwiF4LBKc+no1kiWubTjz
lIgh07qHl9Pgxn8sgtb2dyhURk1iuP1BaTUannaFbYTd2GorgkNTjJSE7G/yA3ZLdIqaPPrncuqL
6z0ITCjRK0GpBQpGt5TRAXrFTuo7F4g714O3YSp4AHJNA2SemXgeUCmB75VVZq7Yce4kJhsUiQtQ
62CMKD1TRDt0oi+W7GmHwvEX6Pd1AMOtkurKuZNQ8UOmxN27R4H3YOjlLQh14NfotD6JeOzlKR3P
qUxLCiZL6/L/FGui2KG1G5mDNpiFqtlQrrXMbLGBi46jTf0Ga++Yig5My39IvNHxix4NuyBVoYPI
aTx3KBSqvRLJ5R9iMCDr3GWJMbtj/WAK8iY9ChQraqlIR4cinULbFRlXbWNNPkzc736nKM4vhkCi
Kr+/WQtxlgBw7NB9aPH9nr3rpRCu2uKhQo1R4bcMu92W1+Iw9La1tqLDZsvnw09m8DK3VPgKb/Rr
oWP+gaGpxtO1nXcu6eEBPVB4wzUynSjw6cUWMoDlclcipv82wT9Q1HwWrhnRDKReNXzh/di2utsy
AEu4xVf0r52YsTcYVyI5xvy6f3xdx0tBpt2b30+GmNAe4+Q6AdnrBQM4dR1WapArzzc4xxw7CgEE
D3qdKZ+kbj504J7eL6HMbfpzhvcZxeS9aXYZ2eqjP95HTQbdKrmHsJl0qMhQBmfGFjPwEC3aMzEY
YnTkgwkwL3U9r2+u8/VeNOHf5OofeG4+B9M/zxQITS8osF4cy6Q2+weuUIwBEFSWTpXkXnrWoy+X
roXF5saqBlvcsdqPnKkysYJXfuupPzWartyto0UfeVXNczXqUmoVZR/rFE//v9V3RdVVS17x/5Ll
i+5bad9DRvt2oYdDBT3/RHVCyC/jSe3Eg76Mr6N9Jy+MGkz3L16xiRm1OGZOJYdoPQXHqO/sY+Tc
UDPvMwyyExH8XYYTWHI2CMs4gcTG01B9p0siQPzJvqEoBU2OzUuPco/HlhZEMyM5W/U8ghDflr6C
COdzPXQZ77+LdWij3dcE9aHovADI5bLq3xVv159do5Twn9hdh6QtwGm4UOznYrJT5NtydYeiA9M8
Th/9ZGs7BVQhR1voQFkR9p8yeQuYRxqDesp3Xup3uLUD9+9t71DAnMWlSaHe/pK+xBkI7VUvtsHX
6xg4TIac0t10ZVYVvhv9M8qntP8ACZkVl/SEyvQh5vbdkVtsglJekOpNexjzQFhPL9iZ8OVsLN7n
1RSTnjUPVnULA2z1GBVXWbwlE9g8kC/VFDn1d6bGeDDLY+nDl53TNS15Zx7CMeT14y+IRuAXG9GU
69J7vnpd0LOuwaDpLzS3PQPab+vJzZWr6vJclgK/iIUtP6Y7VIS2hdDkoy4Lv0lAYhwgOqmV/5CQ
Khol2gLJougqHaikroQPCNo1hP7wHuu/k6tj9H8oUbc8wz8d5LGcAxhnpkvwdiLc6JkInfRyIRYF
+d9tUhRl3QBeSVm6f6RmNf5SjOinF3z6aRiEGtO0CtqJSo8GkxzwWhl5uy3W25oUW9PIkwru+W3D
M/TcBfYlyIaH5g1mSb2Gp87Vp7HfbRlSSegjG+xahkUL5L7HoXvaFVvtEBXv4wxuU2FliQEXc5UJ
L3jUqe7hnoik0bskvhuYgp5RPUshVw4TqS/vxZQoU8pM9pQs5StgNiKcoLOF6TFYJwpS27N7LJ5g
ETGJ81cMH4QEKBhx0566BGi/otJLjNWxgDlKDrtEfxBXKeyetBfTWj9a27dd7WLhj7ywq6SBd175
7GhUFln/958OsgY47zvNfMuHbPgKSS5fzVJSXMOcN3he0dfzDsHEvkRcK6xbUYA8AFWhDa0Finx/
/5sDECM933fnAzvDY1yDoew1cM1UFBU9ynFigdFP8QMd7Br6zozlxRWFobSyh0Mh+O7rFW9pL+GJ
MMkNSXcgRiBIlBus73iTbDQp6AoPpHv6/Fz6mBCnjuHkefo1BE7wBQkOtHvJUJbMFltLmnzIQtRL
yxMCFubtYtoqYvOaNl+dBeGTZanj51GUgDQaUvg2MqXDuk2xqmLz9okVfpgod2Tf6As+WrPML5zm
2yopJJAWHZPtOf8jF/G3GtvqC64B1uloT3TR4qJ8TSwTDfIaDA+CAj/h37l5KDC6KdS+itLHCXE4
fivzameSY8CLxQkzl1iaZh9yZj/yab7LTptww9KI56fFmLW5OhhMhNaKZ70d4+I3xuLQvke6WRU9
P6J1NqbUyQHelYrDpir0fvtJWEYGkNPh6goKb06Ui7+mrYkCRJVjzjU7lll7/mQINrs+jHZPoSwU
ApPfg9jRqRNoqB0r61SOMIp7ATqnmFO93IbMcvt/oMFKrC7Iak1eUmNaWzzADrMejHFEdxwoRSID
x0KstEFvsU6ON4TBelX0hg7bX0KPIY7BUzYzYxPSDoeef5+jEXsntMdjTkUq9OSPn8yDJMpIW6tf
3W5t6+4st1s5DoEYfoAq6wRv2isQ2rigbtyu4k3/yjFWyzClwsakGkdK3ro7fjJZXvC/kv2qSB48
Cvc7oCPB3gzHOZdar9ZA9exAnSzVY7PoeEYrm43rIUVNutcTxX40wN9nsCk5Ye2QflP0GTahAAb+
rp+dtTV9rWExNQHca9OMyXZHUotTZCve0DYf41enaH0By/AGZN5t/BmG9zkJCFt4nbxo8hgZOzrp
JyWXLEITeOeuDmHM4RUPGN653oeV+O4klyRZ+X6KiyszGKk93Ylg0m0fo+nV3M6Ace9SoQvCu/We
fhrImGT6I7v7GSI59dVbbDy/sAda1ytSZ5APZqDXXjd9jGZ1LHPHWabQVxT88bX+EQ9a5JwkR0yf
hXRS2LchM38RX0Wf4PPea2cLCwO9WjuCYrKKdXtBipCM1A/cugITQv8lGOTY7zMKHqAVwgPbvmjn
vu48bqsNhuC4NZmxKKsy8Sepmy9wkvyQiKTBHBwbjRdQ4G4fcOawOweIbeju7iCZpN//G6FB0VQX
gts7Xfmi37/9nMTU7cKpXkmxuZsGlqHON72VZ7TnAQfpc8RoonZjgyqv3AK+LVwKwF9GEhkjru2H
aheQKf+Yc1bMKrTHOfa1R8OEs3/luAaWwStymBGxnAc/f7aQgqnKp1wC1tSn+4iTQaBPi0MwYqZ3
SsBCdlFfFngXZfHmMXAxXFjoj2GwCDowI77EaC3wsqaxeO+iLwy8Cm2jKH1Yly3UeC97r4K+oipP
yt8Dj37EAzLcmp231nvm1TnLtxTkfoA1FKWaCIMwjUmwmX0x+6TQ6SiC0SpSTqRZSOaR3dAYjR7g
ycIDVxMgTjS1WW9a0kBZXT/QgiJsM6W97Ul6NbabRio/q55sUAnjkRA9UGcbf+onvEe64qgB7tPb
HxCF+QeRzhplgQYcRPzkJFV/PM99THs9yNVjyHw/M05PX/2C3vx7heZpLlfKhoflmRmlEqOZ0QmG
+DDUz37awlIbBgF8MCu4QBjeXoV5NaWkyaFEC0526P3DHLFGLljrGOsR30rCYtKScguQYlB8Jj0W
mY79S7bBCFFCO3JKbMxhKFjI+1PnaAmS5ZI/kQOJBJJpVDxC5b7FB7kQuLOLe5U5VsIcDs8TMq9f
yFbxtSfwrOVukMrxw7tpY4g+NGk3gdpF+CKHGAA37LDcujp4qIlTL6deth/MdnC4ox7rUuUsA4D8
uJKW0bzHZy6Faho2INHMMqIRfVhFVL0pR/ho9+9pc1YVW27Dz7weHii4A4DnsBG6Xaq40/o4sX7Y
7w0XA8DStfUL0mHTV5MxwAk4SMT+V54UAf1O8QDejsvWg9y73heXDGed/IFA8xuLlqaRfiY0fwRL
vnPUDvKy/eCzzkoqchJQ4sdImxIjPXaiSgbOwuKRuEjgt0FkCHF01Voo4D15CDErdnkad5al3ugS
0D6r3tXjQAkqJi+biUDSROTdJCQH4YoxImo6DRUw/F0O+zJpWPHZfwruyVyr9zSj9MuPuyNqNduO
J8I+jxRHC4/x9xqH7nfGQ+gm8YOHXCeVIF/SRKJFOOEjX/SLeyFgWo6d/Li4X61PNPw7+Dpoahcg
w3X8/Dp3r9IZxW1YaopBgcMrp/Irn5MXRyJUrhGg83IgJLm2SlKGxzyQtAmFrgNfRJ+n0BslWUTa
iYyX7blL6OOyo8iwPzUk3k/MsQ2pfYiYVkkHDHl+DELifbniW9gKnGjY2e4+2rKSGIi9/ntO0+g8
5sSB/7haJPHqmQo0pH7gi7P73Iwx6FBw2E4XGb0TGvi0Vza9vgCuuhOVl/dz4sCLbiOmi1WQQJMQ
GYvMpFRLuI2XlI1OaajNb5SrvT0IoMBHMUSYzSM96JYSQahWzJaxLzi6kJBmG32Wla/RSZNjyzhi
wT0OpFIbJ0xb4nfPlThsHb39txv/8LGQdkDmTp3tAHkeX92NMSIzuazwGcUDa06l6QOmKqBRAVNf
L/M4nhEwQHbEimMvmCffJaXobxOb+TB1afZtkgofVrzUf2bm2quCiJ2hRDXFNcDFWfOsiGT5eO3N
9w0KyOL0UCGMtQMOi+brjQP6bxKFfukKi8X7y+jT/mZ95YYprfhSZRUjNxzzqX637CsfxFYZBsS+
zglEr85VfBoKLzI73urIhJcnFwhi8QzJhrzTaDyoDpu4OrKR2Q3JzVEw+ZBwto2kMZFiDh6dfOE3
g5sapKl2SrsJ2hvDuydVVhOKDkwJ9xVsgGaSQF3cg/YBwaTCQCxU4w44tqjUuOjTvtDLL2kZj+G5
9NnqFGdvMRLXAgT4ofJqmfM4e979eDxESj7iy6fHqy+foDYK6Wi7Rg3AFufavytxrtiMEeBaQPJK
F4DS1m89j/fDu40almk59l1upRxvEieOj9IoCuny6JgNfS9iB7rxra8aSWsKrANKdQKlEz2zXeyZ
yNgTvNuanP2r3mffBEP5/iQdsG2kRrfCYD84xn7l+CpFDWL/Lzw0OeVpBfBh0Qi8gLQcPBszDoE4
MqwpEW55GNcBIhh26zMPk7SklrzAgqUsnaYM+B/s7mAqgwM6cI4XYbBG8k402IqsqVTPx7ANNhOw
uUQCFtIe6dvqqiTOfrPK2xzdZ0TzMqviFV+wZwwH3FO84jDnHVhRmV7Bd5r2mpDd+O5O4Z1M5RwZ
8TqqsLr0gdaDWPejqm7veHLXNDX395hj1a9glfWdlXthbijWftFVwWopgJiJfIA7pVF2HGlNBAmU
4dbu9bqkXVW+AiEwaNYTzqOdD0EUfI9kDC4WPJJ9ugiAdU1etXW7UbuI3rufQy/UuYZTexeiJugU
yb0athZ0FbMZL4cgnKxV7HUilJrSsqqVChDG2/HVfat0j0lrdBexEoCzZdBuasI/UJwBGvYv0LOe
EPYuzXnypR3VgmXPR0C/JVIzpUYAkBMd1fFziFfdZvkFjPWAvTRLJwKnUH9LzJl4xitFUxxL/eE5
dXDncaAYxQp5bYctX7n5fTeYipwW25lDBEZu4Q9JhgSUK6sGhCzPK8tRccAQ1uU/GJqtoMWy8IRI
F3i2TAyl+V4ZEeA4QuQMi6PQOnGoymbWLNwm3v3Uia+1rWRtMngLcrGKSoZoKfvSE85aGeP8dwvI
Zdx8FjVM3XLyaJHAdEgIXEn9wPtUxPsIW1TXKqh5fan51B1QpPbp7i4UZhW0pKKYw8r8LtkQwBBj
MBgWKnvZwqIL03oAs47ItA0ti9M0q+5aEB5bKfrHsYtMUznTv+s=
`protect end_protected

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HbwFuGRaFcvb7MU2M/BhGkMBwIIsNeZ5fSlF8uuxoE0oA3vYw7uv584vEYR70QyKw6fLYyOkgpyc
T5hGxNq7cx8YhXgG/wUAXoui+C04Zm3yiBZ4QxYsJW1QLdFVLAPj87n7KKM5BqS013Kk81soToIn
MGZcD09/HifLLbaxoesqtSiFKJa+eRnh8vJdtMVoZwroeGNXwTqKocXB6FPvrQZkv/cp3VpakTsZ
fnoWFjJwL2auhFGxUevjGYqy+F7d7lyVLQDVDZ9xclVIEvD4FRy0J79MqrDgT92udk2C8c+9TfXm
sb5Ghvd5b5zOYe2BB34dGlwbRYg5DzxTdeH57g==
`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aj+OUQlpvgBZzH9dgL8QoxfrJAJM5oa4iI+ZssT0vHovmzNAJfatfIoYkYq/rHvcZMvoNGTDtaDt
pUDQkd4jVaHuKIM64x5osubWvHyVrOUG9g8NcUoPvxlQDIsXLSmikj3LFCnc3ZTSN0mCeP8xHOBu
aWGIBIqq3dBoqN3PbiPyWl5QZInWodfmTpwRiZxAjHUgxKDasO8iWjvI2n7PFNmIQ1fSW5lprLSt
J9Sz10auG4Wqp6iCk0SOVhjJ8eOZavn+E8ct10cYeCq9WKCmNa79UWJDkK+jHmIoR/nIeIbib5KS
4EgH51vb5m8i/qAXBGIxgS6fRiMDr/s4H7eWWg==
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Z8hi9RXBCkZkXNZyEs1ys8McWIHm27inhdp8m7Q+yGqQJ1shy9UCcdvrvpVNziJI0EQOFVHEF7tt
tOM8Dr5bqA==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q5/Y3jxT2XGT066NAl0eOzhKdEVSVbEJ02J0SFltdzgZJg/U+UVReaODhutxiRSl43W5QLEmdLyW
k0Txzzk8D42DyVCuuKdapbw6fP4yseQtcXxQVhfnu9bI5zu7BlhH1LekIQ2tT+gOrZ+kKrMgzrEL
VvvO/1851UMo8XFY6RQ=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n1iy7xnIhU8AfEq5lLzzxXZyZHJXEwDGUtZVEFfXBJilgwSAgmdRl6zpgqPQALwXQgF8fBa3ZIz4
puTubFskFM4T5qHdOe4MGCcvZjQtqMJHeV2m5+qh1gnhSEx6W08hs0RRuXxncutTIyDhmqd7x2v0
WIIU0jnsoQj+qXxiZqD8Kl34Agj8XSJTKCjqM2y4r583c2O0fDCli+YEUFCS8GASTXfs7RIfD/Q9
jCMQLiOvNjb/YzNlxgiL2GCwY8jl+Z4HF4fXYBsxBUnggiw/Jjq2bvErW5yC6fGKLF/kVBIMVaXc
B8LbUi9fRbFG7K0KPSYU8ovFhk4+fB8Ke8/bSw==
`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A9MCbfXtzHjSVxrQZhrJdVQ24Yf+TxDUqE68yn9m4KHAYjqM6RQXSsQQLpKtsirU01RDLh/A7nOE
PpUEMXMpe4vJQbto4tp1ZMc/0/a+tZWRPc/0usOKkRGvDvxGblvit0j2Oah4O5muh+iyQClJ0w+6
FyxK6mc0+76v2Y9V2zw=
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lhj1qQJEyyFBjgwbpJGaLkSUbV7+DNNC9LZm+proCJVN8Ot9iLOJHwYcJ8kXQbq/I4FO6SURr+O6
7QZI5O5GWaMqxWF6IzYBCbefJhyyrd9x+gsA6hYpIT5lFMyNRXs7kvtDNiaBuwXi4UtVcAREdZsx
oNc5tj2uvyPqHYqVaFqg1t7N3moCuEfRbNHDgAGyqyyY/Va3pVaUPw60djupUdLO9PdC40+ebYXI
vqrZnbMXDbv79jYzCQrdUagiv5/4LaMxtB4RFWswkvVYYNzAuYdewFa1PzeAj4PPwdfD6EVrUoNn
OjKIFg8ztqyR/kZQOObMDBLprW/PKONrKBGrpw==
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59280)
`protect data_block
Jz8EFAXAAb3I0wpY/4LGRW8kcFb+TjDNYrrurPt86YV9A/hzVUGmCnnsmZ3QIojkgdglT9e4ZFmF
Tq693VOi/N7g0/QfJJ1R1qFGZASy+vf7xPUjmU2lDi9LMd3qO7x2AawMhwYt7Sc1loFgXYCPzF98
b/Xu5EqZbDP0xoz59W/C7GmvTeMzEMYcWDDx25tbmPySlLe8BYk/yUgEMyy1F7Uz4dfB4vavgNIj
RA5E/KlgH9J0f4taor2UUqItdVGGMv2SP7pK6y7ZfXlqM8fsEJbwHn1OM4JXsORe4btZAd0U/A07
mDGm2tuCbewB9loByq+kGM/bDfpwTwHY7GnryM0tsmFOXX6BXiQOJvPTLZRV/AfabKNdNubeXo5y
9dSNq5rB2t/mIV1r55ZWYIR+0LyiV6ZpvIp5FSd2ilomwHKQ4eIWcVrQIuN4VEzcBwfjtCH69iQl
RC6kab25qBHgBYMCzWLE35GgPrCZmYshLJfaZNIN5r46oOAf+iX1jc3kZqBDcURR9oW6994NH8Fe
7gE053ebI/j1dklj6ISGdu+IuPQxtgqV6ibILR+7DtQWBjcnIKHKfKQctIwcA1gRUtjkV1Qcm/7M
rIbAbx6m1/z75AKo7KyKsNARjmcYvQfNsejmnR1cT2irWA7QEekinYB89l1GlKkXt1brz4x7osKd
EsK+uTEUIMmqZ4YAFh4jYp7h1E4j3yoNVnIaY4/Lrk4Nprnce6YYs4h6yymYQF3a53U0TQkz/rk1
wteHPdLz29WLNvcJ3RJE1fY/EUxp9yzrKmGoUJHEZunA39xt9P77iu14AP2G6V1t+PzFWzqHIZsv
fxoOi9nN0mjj6E2vS+QVDipSvV59erP+d6iPSN5RGMspCuQ3ynuP+Mm2g4J5mnnzHTT72aN6phlS
4s77mFPzDvJFb2sz0nf0E8k+8ArAev5zL1RSeyTZI90fNPx5wUJT/4iSW/us59/QiWY2z5HPBDGe
zyZ3nVFUVQv3gAGLGiSmoXIAd8kQHhZ2mNN0h/xRAHMSJjrZQaHN5/tU17e82pr0SKBWBsk5f/Pt
CYCJ/n9LFENykimK5kAcBRoAdI2Rkz5W8wrQ3/2esDnqobzK2JhNJoHWT1kArc8YCSh7A4DlVcL0
S39UxxvFZ41weNAasRpCZMoweEkbDgZ7RfNgK0hiNa8gNonc9B6YSkXULI5g8xXmQfPuAh3PrBff
7IKQDOpP6PLcxiqghwKaHWQqy/5YgMZlq7B9hK8vN+QZRL+QthPt+RPVrnUD93+CoHvbqdBbRteH
XbGgOUh+N3bfArPtNbSB6fgj6d0J/SfVfA5rJiV5ztF3cZA5Ft0/3yw176VrIdFiJx0ca8a/VWd1
JJ5FH0YF4FyaAOJ5n0TMLnCdlpPyAsVrAaOJSIEY2Ng8nmonRoJrGDSqlGATPwvCn1CtSwoOfqX+
ZfXo09FOiu4WYCwPsb4x/PeRl+dC+A9uHjmTEkrdTLh5IRDo8nOBZFmfsAbp4qukWbdTDiKqmfGz
ETDNAYjjMjwQQD6sRR0K5EP7t8uwos6Pq1Ybbe0dcea2Vbf/W3KvEFhU/JOm9pIBrhm2OeIybJgf
mqEY4ROhvmTsOGKdQWvnHydg8O96Yv9wLBiw5Y6Lt+WuLczSRyvdtPj6XU/2+hwpdG5plVvxVMGN
EjyWULhLtnWJkbYvzYHqa8GQbdu/GnLf8/6n+Fza4r23KEb9yGbCWxr2KwMayohPLdlStcoHaPeF
PM7X1LjkwUYn2a6wDBDBd4lyndG0cZodIWorbiceYu0CMyRL6xqjVdgIgNwKirN8ndyRtzg2XjrY
vi8ICweTKDJAJGcpi6/u/SE4FjhdRP6sUI27XeDsA6sa7nal5Nf4jUVf2Ib51oxTgU7j/sfxQc2r
qYezdurJcx/4lZXDPZ2tpnQTWO53W14Fm/oceOh74bb7H944aHgg616uGAv5kONycnhmQGXAUpbd
T/nawv3/EGL/wWHwz/tRszek0Op4IsslRfDcH3q453vlQPZI5aDXbANkGZB5hqwnP1bRYyDsTXxy
Sy1pcnM3qTtAJU/CXBEzlwIu3DPwUlUsexk+8Hkmqp+SkFHM14+toSyucUUp8J7B8SODG9YFqayY
Bf3mOb8m3Mr+EnXx6bT60BJFEYb2jRjpNDmxEXYO6lsX3gP5mF4DWKRPxJ1watN4PwFWDR+AzRsh
scqvKa5GPsFWrawVNX3DS9c6b72akJydQNLcr4SmzqtwKQtbe1MDE25r5OqFiBytXgtn6nBCpY2j
cCNVZ9QDxw/oRulGVFDM9NXlxSu7EwCv4fx0SF8JEJYmIiD2fxMJXITMmtD4gUgzFC7TCSZ1hD0c
WCd4TY1AdDSRdSW5lQFQfzdxc/nKPO7mrgxSGOK1ByhYIgreNkeYdfxKHOPqckv/cg3W4ohTT+z5
7c1mZD7bNVBu63kilojSKTOd47o7dQOa9VfoZCRoq2w+DinGruRmAKP7+ZVtcbWWfFf2mnzYaWBB
iP5clIKnLJYEiWpzMtqMzklGBh+wSwJ1h6dAr0X/Xu0JuvllWyXUoVa+PP+CGpEGckJac03ahaTg
ByZpBz+sNmZSCtIxNlhyIeTo/RtX+lrbsPyAVviMZCgw4tVVUWhmnqiNIn/xv+0hsUdJPziu6Wi5
erqsdRhJLbLayaQR45yxoyQ57K/GtBEBZQM7Xt/5+JH811r18xG9muWyrtfc0IBeJVhbvhchfiDV
hHePyX6R8jpeA1Bag6MQDwjFBC7EpDpkm2DkoR2cuQ+jQxlyKc2PDx52+2yC0oUEVUwgTygY8k09
rVUtLxW0keicT9inHPWROPvluUprapGvlk5DAajONjaCIz3OPq2fJSxSCqD3FJfCKC31MXgD/sFU
uoe7+yfboN06+ikRorXntSRSIOqbu6McU+EVvLZsl3tEQJEt6DUtYnxLLNXjOqt0Orbo+TmdoYmM
zZyB4sKvjw0/VBZ0RV7Eu0XY2ykVNv3OcPsY5g7O75HAwQoTReSmXtTL6ZUf8uj42OsUqVDKaTX1
w6h1rrhbXxJBdMH7twwWRQ66qOjkiG53/ZfLf2hHlZpaOUhAVDgajz6tpN8bn3KnPgUPsPR4RoNb
fI+pS5UFY+Beqh7w7RsEIQxGnqjCNGkT8Ox6PL85gnT6UTLs0s3UmBRO3o1tpi9Z/awqsP+rXnId
ueqM7Xguh4N/8SFi6lNz65dV/ycvqS98B+Gw0UXhdkHDo7UETJCXBDe3vbyjnOwLG9pKTlWfMh65
w+EF7l4GZioIr9Ayb0N2P2tVD+/FHnPsUCbk8f5QeN+4TM6SbFwkYrHpSF8YNVZZcn/X/8YKi1jR
Ykw04+v0rcirBb2QpB0FpE6mLzXj/sjKtJxRE4Y6mGccRUlFAX2ZF7agMl07YU1nwnYHKk0jLayP
koUPQHcu3fLx7ohVLm0X/7DspoQSPf2yow4gqZA9nD66wUoSzLswCB1juFhLChoFG1YzsyEszY7v
MNXKVtu2Jkxcyv+/875LhQ/zahJ+vvZgCL/8IWTclD003/TUPZt1KAaGdCpm9keY15z9ASU/6CRy
v/zNLjK0HsO0hQI+/ktaJMZsKoizNXFTZwhX/q8j8f7jfHH/dlG2jua3Lxl948LVXghklcYHsz0E
N5AE4yfUe+UbcmVxjsTU0Y4Q5PtzZc6kTJghBf3Qd9tGMlBwBhMzXyGnacytXZv3L8PVBbPkSvp7
/pyKoygvKw7jBqR+Xlu4PXK25P0V3XFuNKXZSdc1tZRPUY4KrcvrIIFJ7DDlYnoI2g2O6CRYggrO
BclFZoCKauaN4oEX0HMyOHBTkEQ+i+tZG0OpqJ3sRZmDCr80JlcUY7cDBBl2X5IMOOlvFsPe+53Q
rvFc/xgB5/7DtvC4NASAQqf0hoCtOJaWmtWpVo+siCnkvoD3w5UeWjsOq0GT98zPXis09R1tEr+5
W7ZB5VFU99JEI4EhXmZ/PbGRqOT+DNXGhaWu7S7gF5P5/+oF91vVPFUQyx+y1B0KWUXlx2JH1IE6
s/+b01fm7kq494uxHBtBZqQj/Q7gC6TyTsR2g7+07ED+M+PIjuYaFwsw1ZWHP/TPKqe0i5t0EaCk
Fxf++g/LAM2tnTTg+jqHq2MVC6GB+fOk6vJ3kkJsMnUa177lXsOUq56KSzTwpowoBpe06HMbVJIb
wg8NejdBSOomSj3ZzUs8IIffgf67k7aSWUk6Cn4Yk680PdF5EFTOizybUcYAJBq0jmkQGXZlS3E3
dQq88CokyoBJCABCDDBK2QHS8wAjj5U09ScAOZsHF3eL7vGh9z8/0J77x/uuIgNxRiYF03KbMjVQ
wGpQCPkydXr0SsaLl56xrnM0DDYi7Vmc1Tamd+CSRBwYtl3gtMknPiY6R7sueQ6k8IE/je7QP2EZ
2DtafXO1znwKujhCrOeBWP8depK53uk5df5YZVk2k1M/inoFPB3IwyL8SmmPY7T+rxx/B72Gk3t7
41qm/EOyX5J6uDxOJeS40odcwcwCADKsw3C79/ZRWIxntFaL16ckIJ+PgWtLrXEAyJsqrRvUSVFz
LyAKiW/HxMtJDC+QZMaGUGhWhp8icZsPeH6xrUDMCxZIMmBe3hq6DTC3ibcWh7/d/ajDXJry0YPj
bPp/TIoTex+vw4yBFQJ4z3Amc96B9UH5GlOkfbonhpzelXsPPbjU5aCqCQApgfXo1A77Xw5qESJb
48SWS57qmD/Om1K4Ns1djeA8qzkbznq9JtuK638vWEZfxZjqWdcp+K37L+IfGIYjCE+xa3vcIR/R
FR6OtVK0AscQ7QNjki3LOXyKv3s8qy6LHT6rXIOVMSyAXZwpXtaokaSrFlEJLCredLhgZYHiUS/Q
GM7oLh6thEiAo6r9LZ2Ok7MonaU1IdwIVGn256Z7qExxtfuIFcJ5ML7Ify3DIa45S5IxULYzSiqP
n6Ai6FjxECHiNesha8kxHkAgyRfLk+i5DGXu0/rEMne+ZEhVoCm2HHfaTmT3C7/bmzsH9pEhA7pa
I5iH3g+HWed9BsNLufsaqu7pozPAyFySa25E4oxzELKnhEJLcmfP9aCihb1YxR5rYVXVLSkcHn3k
vZGC6aBZnMwmfac3Qn1xn8VJEUr/2UO1DZu4Em/m+dfoSiQqZ/qBgV/5blFWV/wA4VLQweD6saST
LzL7W3PAC0PEHWUedC/8QD/IQg/+Yt/eu5wM0ID3tJbiUK5LdWfleMdLtGEk8nkkRu4zVznjODeG
m+9opRmPjRVPX4LHUQv9JNt2qelt0p183QjTWWCKMTdT/D+y/YFRl4bknLfHz7+CcioaVoS22v+w
PbjWumNnE+e0L/zIQGVlWtrGbdZiFtq1Oe/tGEY5VfldAsNHZerVCccLzkdTs33lltuN16PgijwJ
1vnoqCGQksNjL/0u+Byc19E/73vJTXJBdfs6BbFzmDrGF+tNKkoV+DGbKR8YU+0yWm2H9ZPDjdkj
6v4/3VXvYfpL9ld456MqZzFqtw+2yUkJwkjnMmC4XtQrcaxftCOf+GlCkNqvBlnYj38UUaVPmEB1
R7N3tk9bUAnY9GI+ImJXIRO1dnC9O8aHGgktO/cdf3+H1PRB4wiTens4dM/Rxuf6Gp1KNHsSg6sX
9UVhBThMGWjvAB5gLTW+QC4e9SJslt2bVjGR7r4PkCtGoT5H3lBlMoFEcEnOq0CqsFNAIF/qsH0x
cC6jehF4KLgj0RjiJxHMVeY9M+yLCu5YMAXuyHUwYBFb5g+22f240eCHqUVuqacod5l4Q1uDu17J
mU1h+UsbedURfSJPPYWp+4dbYceedUE01FLnfcP8nEOT3kJPeO4ZhRbmWkcSb19pw86pvQqGavD2
Qz3S8CNFKpHNz/56/iAaTnxQf2WLvRov8BPnu6dQt5ZP+d2IwrKGhB5RM7OHsXtElqkXbtJb0SIg
8hU1EMK4FznPQmh+islMshk1GWJw9G4up5FwqXnLHPiS1879Rb8QNIGQ1aIgJvaZwQxec1WZKanN
5+G9z3n30sE5+em5lgKls9x/O/N9xsIB5sXhWfdXgiR2EWwrbzCAp522TRMLoTEckBWYWd7pdKbt
sljsQ6O4/qP+eJEPgCylPIa6LmJV1QXU6lPBUhrJImBYFz7XQRI6YkrKTl0h2K0wsR/m9ym9Eqgp
UJq76CV6yjAGYe5b64lsxnSxUFzI3V5NmKlPm4KgEqaxY9dzDSN2MUomBzmG+Em6MQKug8ZL0vzg
brw/bUXjYrEtTr2sbjW1yhxK9TtCuxZU3yVlzm8/9MaOUTkZOwCNhgNBgFLj1NjlT8e+Z5zjXvwT
lFeE7Gw/Kbz3q4z/atxFHlrOi7+BAuCBhyBYW29cLt3hBbNPiaGkpFwfhZhZKrsCvp1glrsNZ3Hh
nQxreorR4yiYVcZx408LugdTtLP74KcxuEKUy3Qd03S/jdS+QW+2g1twITd7AAiMmiVS+lxvqWbG
He/OWpJZAlX6NSSFXD113r2TyBpMJWUVpElWtUpW/zvblTPEUkY6lAyhS4qJPZmMrXpdKlK/asXb
ojUq9PaTNNfJmbzr2I7iLIiApfaBfQ5GaPvI2Mb1/yFa3qpKDd8OIY5qsqF97UDCgb2eMlE5qr3H
esArONt3d2FxI684dxES77EENufoYKusZaVYspZdG4b/M9e9Cd0hMYsglg/7eIgN1pPN2Dd0YO2g
lFk23QNDarJasQJWSCtlHExij6JQOjckluzk5a77gn01Ju6XV9dlb6lMp2NwucNQSWBVByn9MiRk
G7G1abigIhQQiWA5hz8/KrtiOYx8vTQ77POIfYOueqCctz6eOcTXfa6HyUYJo4CiJ9n2oMp/B/Yd
29/rYzBfc0LubZfDv0tOIgO2HvJSPgJNluo504Re/AMCK7TLUEGrbefd6mj1E6yUDxAtlncKAp9G
eM/lx9GUT+UTwvKL6zrp7OBpwPmdJqwjKQOPEQp8ofU/fsFvL5AB9Ro54qvTfgLIB4d2AliTtj8D
f/Dj0ZFhttqmCW12NGBYokaI+vxcWAU5Ei1DoHuqUoN4TDkdCC7/cGZknoO7eQwGlRHCp0X+WdMM
D3DIFHC1stOHjN0EJd4c+yLI+saIMXg2zWst7CO2spCvT52DwKkzQ5gxZ7X+yQX5J2SJN2/0Xho3
IvhEZdy+hQCcSNv+SwebJhnTSMvD+cmt9gc+CINjldIra8R8tDpGmhJ4Y5TCNJphTaVMMHkvo4ok
tXmtPALEm9V7Z1TX/14U8FJbfhw9+O2jSUBEdFj+l1at1Ti4b4bA1uIdgdg0PodpTxgHMeIKq6Wd
KAtMooPNF9/bVZqfcu6+o8CKv7TSjXCYNPOcselcZExKJ6Bl0P4Y/8gpmRNOeURxp0HjdpxNlppc
g1h4d/0P+CGbArCeI5xzsgf4r3+uBIzhnLuPhcUfbAFaLuCGWBAn1gIT1tn0i+EoL1KJJmhJW6F+
+8dfy95teaywXi2FjzGAJyATb0jSneG6sraEd+irQTeVmfJgb2XunumxCSUvElA6gqGzcvvXI6qY
tue4/eQOFy7uuCJu5OmSMhX6Tb7ct0VXV45IJ8Eh+UrIyNciCoRICztDTX5YWrAKHdz1L6QZAfle
GC9n11PUuilGazzg5G+QtrwFMk52NyQ1Fnrz2ojMzxNWfl6/xdp/P0WEV702ewN+NrLOB0kjpjVt
ZF2H3bqEtgkpfJDVcDIux6MG3VwhBhk9xk2eptHEyd9DW+xBFlqCKMLeyd9jeHGaK/Sg9F2ek11r
wGgt7ZjxCXHMSpPTh4h7KEgVPllaU66LRcltazd7iPNnyYIYuWshsYRzKZcpCzYVXwlzZ6x3Kiht
plTVWrL1EEMV6vb+RkQriRU+4WMGjbJmouxhHojQ92SV/DXMHD9uBphDyohk8yQNTzTuWJ2a8bLJ
uLB/sl1UDaDvAbuojujtvlN7PaVdOuT4eyE9cN+s+mpFHp4qoM0MnpXE7jzrHUvII2s8GeushZxF
Q4wQsJi401BJtF76djkqXwAXh8zFZ5EG1eEFVnVI/XT+tb9TGHkyJ3rHBKBn2W3pKyrQWdbTLktW
fZD/A1RfiQl24N18gHyTVI1z9fVz0yaE0Vo7t6tjhxWZ2zr2O3PBgCJz3rYM8iwqzDItk7vBNjNa
qrGdX5aDiW1Z4k/3T32G5Kvy8bZazsNo0OoXdiJt9AXFi0lH4NcDXqk0eB+DtaAREGajO/ho0BQc
TdD1e3SDRMWHKnb+JGi/AhGsTsSH5MAbV/IENvO0SiAyAKTcTiEJ1RaDrl6JGiaLYNWlBXZlLgp9
Qh4IK0870Uw0yRhdwY5SNQvyc9qgwW36fE6PDyvOHsUI150aEhhSP+SKHT+tbxE+78V+magxiulf
q9kB6hR9fvW56kSuEdzCUqfwOQFEI29vBo0cRKMe+FVHlQLilPJ0nxASPlIu85rzUsT9LDMOErLT
rBT+RsLwQg/wj2XeANwNGVN+lv/ORgxaUTtOCsov4UcLXTmbxl8bxG2YyHYB6YDKA7RYr9YfWrDw
yYJ9ewWrCmuIGd06IUuenBVw5pQsBfk8kFA07zQuHVnRZSOaBbwJn4Kuc/wdKNoiG8dGyg+I60dC
5YS5TCCNj9LvaFBSByDRCwTyPZt129SjgEu9RF/LOD8vzGVwSJfmg2PyXc8O7X1hnKiAnGNV4d/B
oi/oFl4RYjJXJMuyIMJ8IlNwTqvDsHlHyEl7aMy3fSXi86VbZnagyd1ZWT/coJAjVYNtODZNUbw5
mwwV1TuBauShK+wLlujXoaeJ1j69iGsNAN6Glo1Ywpby0QGUhpJc/UM2wtLFm3TQPu8CuxEtKFmI
KhurYWZ0nhDxyF5ZI67OR87vppfyDLzsFk1Jiz4WaH1rPP+dTDd7dFGnCNjWVkQ0PPQct+EkIL8E
42lC/VWvhMCjS5GWmyBpjO+PZoOffK3zRB5JVaShxbv4Ozplxbb3lPHcaGZ61ZwnquSvMrd4kD3p
ezhCPc+1MIElaf8Z2+o78UW8VIWJHex0FvDeMm5L9w2lJEq5qy6U1aTsvBh++HEV9ZSLvcp8jb+o
snH4VaydEbn0Fof+gDqsHULglRZBqlpY/s4mY4zUvAJtDXid3Hl3SisjRY+bJPmCDppElnCrF7ZX
ZD9nwuCeIW3Ipf8Z2j2UUdl3D/B4VzqNPQZ83oSU1fYj17S00R5a8AL2yB5Wna0XGOr01vjKoBSu
VaYc7kDw7FTzbaIkwX1evl9TJF2JnVeSj6dwUnYrPF1yaYsqR023llH3ZsorCCA1pwjQdqheMSKx
1yNPk4wYcAz3mB/goG+aHRwDdgb/5r2E/iDcrYIVTn55XAgBeJFxZvjBS2e2h1XfIuIfWL/Ws9Ue
8zLAksWQ1Fi9fEnTtqujTouzq2b2yYEyr4Gb7E0jjBtUPnKGKLvDCupeMzLqY4fjFw5bV8S/hsQC
8cgfsPoBDRKEjvfRE5dBQq7UUbc/LWNXO0giyyoc7SO6SFAFLPKW6kYISS2SOrFasEX5YZ1A0QNy
wf8TmS+rT6HE6UK1fim8ECyIhc0PwGXZouW7G1HDaMBmM7dMV0KX227J1I1yLAy7MQHBP3dz8opF
VLg0snb1MTT/awlOj25JWsOjTE7skNZoVQnCdHcln+isyI0R5QVF6n6om+UzurrZ011qfLIPf7cn
KZrAdBLLDRIMVsOu5UZbXRiauHwz+8RWe7xpIgi+WvdkXjs5fIoYKWDfO7JmbuxuafeZF5BowzED
dVZsWJ5CBJSv9BbI7Fjate4cSlycvOMaNX64wBZCdZ6YRE1c5IMUXnOiGI1nknWbhz0HEIvO5odt
n3nBBgvKp+omW47r0Cfv0I/GJHixhDs2FbNhGLhNOHAcMnL2zQQKURr5DM7ZvUda7ToMyiArZMml
iV5HYwsW0GRh72xBo4Zf34DdjBhxUrkztcdjA0t+I1iuMvX4y/F1ME8U9m1Rm0QU+hIPfgmd2RAw
XCqcl1DM9fMaPHhlNjVnFztDNSJHI+FGraGM/9xiedStDom/IhI3TCpwreOCdWP9968aQg/Yj1hb
7ovlbtagGz85KbyMofjU3p3QrPl3DSi5IGWMsDVmwZw70dsoKCGBPkFZ7exSQqM4Ta9VxzHBAQrT
RFlUBLDH19Y5p2wfCgVdlIS4DdQJ38lsbHXTJpzBnalxkqPeWrQG0ax5uKESwvdAW4/xnDFn6yeF
CY+riwRPB6OGCY7KhcgGvglYaVjWATjPcnSwMR32C7ZqyaRnyR7lBGfUCkjlVlaG05eVJz8G8YNm
Cg0fhYdlorejOko3Bn6cyOXR7mMH8+LTb77dvuGhnSUvchpI4OCDJNle0524ItPpyGqQspig/CHk
mYeR+gHhLlvknbBMFJ7xwf1ITLEM0eSbS3eBwirKuQ/PAPw9ox57I5iFqRBgWNxmbQM5P7SqG+aS
G9TfPbTKd7lfqQOZJREVH5pdNpl1Rdl1R7w3HFPFj8TalXbrNPTN5as4k86pIMhds9xLQ1cC4MzB
J02iyUQaRS4ENqQkU6y08jzI92/4Mv75QN4jhG8frCLdX83tTDocBxMEOSb8mZGEPxO6tv9Xa0W6
VdxNnBczT04EwL2Rx1t7crJRle9jNmwyp+pBqwY3ZQMJfWO0dd0yvPGKS98k8OEE4i19kbm/UqwK
F1VHTLVxp3fFTQHySFaJ1D58qs2GPLatpIDFWdfXLDCu/OhI+3cFEgXHymSHIdyvGD7JcunfGQjj
Pe4x+wEv+ZloxwdjNGMDFpARqOSnMdJi0z+Qzh4joRxKXQKlbN00t7n7k4yJsjbLfc/W2AkceeeN
u3+MZVb8A2De3m+rKXW6RJwO3HC4qhEiCbtDwrwTxjfPPCq5AvtfTcNXF+GPf8vLGleWR3aSUlng
LWeQA7ukBlvaPM/EmNmFDLqTMp3fwBHUM72R6U80o/Ro+5BFZvyMfSDLYC+PxLt8FrYtSfN0sKPH
EZHIQS2DRu0rTkTHxvSQB/cLg/PybxwZrQGPB32fG27NkPHUqZ1JDM3upqbyC2pTK0yZbYvkBMB9
kc1nBL5KNC6K6jP8YV4pbBmoNwsVv4446nUUKzcdAGE6OvSPpG/RwxdzjkO/Rgekm8BpdSe7dvaM
YMGxCQ7r5xNk13KUIG73MK/FPdqbZ7u/XgcwNcb4GIpsIZKfkX1l1ydGtqIT19QnMOijpqLVm/a/
bK9Km1YqTn4qaoHjw9/Yc1cbU+OZBT+FpAnxqsygp8hNljEI5y+C5Iu8TvjfxJyz7vVkHFgvxBXP
Ml324yhabzyZFNyPd0zZfJUQ0yKRd9/5q7zxc11Ot4ka28Lq+cfDWlLubB/QK3bSZ0jgtVrplpmC
qrZwjEx8B+5B6tVmu1Andzy+ZPsIhkU7Oc/P/okOocet/b2arlBc8CprXYwNG1bhd9gRy/vktHgj
5sRlilma6rO2oV/PIiFNv1IhAKMnDm3vJ86xTidoFE1m8JyfH/lE2pdu4HA4O+PT0v5BlDX/8HA6
Avkq8gpNIbW3HMym7n9chhaxvF1o8KYh+9Ukmbc7CeuRS0ukudaYEZzXJUlvelmwHoA/kIXwQ1Tr
Xwa6OpjMpAOEpoVoEnkFA3M1PsAyT57F42r85FdOdng7W+Ci2/URfAvh37VFtyUafG8C4+Ix6ehH
unhIKkWVjmyTWSadvOm/mU1sN/Ofc+4JdKVEfccPNnV/xvnbHoQwXr6s9jR9z81jywaNEL4rBctI
go/JiS6zHsBSP44pW93nb5d0Z7eBksoqAskFDlB22GR5SdIYRhzjCcdToOW9hXyV6OsQ13utiNJg
wGJdJR/CBplMC35I2DnFzAHbuyWjNXDe2rpex8/Lc2InSKIQhiyy2Q5chhnhr3Kd5OIKJi1AF7Rm
sKQYq9vTT9M5aUo/wUATQPIwYgAIrtWcq9EYTMpxMpNt1rxxBl7K2dsBDa3Lr9j1+gSAq1u+ROqO
lZUdN/p1b85GmMGQsDksiBI+MZtOgPhK5bQsZH0iOT8DZW6t8AO6MDA6gsRcvyF7h6OsTXUJqAQC
SATZOPwzOcPbdv59zjk6kq40ttLORbwkXQCzlmtq6QkI8Lp/Kn5mDfQVqI7Cqcuye3yQVPyhW1NB
pMB8C/fqRfXJxCUdhfh4UX16oLnU3Hj3E2NCgtRz+CokijIByUZI97TzTevUcWPKdirrapQUS0M5
RnlSxUDB81IVpUWb1uwGQXG3h54b52ZqvhekTiFACFLuXSx7h5EZvVEG1vVtrGgLby9R8b7jySCE
dCQKYUfpchBN8IGnTgleofw8xIH3nATPUxClbRsPAByG9SFj9ByX568YyYu3tNQ2jPYF1lxBd1He
sXmJ/uL9u4ZOtDASGEOmePHj4O+BE50XucjJ3rx3/DqfSzR2hTaKwArFwfOmy+oSo94+OxApi4lv
quFYeqktZP55k0fNuwwBm2w4pZcmFXc0/G/MaY/zIC8y1/D9ZC773RuOIAEHtTCshFFzIo/KiIsy
sMTMfcX32/wfTUJqGB135ddbleGuBO93B6ybxKu41CneE8OpMjxCe+zwzBMa4vajVxYgr6Od438Y
kZmJiHvCjyJK1vFAbd669OXU5fWJ8qf4kpmNgbQcS33laO74dzisA7UfUfS+k89szFt37QYKMLsW
Uq5d1NrUggGBfc8DBnNszrjxW/yyIphKKhRK9Ozytpx9nIi+IHT9SqZLsiEcA+l5VO/MG/haZjz3
NEnDzRFB7dC3w4JOQSUvsHleBaW46C4GyrF7uxScq8bTpok7l2prA03dmJAvkeNKIK/apncPAHty
wbgESVhIXsRowh28W6K34RWGPDImp80sepO4AaMKrukT9VvqLHreTHNEmbfPzAvnJVJDrb7M4qO2
2qDjzICEKTsjvlhGrojgWOXXs9CBPWFw8x+joDkCEm20wC/dzdC7L9TKf259GoSJLTLiojLPsNSW
W7qUzKSyiAxW6nRacmbQ0VVL/rG+XpAH6eN+RhvQFV0Ui9Qdt1BWzRYj7GVIB/DxIWGNKBy/rSo+
gZ5Eb9PYOvUkmECjR/Cp8PygdeX6qQgl75ojCeur0JdzljHg4B1ygDnhTEWLvLyfSg3XnMRjsYHQ
MJmUOcyjR3aYOA1AZnmmUfYnJrH3kT7T1Lr4jWp7rFPut//CZH8Ri+jak4MSKeybkk+pWI+Jc8k6
/zvF9MtYCy0Sxbw4pSkQvW06v+Y5eBn8Bkp4Q9qMStIQwC94VmhhFjCxaE+yXKwgUzv1gw4h4W6+
UtsYS9jeNSwrO+Kfy6wDg+f3h5e7+OAtpcKim+vLjKUwSo/KXX0eq9P2kFSCoT+FCLoBbGOQ0mK1
Wcomw48vmCV1O8jfth+bTxtAaFy/VX0BzrYb96c53jb6s/NakhMlJ6jXWG83D3yTNiEF+loTRnRL
IypvGq3CVU4gTvbdJLPJUMylnbJ97rjv81xheUjJmq4/+AiTLaDRUPMO29ZqDwXFtM7kcVvZxNdV
jQ3hm4PRVAjRwuRxRl2ss59rE2nUZcVqOEMpKNExEV2X+cbzpE6TXrZoLDPtaHQyKlGKxypKnDHQ
kIvWNEgN47uKtA0iqBrCk4iOH0EDJ3lmevz2UrhFAJk/36yxDJDJsW0ghB0f8zRtVhz/R33IWDL6
XdtdydyzoyGhG95cY9eucqNqHTVXl1vIlYCY2+k6T9tnnuwGZCIsV71aHBjpCCww1nkmQjxFjL1Q
hmu8MhBMH7FvS89CloHWqxN4myald9ZxrOgO0zucB/Y5/fKMhb3ge/tIIqouY6x/Op8zNDM0u/sF
44IEL/LK5dBchKIvqIQV/ih0OGazXnTt3vkDDEynLVDIkcDRyvFAyr4m3jvYd8/onduSngbEPGZH
rXHTEUqEGl72piPlT1nkJp/NGeiR9aDOSKzYiU5roN4it0Dro4mol0i38Du7G3zIN+gtVPWYNhHF
fRNNm3ELvTdz3vgtuX6YWFHhPg4nV6IlixDSoX+nc0m7ULaYZl1n/f0bWk/1lL46+kXdO1O5MMjL
qqDKn2LclZie8TEIz2ar/Zs69lpo4Q7kvdZSJp7Ocr5TokrmWBXpoI8aQEReTeQBUmvarL1AH2EC
q995Upk03BPM6ZqR6X0AMTRfMlyrSKHF/1EBz3ELJc07MlAtBeCfZCsLjV9Eo7mtbOZmZ116z/iw
XWbsF3go9eM/Xe/3ZWxJb9Vg7eM5Upfoq1v36Odykk73aSPjEOgi5xnFbxI1uJmKK1y0R2a63bbK
BE3jlLeK+WhJmUt1+ZEQAJ/LyaKxKSrY88/8CQ1Enag9T0e8tRXvJmkAoQPyKWsXwO7OI/U5elti
tR+jNh4E33/TnM892CUVSBl+45RT2N1T6Zv1bpmYZC9DgTjp93yhnn3Q0349/ogU9bmlniwVYarz
el5Nn9aZ3z4MhEGSc5Pb79QR+F+1usthc90vRe8sfY+kYYBseC+wj/KuHJcJDjMhy0RMaw5IhMP5
p8i8MnbnZSAQOaQv0XF2mcmPhZ+ZN7vCubAwWHngi2ZhZ6wLzJn60jOPGlEInI5eM6U/aCkTje78
WkET4G0IiCQWlhOou99X7AcYlzcvRgEDS/E7/vZDRj8wc6ykTlHTJ/LsH5rJRZRRDYx/wDqcVN1a
/UOSx25maPDZD6zgrG5I4b77Sprv6eStBjnL1gK89mtGuD8cXcvmohxbYje11CXML8gfwu5FXBes
d8FqphaOteQPVD7lLG6WjeeoqbLN8mTbAFka8/6SQZ786+WYvYGioRcYf4CCgyp0cMEH4xaDjVxE
v1wq54RRNlYJq27sBaFuLJll/oxXVlau2yeiYkEfqGDmUx6uR39OxBEMbwUFK3ZmYg+xWwYnoh7M
2Xhr+5dEXY07nwOfmM5wLlzvAJm/dRGKCQAz4WVP9vTNEer1UMfcsM/KVGn7UQttYwQTEVa4zxcZ
Bte4tOtzFoY/KrcaWZbORwQ8xhiK67nCfESVEZY58eIfdberJ/zLPTkK1DHsJHFT0jB/sfaWG07P
SFmkrTzitucGBTdU/bRrzA9I3UT/xmXJ+/7BOi2Yy/MVQS1QIziuGTvubNYlr0ClhBVzf2UPEoZm
Klo0a+GAbg9xPIz+DKCFfm055N7QJhvIzyMqci00KlWO+0SGWvhpRjESbGEoY+kC/L1PAq9e4WmD
2N08gqGDNB/R2Ssx7OP82LZAyGfcDxxctb2f4bc8IhISv2JXZg/+LrXBWSM+bGH6OvshVS/57nwp
86KnecbRYC4VKpXu/liF+/CCf7R/bfk3+Bu6S87y/kodQcRO471GraionG4gBtjBZOpjBQFHt1I0
exJ73cJnHheohMmkMCZUwQvaxUQrCNFciSdaqzI/pT5pXI5CViQ24s9CDOuHseqBeO5h1ER/Ihb0
wZlBw5pC+niLUE37NVQimnuf3lEGdQdm1WTyd8EvqTsR/NMYs5+r8w3ZBa7RWGHOso+y1mnVQwDe
LXlU+eaQvFrIJcSxP1cDN6qqxhTkacPNiFj7PSwxT5f5P9cP0TyEdfN1NqH/k4m6cJ0cWTDbAaNI
WicntUbIbSRyIToojLxplqAq4OoSgHSMkEYRjW0PkazmhkEabKPoNOZgIqknlZJxIqXSjww6hZpi
9jkHMbv6Jfv2rgziS5g6xIiGPLuWcixWfI0EV8LZaWksgT3tl+7xdOQYUZXsU9RzjgEIYFmf0aWZ
Uo10uGb0Ips4git88NfPw+nAgh1mAjHyOuCEtePDIXCIFtSmAYRmhy9KWPm5hM6xpXs3UCB+4eIe
SD4llm2x4qbaDiFuzKHX80wIT9e/yLGarzzvug9O/Ge2bArtw6LUQmL+X7PRxo9d2KsLpyMUf+Jc
whUk7BCk+cv0IAKtU55Q/idmf2yax+khlst1jW1bmi7F8+zaB3wCJfLw+M613l7P2Ys8rGET0BvT
6w01uPrKzmSWUCXpHX+xyByhnLIFmmLPz9TVr4epKxZoJ26+AzJ9PhPBao7+gZxfxC615V48IXq0
v9zvNZN+LneTGAUZtEzkb3en9SlcZmOL3p6CdjTAZFRXtJEV7bV7/LD6QQlEpli3J/xSya90c1SI
fDWMw7wLhJzDSTtFyT2qFB2eIQIfzg1TSmkJlYoBU8gfS3ODyLi1fB+ol/dhn51hLYycMuudUqFN
RaML5gx17djbI5eHmNvpP7nDUR5Ms/cGnfzZPaIBSIkKALbNcAD/6oJYcVK7fRUSXNrW/uT5ygd3
4Y/bf49zUJh2+6PXtYb9tuqWZKezJCJVp6mUAxeNhGkPo6njhMS9h+Q7qiu0GeDAcWdeoSVtw2go
Qg08wl+ksr9YKM4tXoBwGjZ7gXefoSe9UR1+P/hLV/V3RNWgukIOEqfqQkCgdgFXoCfIp38px6WY
/vVbhsl1JKZj9/Ia8b3qa0rRuOKAkhTOlprwRjavIjZK1oRaRBVKJWJi+Gnkh/6p0wmtCfFDFTWq
pAqNI4exe7DgZQDmN6aZEWSWnpA7Y2GEZId0zLt832G8s4IxfKekKdqps/Axu3mvpHVmoPcbaVLk
ajvc1Tp2zD3jsJx4XtCB2DUt/t3GXB3myK3DofNum02l3i9lChWhEzR4wH1Ko1s+Veaa9DXSyOqW
V3nh0/fAqRFDeOpskvU212JsxsWOB9txWav1+1sfHXcLTuKcttpmcyDroSEI6UGBaUBw1HzuBqvf
x94Sz1771wPTOZ/7bveeqC0a5DwoLswYTPSnRXtaFoVRkZx8Um530yuLgW4U7aOyV2fmLBns9cb4
33kO6Q2dYyDdjF5dlxdmWf7q6+z/JSBR0Q6Zpra2ThBrH2YnHQ72u85aXpG+miZorFGPi3Ft02Jb
P22UE650VF9g78MCItt3B5Cyd+G1SS/ybOoJ4dzuWTCg/xFX+A/ka7l0ZDd4fxHb5y3cVukeaBvt
Np3WNiJxnETwHBPeZ0i4sEXGz75a2FNSGKIvWlX4rWuZhSHgd8A+Kz4kk0/cytfNcT4d7ny9RuJn
r8Ds6n+0+fOURIQjI+8f28hAOb5tz87A7ZuTvL+UiP9gj9RPbr9bvSPzdAPRg02lpCRUT/suZigJ
JX77czMV1ssnQU6PO8qbfOk7nD9vt8qGgtaIBg6QLA1or55n/2hpRywVJY6NN9thEGnXOozqkpsJ
Q34NeOOwQaXTZVW/Ey04UjnA3zvJmktBiGpbHlVzEW5J06dGI4d+T28BZ0qmmAh5p13oNYO18Du7
/qmdI7qEaMIjHRJDz6y67KTbqlXy+VXEZ2owpCuP/lJhHiH9fIPFu/b0wsEiKtT5eDfKZGOs9tFM
zzslSS4r0aUnqmsgOu/BgzIxpvo/lqPNn9NfhcFvxjlupowEU991voqsznQ0XyWkiYR53iMEI6vs
GZJ+JEDzVlSWyERlPjinTQNkXlLF5DVCcGSZezyYkr4eAK/K/M97D8onLUDobl24R2bCX+zmOHH+
WG/hghHRmjS1JiEciyvSCc/0LbHbRFOg24XyZ7xODMZOvZzjY+uzeZOVhjflNg9qQF0j8PER1shY
PQR+TRN0axPef77wPtAbwa5C9H1iHh5/bBSRuWsC4PwVvGumXdlxNmHkqfo/tq327TeAjjAAxSRE
lc4B9gBqmPhgYE19cB1LrNdh5nJszyfINCSI+sor9MPyodIBuYI0IC62xWKa865rBQawpJ/us+BY
6YLwWNZCCMDJa3WDktJ753Q1GdxlLRRJQZlDRE9pO8GWZH1a1d7AGFp3bZwP7LSII7HeOq+qK+QQ
O1RZ0FzomLOTMzdD6JbbJQA8W8SgfgeNH+g1nmJCaJCzAnhNQMd70vN3ojN/Csrn413fU+HjZPat
tUhvtlxqjdwISIBkDcBu2EqYZaYe+EHHAtiFE6ZWzUbpWD3TYH5mhT5OnUp5ofdSTYTsbv5XweGU
oQp5+lIwJhi4txMlrF5qFi+ZRlm9PRjVt2Axui+beblLDvLLQWF8b5ylMxePpO77He8gq4N+h+oR
Oxu8G+ry2O8+IiohxiiGMjlRAn+paWZabEb3Nil8Y5cEpvwtFL7dggl2e7x9H1+U8ysn07orysI4
YKjsymrVBr0VKjPfPKjyfow/SSxU2gA+gOq5WbkHnVqfnL+OT7mtm1nMfzoVBm1/ox/ym+I1v1tL
teZgSuIadH0T5G2+6dibIVrVgp0dm4TRDb8GkMOJcJuePuZEj5cvDzq2ctQhPD5h8A0C24NWxjx7
vTXVLmxvNP7yxyBiaCdRgeL0wWbT9b7KeaeaaXC1H1T/75UVec+5w7UkCZnSTH3znmSXjK6ZzKRC
/G7kLtucMcI/8vXHmvCfHTGJATXgGHKCIHnlMFPvj6h7aCAJLi5Uy6N391jER+LaeaLHZVW2wzGY
LwaMAyP7j0F5dC3xn+MyJOFreJ3u6YYdhu43QYbUvpdbaR7zA19Uo/FiLeM25D5PxbPtrqMuRe7V
WjrOJXsWM/kk4Tf8XNhaB35VfnI8Ajb4jFJTSoCvSzWwD2o3TdC6omkKg4TuJ8maKBruSwKKBPbm
oiLpL8R2E2O0BtnDQCW+Wg+2fonweJhA6LeRCwh3jxq+PnXSL8LaZxL+JQzoninXRN+/wgXoTfK6
FCgJWpTVLuol00D5sjrASttA0VwlJukwqnBbWGVH6aWtl+y/B0/xbmT1vB09SF33+4ekMY4PMtVW
l9yn4SHDGcXj81VbjWSIAGpNVquK0dhYlPlEmJ8LjFjdqpGx+bQKFeYuc57v6i08YuQ7iwfqI+hv
nVWabbfAevBKZW9a7x2GScYTHad08Y8CETo6ckF5Z/Z+Y9JbiQhflT8Nfl3mJMy/xI1FuR2S2XHv
LFdfnf8zK4b3obj3KmTDPatxFbkoP5mxlTXMKC5RAXYD61CxMk0tXVrC6+hFhkJrbyMAx2zFuHU4
5XeksRgcBmLjB64lU33e2oLai9qd6Tmxi6jEyeSWoInvuatw/WVbdGtJ2Pd4G35DQfh9WiP+nvy6
0WiC+vo/VBRk9DEYpSUnxc9eblQ+Cr4QOsPPDhH9ifRQRCiInFxufx8dJNeguSre7Nd+qXMKtXzs
+9CeOLkk1/AQ3+GjSyzi5DaBuSm5/p2+50ZTB6FozDOB2RNd8tKGcZJuxhAMd1aZq/HZjHdKvwuM
GtmjzbdmAatBcBpHmtDGlnmBEN3HGAoeKsiC5J060gHWwe2bi+pYeRhJQCyJFl54UhaI9XU7h14M
pu3wnv7sWVJah6RpTEfZn437B/GoWYlB9jpFZKonQvmJFad6NsWh9VS9N3F67PEknKJy46e61a9o
pMnIpP1vMwYlpW8tp+IXCkgcKHq01W1/R8Ccz7965FNvW3mYeXhUeMUj1fcms9EzTZrOMyap9IOd
PLOMUPGDm6V1kGlAk6vrd3krAfN1DDOZjLj/8FrzSatk5gq1soN5APFVTq86QRWRW4N/Jv5vqHPo
Ilg+X5cXz7kzf2cNXq5DkXyT0LnMHLo4WoP/wjAdZqS9XMqZID89kw8PriUPMuc/02SX/kLiKfdB
tIKIywb3Dk8EbUoM7k/wlxhhtZMveD1D41qfXHCLhCeWGPBT4Qr1UzhvIN0tv3HH8uHsFNgz24cO
CUQ6IC1iVFejP44BTjmVHebOUKKuphB5T5hmzARkVKRb7j32kSZAlzjIy1CtPObY23ML+TmfoOw9
WFNe1CcB0iNUNpzhSQ/keSYeIqIo3CQ+rqLJGmmRaZaJefQKnqlZnG7/uFRqxfy+4GGHx7Js/93x
/L9wX/vtSWeJybso7HAeBe4gUOnMUZGxOplFGf24wXBYNNknaRUS2s6qg0XYwNh81Hh7mPFgZZmY
dTODWn9O0PTTfs9u87Z6pHPTTNS55bPokn6yNHOXse/ucZ5lFkkTJBcJOW7mdTcusLDBkEyd91sV
56eG18NiT20Buqbeu2Nl9JpqwBt8WhG+znVGckBPibB+XSzFcS15YaN8s4Pb6MTkZX5sYSI2AlIl
gYFlKpHP56+ZKhek338gEapRYY+PbvW1AOw4PQYW4CsRO3nFrjknu8BNz7tB1pC1TYr+boSufZNd
lwRGrT21dUEqWEOK7jF1vW/GTScN6S//FXXX+JrV9AGXBUhx2Rt2fer2ih8seYOL7fC3cLMWJN8A
q2Jk3KE+EBYds2gOBtz/KG7Ale0Y1lndwHEakhYyQln0AjooqLbD6bBmVXuqewsLGuttuuDtwJtt
lw4+YaYB7dDqy75pxUc74QDJLytROSf0RQD49VxkJ8bAEjPLfciPSkyfKSOSCP1F+sNpmgUgWcfJ
VgUqIQrtv2Ec1s6J0sWJZ4N+ddD9BAr7TM27ynx23GaC0srUYZFfLKS4z2cQ+3dYzTyhhoiW4Vvu
n9RNaUrh5nWVuJRStFegCc4FF8P3G0b2pk4fXLbtsbwT4tz2pEkgRg72/ZOdKZ3JfzfcmJZYB75j
BcaLFo6pC6dDAlvI0x15CtqcxH15cIjxlXaiKtcX+KTfX7hHQA8LiWH1VGuq/VrO2glQkgGkVkNm
Cg2K+2w9Q/a3Rc/IJBkkMWtshYpmatZYxzNq2JckN9DlMhRLLvGcXxMLZDDVj/ERMC8LdmiN5Dij
jSEjQfzDNODPG1boYbBuC+bWaEmkjbWCeIMJgrBWZeljHqRuIurtH2i+5Z1278TbGiLxm2HI3XKO
a/zulUG4mDyLRW3iTqR+XeOYSV8jT2IF+cy/hDM9E5LfX3ntCy3SgOgLx5ZC+enZWlTlWMFYH0Y1
U1E+TbAVoLcY7+XN2xCQPpgCWAnMbd0yWSz797wmYIoqG7MhhAIlxV5pFOyodajfWhndC6cUgfT1
eOKt7GC38tc9+M41KoLORnxVKLSLr5YpWHNqU+VoGu8KMxpEub8LjGg8c/axY04D2PP36kxXbmcp
E3t05nks4bR1Kz/skVp5UOhUbujz6L/FaB2qA61YoBjBJw93Fn1CTcvciL87mI8moYJJ4G1C7cX0
EPu6LqBlAw9BtkAuLfeWCjzj2wTt4pO7DEdgiK/zMM6e5yzk39r2R23khjtwLf35Jp0Wh1ijkwPq
xFiXpc4fI6GwKHcXrkDB2ItB/3gYP+7pEsSKaeEPxXmQ+UpXw1DpIZ/SAqZSOn1aq9zkdK61d6wE
AhxUfOYmphCTuF1ODxLxaRUi18D1DreTdpOBHEgAE35+OxPFZ7K546yjWqApj+HyMCPJcDzrfHe9
3wkmS6Ul1O8FzPAD3/a16rCvV/RY6R1yT6A5tPJs+b4TfnNbR7m9eKg/0gWi+X5p1G7j3YgdJsED
zDaaAsVHt1F3u5UZlm+D3jempPbVNabDEiBvYBKvAmoDjLfHaJ/g91U4ppjEYYCVgmOJEWR+PgE5
AoBFsQ4EaoP24umTYv3Msfj44PicNZmvTirCvm2SEs3O3qmf4s7vRGpKJbDY19QgHxrovk0OVLx+
DiC0glwaXwdNxVNGdf4rmvu6QG/y0ze1KrDb0PyjqE18Ehn5npUTe7H7fU2i0iwLPiuBHpOoGnAv
vtwW43LkXCzgbiKP+MDEW9r7WbjTy2AgTMgN8ylXp5iz7BRRCgetXqnVgquR2FCRsrkyVs81Nii5
6IDNLM1XayH9gqJVs6XAYtT454YoMnCwEbCUQG1arrVurq58bO3MhI8Gd6ede84gGJhCONI40czh
dN+Se9VVgA7Ip+MQqvLBSi/NBBpeq2qMyGXDmqeFH8xHPzPVDGdlB23KCgSAemtDt+HYxG63KFHa
G+jMzD/NmtQmLxyGzQnk/OTD2dSmjKL8Rdc1cpJfjWtB2g93YjTuGH3siKKXCYsXsOBahg0Kqq/I
MTXdwH/BM4Hqoy7NviRXswUq39AYBWm6x1POJ6NsC+uNlEEwPxNUXUIl8O13AIyHAFAOBBaxgDWb
q/8V8IZAyj7hURQIEdVZXmwxzHLR56Uvvx2sMKNVc+DwZa0v96FX8wxVzVQJrOpIopnAVOkzDXiS
BYvO+iQC/nBcAZnddzC+/mAj+fAi67ZWdT3mu6Nh0jn2tiw/eXT6Tv0bPH0BO1yJQRt4rlXSTgHY
hFixN0OtrSlSTA/eGoES7b67zGarfgF/CI1dehyoZSWAVSKcl3XZxndhYo5hu/C/KopzCnvDOQkW
T2islgLJc7C8P2sBy2G7uoZp2r9rlZRpgaJlNR7q/F2H00xUIlW2gDaUd2vqgsry5MbGo/mKdtxu
bD9RtAkc9c9VZdgBiC3LdrTsB94KWrPkFcOgAetC6SHGobqsmGurlC7q3XdMh+M65Z+YZT1oBoMi
Vu06m/81dXzKMWe7TEeUzNFUQCxq1YfnY4pl1HjmO+Fbs6sGAVu06iWsjdZJ0TIilEPNdpYW499o
XTC81EJ4tt2XuXXa9C40iGQLPoBTAFbBf7X432UFFYRL7yIB6M7DM5ryqpdcv1WiTz7NI2h36IPz
s/ogNrTuRSw0x4r8GsOqYjXvSbSqlYLcpbb2zcQiwk1QTtlrixSCCuZSGRlOerUTTDZRdvx5Lr+C
zxwlkk2TwwO0Yr67GKU87GN7snjvH3e9UobOzYXF8CRZeRJVoVbhC7v0xRSLNz9Ur8q+uTXQutUK
ahoqOhgjDl1XismvywK2h6gNXaWFCw0kXq0eyS+HkliUU+cQrpF0BYWWVym2w2x85i5b92LNU8fK
xQROaAxzvt4++X5cji30bgGE/FcD28BeGyH7HZEe915BpZlXBD+UrWDfyM4fQr6wawnRezH+N7qY
xj6ehEAJFGHKheShF9b2DLTHSP1q1PJvSPScDX+b1torU4frrVS8dmaQ9D3K9G7pLiOKJ0ZlwTtX
WCxU/tdUjTK9ygGpRm2B5fovdHBffTsueqkBpCyYLKJ0XlbNnrHSkpcjn3VClv93+ceo0Qd6gP/X
C08AehWEoiHxGKs2SSthpN6XjkaYhbEFerKZzJ7oozKbg4McC/uHbxqR6YWSHAJjjeoRcK3b9F97
144xf0KJ3XnyyjjR0p0/0ehqx3HZ9V9pK6dUagBQORUJB+sXMg/S9aBxmuapm8CAarRL55iTyVN2
q8bhKM0gwyvTF1zVfPVsT56aOXjMkz7n+dA+MxckwRxfyJ32ROHFuxSdSMbHYQ23t2ljWDv0Djwl
Ttr8Z6wGYrZbjn1pUAZCarX3Y1cq/QXERXJifBJUVd1fOzyFDNnDWinldyFKBqaTXSU8foFAQXWe
KizHrXyC32Rgs+Gw72pGR/C5tgLPNoHUyhaxXRE7IRJmLkgTPQLdO2vPz4nCqJYHNfe3bV8MRNmc
gAxzrmcC7snh65kMzX443xQ48D7ru5lJLz/EFHhVLFePprxxZ0fZUTvBkTBSNUeSdBR30ONNZpJZ
KSFb0Iuzrr9M21M6wZOVaJXhUckLiLXFHkYHnxfsHn/f9JT6QYZf8ajBclk62T1EZaxUgrZcQtko
xQQfuzCXxdr5hMp4CfOiiwWg8HLiWGJ2L/kKPj4QhvOAEP+fjsYzY0VF8HKNDxNzvYsDQNo9Pyhy
l5V8FLn4ygThhjrVGev16Xw3o7PgexkhQvePDE+9UbRf7Eii3vrWu8aWryB/OGw30RAHIo8tCr4H
QtAaw/sPHpqbgbqsWmq4a98JUBOnU2JLWihWkNoGn19VfX2iZ12QApvKszY4KNtxtOERsHDhZCtv
tQ5uGvdN1cGPMPUgogNQ9a3J2TVyxDTV1+yL1VSETng9cENEGHNDRa7TmvPoHIYlT77oO5FAHYba
qobMlskUkf3GC6wZI+p7U3q++zKe7PjEE8eDxRJ7wsvGsUCDL/W8F7IPhMG3q3OUptCiEFqTbGn/
ax5g8MK0dkhVYktw87Nv4pB8vLb35ulE5r2TsqRbZ0V6D9agy0hbL/EaKyGlKcTrQfq0Huf0USTY
6euDQsYpBZDVAlSnWrYb3QKNJdWheEHZsdB3hMJ+zUANtmxtHFBAtNFqRkf/SH4qqYkG8JRNcjtA
wq+TakQaxOe4oNtk/5kAoiqYqCZitB+EXqm4o235DxfNeqv2OyU1xWIiix/XLyotnEr2h3tzpoQj
eAKCSY4r3CmiE1tTu4TNFFckollkOBBP3HLej0ekEN46Q0vRkq/t84ZUYxll62hoG9YOPxreo3MT
wDSFyYMRg6HiR1H33OLFuTn0kgcdC6BuL3bj5+KIJSUrEZQx3aAkUexA+v1Fa2joXGtcG0gs0FGv
KSESTqTpKNklqIFVYMRO4CI8FKF+IO6v9Fcap/UAx+nJ5Y06BGb8ElVNr5R6uAmVCorW//UpTPaw
Pb44KBvo+wrHqpeRjypCy5Zi+Csf2YWMCcUQ0kfdNYTx176fQ491TTOza8wNqifDfCdsyV0dkyxa
AEQMRdo0GmAiHfMx9qvSRI5qeWW6E9xtUSsRt0nMAGUnYsqiS6+FH8lJ4RMOunstX14VBwmJpscP
tpcvtMI0ezZL75+roq4I6WWGlfj9XXnw0gytOJo3VtIzkPL7Ih1WqpuGc2evv293FEywoj+96H7k
29GfExYxAmu3AoZNF2igmEMEO8JeSowIpx8iM6DJ2XhXn3qEwgA/MleG1PQf4ScKMJnmEL4ngGCE
v4XSiBS79uWF4wthugRYDRutPyu0feB3zM7HD6Nqtx2ryUlxfTWMbMw9YS91ChKCQ8bSEkSM/p9K
l+rzNfQ/zEm7DUgcSElp7PoYeEkhtHaAzBatmH1K9GN20runXrx+313KSm/zWi4XuZH8sUymdVg7
81JJjerVIdnEWXZ1GlAjuMMIjNtxQnpbhKZSCFTcuk46YlsFiVKyIdlpsEFm+HlSCZ0h14/diorI
n3eN12k6XlTypKu/h72Rp2x6ZzdTO8nCD/KgDa/CaMAlXiRqMwDAkuRiznxO/SzFXQKGcxVx8WiB
eMhd71RB/b7CQSAO0MCvEP/IGSHLLXi6MJD+aJBLUvOZ/RhtuNSd9zE6lzV5oND3hXsidSTFA+Xf
T2Kf7KvTPjRa3wOuaTGZOas+dHK2fkofc8FgRtnQqu02czhLWI0z0VPrtVgzXl1lS7OKSBnWET8s
lMR1ikAxWcfT2Wsn6bWrBblCqsGBTysmXj+oxErs6NL7P1wWSGPXMzwi0TBzxGFC+/gwEL6FVbYz
dYEut0KLZNXOMIYPDFEqOVgS8Ih4q+0Hz7imT2YyEGzFGubdCj0xcUUS7tSVl9+CIdBwTZZ7G/Mh
gAl7gxRxx8oHFlqN5COeP5hWr+pmv/Fjkzcnyv6sgf/G9Kf1XYhcTHDtEtm/idEircZV3T55+2lx
cqlFkLkf+Wr6meLgasliEEbQ8eg3hfTAq2Z+OQUsAu6m6VhWO+1HDDf3H6Rk+2aKGGm9PiBzbGuD
EPo0v2YFRbmM0asRbP6zwTqUmOv9bh/C10RgdxmI6qHdMHW2cZFESZsZmSAdD+z9aPefxfeWJZux
S0j07CfSDTdg2p5UUMLGs0o7dQiPCafDmow0tOa4f18Sy1GV4vmGS1z1sTuBTQPm5QQbBmeBHil3
ny6kr61jw/xA0upmC7otZrn7MJCKb+y5mVEQFphS+IxQwxRiOIMwIBuY+BIclPiDit2NtWb9mtiZ
6mGkBHztji6U9BSt4wVzpThna/VlL8TDhfjvNemE3eDvRymFhbA/k6DRqhFVttgRN2eWfRhMALXu
2/Ps9RpG4BD+anQUH/wnmGnDYdHEgQx/tS0xo3EmyXvEjMGUwB5dH48CiijgTgDqH4a91Mq5jqMK
D+rHmCVvlnl/4IVBy0fMPAELQJct5OFLIoYZpKWb+TkzrZElrtS9snZyQxviGHq3CPs88JEaW8Wr
3nDliNK6nElAJnd4IXjAhdnBrqJ3PGyVACS17tFlu/N8/w8JCFIq37DaTkTQr6/ftJcuDH06RfL5
H22689MqgozkGKTFtNRWckpTbufpJDRfwcRzjdkZLiIkAjhzJ2rhSeXBd8wytg4/K8NRS4jkV/r/
zBzyZuDN9r2MY0dcd5z1jTG74/awYRFwhkFjkRAuQPMHe5N0Tic0tQ1rLJDkDj1YX472Dj5rrsan
tzPYjcSEDDrzm/7HgJf6yepCHGzhoGikJTg/wfrsZkcEnSTxS+xdtYjbpqxftPSr6jaYuT3bDs+P
MieV5/QaB9XZpVdxM0x7d5cXfm9YrNZgzZOnWbeG/XklPkw2AZKhef2pSjZ81lnXga/JOHMGJ5e1
g6HPjG6k4lgnEI9SkzCWTz7M0poWYtVq/sqdI6IPSsCHqChSXX+MI5+SVBX8bXSrefvuaScPtTVg
2YXqput/H6EwkwrjRs+fq7fI46M7abNCiaGb8mK2cfUlQMhKK1PWtOLmB+NfK08bd2P9s4N8TM4k
xDt/zEG0I5dtU90QT284d+752xc2o5mP8J8GL33yXGn2MtacjJKBnwc9yQpm324hvlKHR9zNgPww
6R96sJx7dPnRvyJR93LU/UPElNSUypkz2ovbhnH2l91qEBQiP4Q58vUPM+NNUM1M1kIfBTxnE2D9
vROxVyikHyoVYrnGjfgmULFTiicGgF/rcTFovPpa2/hHIa2VB1iqsACJ8holHsssfGCOeLWTso+w
gO9Cq39lm1KXIClukt3S7L/wFgivKYhkaa9uAInXc1fVeoCAOUg2el2IN3qyQuGtJ6OjrxjjdxeP
rZNrK/oeFMdeZfleSqkQq+9rSxt7Zz7jEJlTYCIu8GpnUE5LESolfaZBK2nsrEKFw5xpiJDQuuzE
EVb3mPL3EtBHaqsOelpIQuSjYdVZ4lM9f1hzyo1VYpdqPWXfrdr//WOymR9tNxLpyYcfmLHv0NVz
Z83NuwK1RuMN6pHeoIdcrHGyXlEN7fTQXvKBTMKbQwDNEuKm3c60vOPnEGB3B6KqvGKtESUX+BGz
mr5NqjDkxvrPRk85w2TUBgQAp1dNbimkxiDGqlV+08vlrJSxAsbWrQDFq5N33aAQs6mHqEZKXzUl
NqRKCspkJq+VyoV/ubTLqQy0cjyPPD65og5nXW2mrDKpK7teYzXKonSiir2c6yzhAeoPBZPwsPRv
Y9VQPRy/EvfR0hBSZUdvL4fuT/vc3nJRLJI1NYTPiMFvDdZCeqwmxhxuFXlFl3SkSyZbFaVgk2VX
p5zSqbOI6Zq33u3fqztl9OwihKY6WLWhPXMAyl+1WTHePKIMF04mQP5POpe6wvNYMfX55skhSrZv
TujmURTpbn0XMxtSzMJTY7sCsTG6VE6RYO5ZXov35mWVdc62ib9cI8cVglwZZf2ReU0libID4MPG
mzfSR8FMxIbZ/PPU33qeXrb1Ygx0rnnFVpLaHLwEs8jCTul6hVrKdneil9EAavCHNRjFNbcEMs08
BiqpRqIX99+IBCgjk8ON3XxtcrlnFWZDXgn/w+ifd/XaTKkphAZSf5fGMWcpcLjttFRcmNv7Mndc
xAxtsBKJAvu+SdrvQCElO9bM6ELHxNxwzcBM9qvixwp1XfpHk+7R/n2djbGVEw1O39o4Afv8G3jA
0sKCTsLUtmQPrwrP69a2XWpTS4UHUq0mvBDDe4G0i8biq3PVQ42ohb5ZODNh5TNsgj6vJgsEkZ8n
HPU/du97rRqa1wz9TX/UXTk0KZuTx3j7+ERh1XapVJufIb6K6vbhTaJ1FBt3dxZbjl9DmO2mQnHe
URaBLGhZMSeXNapnTfEUsUzZNw7UGr00TdiG0mtlVekv75r0KdSXMaPni/49yGBu8X0ZsHQRNwSU
c2uYtpthAtrUWh8kh1KBoI865fy2bkTuF59SHeqbfERCagy1NPPucr8XGcQyQNlSilTlLIAN+WuG
F6xra7559HAIlAGz58TDIJef9jRb0QXvguqGD7ypJqOHdFM55eF6gqFdC7IyIPCSwljmlqhj9RSo
Nr0wNZA4pOMfbpE286PGELj+JVGVo4lsSWBAmxl54dGat+g8tpA92KGk9H+hUXR5WQq6YPgPsnC8
YU/g2ybeD2ELMC1xJCQKpeVF9+V9+96fKU0/r7S88r6SUREqqad7pz43jbo7QNsZ9nLssRvoZErU
KRmUGOGaekTjAgesVLOpA7GSzPDGR7mJIGCQAK2KHdoHMTuKM0SuHHltbkAwmiLHMqNWw5pkxrC2
jWN6wmvGQeKfWdxr8kZ7vw3iFWeLVbwurhbOejbpiJ1JgUmp3FYP1qfsD3HzUe0MaNwaDMrnotaj
MUG7tkrYhQRTpA84xdbQZYoCwRq30ZeO/wmjcCMp5XsIkXKDlN9xqfrzj/5mQRE6SitizWgZtgSu
g4c+c8Lyf3BHl72fG5QJxOdMnNtZIyuksrUg+fM7pndPsj7BG7p2H+Pphc7sjwSV9UHUB7HLnZ35
AeDHDpGAJ+j8G6662wY40wQDgSmkkgKI8uGv3IXh0cYI5D0egYSJVv1KqdZm33q4glFA9budPmdg
o9B88THDAlmkgMB3GqdAR1x2gxaWZMPKnI0tUYp/s5z40CAc6uvBmYdRfGUfU/poEDEfrtbbjwWm
qxu4IaAztpsfvbBNfQ1wrj5vyJsxToN9Aj4xLmHmUHEr1S1muwV0qa0nSlFSbzmZg3ETCcYlvER1
srxavibuPa7cZ/TUKzi17gcnXMsRt4vj/KdoZce/O4A6aDnbgu/vrxkMmtAkgmhMaog8sCmniaWq
iQjTN7FISIMCToFsFKF26BCxChD2+FwIfKJ2eQlSuFloH/RlTnO/H6TxtaNkmRqinEIliEeY70TV
14CQgtVbo0kAuIpWfw+4S2+PlvgNBAKlWu7KXkz0G8FvfweSFZnQmpnI0L47ypKB4L8CX9iTqBhV
2ypnh3CfqAr7rx0o4uXmLz2Ozr7KhZdd9HDzQga2qDgm+u4CbboKxng8tgCb8qcVvfnPBTLONGA5
xt4FzEOsgiijRbAeKP9tMlxLjbMgpXySAUPJbo6GFE+VhqRKPVrHF8aZDX1SIakDP4XROLI/DkZI
wOCPRddrFulBFWiF5Pa7TxFLiu/9JSIvUVN+ZDArvfPJXaYkoFpg4GdsJYdtgkj/28YgbOg7Ke2x
uK4exIBtXrUuWVHIe7AGirkkkFpDYlrNKyQw38cdkPMgQcsBigzxQnSIzS3Su/SSxv+hcGgRL7ub
mTd0206y51ow48sjrx0ycV2mFDJEq6xWusLj4bTbwjRZNbXo9F7UPMqYmSf/h99tAHNorGL4fZcL
Y9I827jKiSUIGqZBa8H+4oscNeTmcq4V1g4+nMwF8PU0thyNFEXv2/JAh2140x5/Ot9dhIVcXE8J
0vXSbChylY9njEYWTxBpZPrOnz7V4ltvAduh4yUIjTLUVW2pSVgaJUfF8/W0N9O/nlJq6dOe3OFU
VhU0aRz3X89fqhuHorFu0FtYFmHNLtFST3x3U6/FcwMUsKoU2YNhK5nkXfeyWCfuZ/S9Tyxr5bg9
cr7imU48Ga7t0x5iVMl0MCQjKQdLPPGWFjyprxrv+ym2gOJqTONiimEL5AInED2Je7o51yFLSWhU
FeNBUTxYhTkGLuivOuVTQQxFE959EMp/Gi/9TdJ7RHi2cvIgnFE8orwKLidpYj1B97FhJIN6PYbp
ZP+T4OGdenhrfnx4lUCXaEY4IEKrnAVgnfoCU5emkhAmhuKhpPzoyhhSuQDQhf26+TyrfkRFVDBF
VyqlGbHWghj8a3ocuFFak8VQH7TTQl0mHPnHTLroSJ8k8Op3+rZjhtosMuc33dgyl2eVrmoIBSgG
nthNsknO77PhbP4FtmM5Y+s04VRkHxEp167H3r2oAnhbgyd0YUagyxX7JdqcXJKyLPC721G9yc/T
gl9sfgx9LMjALDO+ri62+JJaiLJ5+b8MiDtO6Bgw2XruNEFf7XhmtULAK3rsHAXV4E7unhOGSmKb
vs4r35oBpycG5YqXxkDh5CnhguimgN0Er0u2I/jYcX5vBXWHJKB7v4Zyrf29NF7WKmavrw/7C5Pk
4Idu9fSrS6ZqkjhlNQK0Fyqpd6hmT0j7OTVgXTRwfoseuflMd32GLObVzh5CffkcGZZccQsX7Noi
DBTHx2fu9rUslbRuGJGPxGPzRGsXjasSBzsQmgWURDNhUgeHdO3Ktd5VKRTbz1bVysY9bIwvdxjD
zRDPerFMKK9YIkvuoXNS0UakqLBwKLOHxPt4/SLacZHWQgFFO+HAu10RkpKhpk3ZXzbz8EV1GpnW
PkMQwEdsgd7f5bAapyKdX1QcE3H8Rkhmyy9W0sa6KJGxwx7SyJgkEYPIu395LxzFocl6hQkhc+Jl
NugE7fLbuWoXj1WG4iGhY25sqJKWRzDZ0+JxmcLKkDySkSqF1ox7if3FiTTN2k7mGvr9bo8Hn2oW
FHdl9e9Or4UCogaLi8+yJPi2bQ+DTiriUD2oCLjV1mE+XMKBTEo3bfRuBIai6ubvwfD+NVoSwAgl
SYwfrR36UFsQvyukcyfsN3cNBlPbzwpAKLmk4ox25Bqxb1btvKq6he2kctADiqicmwufg262JZlV
8YF0JQny0EU4hGESm2W2KrfYe/dWkf2TN5iwlM19wuFUKPg75h89ZqcgFAY7SOKaHB7KyA412/2y
EoFk6OId2YO4Oo6PzfT5tpwfjUY9KB0kDuaxxqL+JSaotmLAel9I9JdLRUtXvW/ZeJ+B/zn6vcO1
VxKYnvGGPSozY/wA6NA4rq9dO9QGwnOINIZiuW2wXmCQOnRqUrtLOIz5IVTkhYYkd6I6rpePxekd
oscR85z5/e8CvdpiVKtAnnwqRMQAgNCL5ZNFKVNEdIu3XN/5aZO1wsPcCjsyZXz0LuyYauPaZ04q
IVonl/lfO+y/K87OvFFdpdHT3L0g6X2SBGgBj3a30IC1YRNgsMmI6vpBHyfHFQBnubWs3tLwxvls
tXMOPvfUe4NgbfolsmzBPTYDwJuMh9Vyh02fiZCFn5ZUNr2MLYkzV7IJ1wxC9/uMImryZmLAhEhY
6rlT4du+ADtPd3GUwhDU1SbkYW/FUrJ/XwxHtwi1AuSqbmLehPwrb/EZtw52RrcrScUmtroPaUAb
hOBPCazdmYaTkqNweOOz/5A0Bo06UnMLFyJKK6kIRTA9FPpjrUyqF9a6p/D91+K97ADvDUEq4Sl/
5BwRtkAsAbMZCSilhlC7dn9OESO0I0OhWG2RAcMtAsy4877Etpihz/wtYnqJDibBj/e+GkKsdWNh
0tvDE2WV8g6CCJ3Pdlvc1uHz3fMAHrdv7JShx5sZySOjbtmPeFQr+qALKU51/sfs+V991v/S3jSa
FnruAK1usrNKJuBfYBKoAyg6naQRAOSnXR0OY2SsS4u89t/S/690Dy3DBqKbyc4x6mLZrucDvPHO
Gb62RWhPLT0frkVYOLW4ZuRgMX7Z9pmRpr18adADv6gJ0eFczUqN/VGlo30VpF66UV+CmMOrjQ0J
ppxYfJtPVbV91jmFx+ENBiHbDHE2XxYMPinIT2ynS9LmzCsGf1pAIZnpLXMIhPsbAnNsheT0DNUY
W/heFdelNRivtxNXjKKoJD+abde7cbsTT6j6ftvoISoauMrlnIxdLiw6JSHARQpMiubXk+VPc91R
H1TY1YucWxCpm8xk0ToCr0soctlDyhQjML6XNcU0ofMZ7lUAQJhl0OIGNZNJ4axJNcojsX/wQRWy
+QCF+CuWBeb+aQf8YiXfRODRrT2RDUW9DUILcdX2brW2dbm6izSF/9464NTJGEuCY8t/ehlQLWba
6e9eJFdc/aeUMJZ2xnw9MiCBtN6c18r0l//J7GnzCp1xTs+UCqMC4M3C+VKIZ6/IleiQX0KdAaxT
4H1T+urr4tXNre2G968JMVQFi1UKhKsX8P/lxLkKKjB0Ajz98uEa+mzdWj/BefvRWX9wAHvSOB5c
DVlYd7sY5GaxxW7xvh7aIaJ0vt730+UmOm8vYfiQGeduE7kEz8N5x3hHmkxFBdjdHOFjpWyMaQwC
Z98qYLpl0BszrNLduxcmzTIBUxpOqlqUdt5/NOJCw5Jg++h5AW5WeHV2+b4hkL7GapZnwIc4uuWc
g0L+Ny30eet3O7Hd/TWmznsxzp5LK+haWKU2HQ+Q6ah/pk6/bOfT2WdyhJS4k97nGQxxjjA8pfT/
kV7lsVTOuF5cPJznV53pebbezwrli9ZeTnSW5cc7rWXotyAIUwz+fh6QCPEY4MFlvyZOtizUY1Wt
DRzwylt7SvEvTUudZ2XduyfsInhTMVK5FlwnsmT/ffcJajeewp2W0qo+44CzmiDgEKH+6/39KYUA
Z9iCyJTCQsi1LfmsznRfjyrk24+UH6T8SPW3mNKNw0J9FQDbVMqxP0y2Seaqr/Sz7d97nl+/1PyC
SqyowAy/wCmBIWjdkoOuZWHGNl9/xIlaGRYJLSuRybgf0Eou7hazNJLBSu3vp2Cbq852MO85R7dd
Uwas0s/zvdcr5+6/zINPzajZ1zwro5WHwX6m/kAWmF6O8aUxOqNCbcgThp9mhRaf646HcKCHFwMr
geupCcXdtGaAh5bvSkSRB8NTnQYNlGfjgsADiQN0BJ5iGdlFg6zMvS+gj86VuTI5ZopriCGcquSM
ZWIuic+HKeH+YlvLxIi11gNCXFSfNlz+yhqhYErHaZG/l1VkiGmPQ7MwxGQB2hI1nfcjj0KWd29e
KXs0Uw1l59Y7x4l6LFNpXMjcalk1UVOk8fFbGUkbI9Tp5XLAdszpyDPdyGRRXwQT2b+7GhZa/Cfv
eAJhwqT0JX1YR3Eplv9vGXPw4UpD883NOKkpJK2eoCN0VmmhqTMawxzOAuHbzs36dOb8Fz1P0dJo
NEDcAcUYr2O0ULb0DmyaGQFXovMUL4Pi0hIsJTxZgZ7zv4zMgfyBqJvxpBdH0pl7nztr7G7TZ5rt
pRnAsgBADmgXHMOt8/Ytyq/Ev9V23zR2rMuU4jFvW3pi/sJdRmfMKrrvDHuv4kp+CdiTUZmgc6k3
BwYWbgXksmZ0ivEShU3grsS+GcEDV5BK6pckeRBgeXwNq4YFf3ojdz1lXPkxHdtg7IgZZg0QW9L5
b3hu5SqOOqrwGoxH0hWT++NKhabSB6AVnJN8iC0Yho6dAaq1ibrmOtGA0kpJjZSpIr2H5TRIdWdz
CdBm4FynINFTh2Et4O75YUjIx9Nqd34KMyIH8j/dToQG09CYClm9N1tYtg5tw+7u8LZc2Emuph+d
3l9OBpIq+Xq4q9ptgiGC1q2aEXZUy1bJsGGj4BW1hMzzrbI4iD5VK3mDPZ4senwIX/O4cglzelSt
fr0I1rKpngUyVNYtW8b8wXGP9eb4aWAacJsFTrdYnTer/PdE7+3GPCxGjiXQ2RTx0IlMeFt9fIyR
UuRSZASGS/LWQr/GJ74gCTHgz+gZn8j/VzIkoKF9zVWZWNMBXpye9NyYxs+C9ETDHl1iYtoXef7D
dddwd1/hhNZhWQXJx0m3DTLWWN0yhTY2oSQHscFIwkAy2tNRzvmQKdscf2FMCiLQ9gSZHilL8LEF
o8Gv3+Ye5wOFPEDRuO2Zg6due4IhmmH8Glf6sixqkZf5/okW1xIqPtEKp1wpwuW/D5GH4Y2/bVgL
Cn3Hqpk5AyIjbzKVStpXwyQfmXK7trRuVYAOxdmoDjJ7BuPhWTxQaNQB35xcy5GQeuZcP7KanUFC
9oJQbqiCoRQKgglGfoGqDEDcc+TbUfYZl6RP55kpZVNYhp2yRKia8/wSIzTm10JMWrqFL3VQBn1t
raU2XYkWASNhFXt+thviMzCWiCZEXFlSWIAlFiEUMok8jNYkiYeBga1G1IPd2Smx+YERinW0dfM2
ccU3Avf9R2IC5hAO7XfVoF52JWeKKY8QDLsl63Xs8/5BaNOUxFPBnERIrtgtF2cjah+GqDe0tKr8
5bPfJisa8PHj9znYgNCrwzD1hr0zERe9UMHqkIg+5D6AXF0R1C/hdoOXS9cZ9Tr7JoeLUKhW/SoC
MAph84Jd+YpsLFqFcLuQkGdRlOLOF2YhLse24lanRWUVuklfXiq0zXz+8MSdnSj15TPgmR4aVmS9
HNkgvhHcKiidpEK8gjqq5l5uBvsR2+Kw73pKSu0PALH4zNgERHOMimNSYcxD3N+TXhQdFCAICQyu
+4aMQJLIe/Uk1gbcwDkr3LKmgilInp+mhhbIQx4Wn2ITFILgadDxxf7SLXT7PPFEZa+59r+B59tB
v0KSzTdSWgnzRyMQhTCLQxK6cbI5x+oP53kiISmoEs+2q1Z2jSZ1LHolui2cIqxEG/qW5xTFAKQK
xybqAcJHzij1B9IWryAT0zmpYc4n2JklAHXpUn1CRMLSXzItzZS4XysPGnjnLrnFstBktPTZqQ1t
fcbumIDd33k9X4lCOoC+mT2+nJ1+AyWf/2Sff57Azcfs9eM7t0NwbPQewLXHaGyz5542Vyw9vj8O
FsQhVPKHAPieAW4xYmXKiEuwkPHKTHW+2iFzhLP/dU5jiV7XENWNpqUBAaIf8k8VnFYfrl2JT+gV
i9lOlBv/RKuzI2n/3HAfUXOKLa+pdzW4OD168ot4mjIQrH/dFut4LTendOOHwII35YTGSCzevnrw
yF3m5kWu0Ulu2ZkDZ0JXieDmBWLyzvN3DyqzCjRU6CwougtKQSfc6l1egcRPulSWQclMtfrw2sH9
nBmgizey9cDG+E78K3n0JIwcrfzkAZoZnqKZaWFCWmkyFzqVYG8Hf9j8NoVfhX+tTXxR97P3S0c1
8ablHMvgID0twyuKF4Opl5zcv4IJpd5Ds0gK2qwvBHQdae9gXJ1rVfKtSZQezP0CuUrP40Ioknu6
udyhDS9MVwnI6QKMJZwEybv6bjDGqZM6uFFMnnS9zWDo2ya8C5UxqQ73wVOUNYwK1/1wG0F+fFnc
nHQt2+qXFV41XWb52Bddr8/ZA52h3TRyFGHl7IcjYaq9ReDd+sf6GCR/euNaGRcIqnrDIhXGk4FV
GL4wCe/mxmLA7AWm8dBWYeHX4p3NbpUk/ApnxVkz3XVB2jZQz7nXY4SiRdYhWsyiUniqhR7Oy+R5
K/GQDyXrvGzqU05dPfV4216lA4tBn2n0sPj97eeJu0kC3cyBityOjSkXqgEenNTjJylxciJAqteH
PPfn2IqEVKafXBv2ik9hhHDrFvxDsFBKu+zih11gyi7Rh3PhM3lVbOvJTaYt+OuK+ZSOP8AEwgqK
hxRuRWWZmtQ1eVB3q838dJh/UnFbfgnZeJQDDS84eSAIvaLO4RfMyzV9T1luAPM0x4B//vP0t7HI
iz3CEdLWbjY1j6kciTEWpDughr3VDd5jnjtYHCKJ3Amw1w6WjB4I0VLGmwALuvgFOlyzuc7W39R8
BssyDEasJ5ocn/627Mv2yM7p8nph6o0qEvq3golIVLQJ3i+BZ2MMuB5h5SQyDJAWWkWyNorT/gSM
WJ0jI3C6sLdsBjtZLhKfnacUqH/i/y75jXncVnZs0hbuRR5jRe2drAo1unYI4zaD/PE+mYPxVA2C
FO45XjNMAKvM3tPbaoelaqaqN3+ufzfwFBB5+/AdopVcCEDMPHmGzjWxKzNv1Z3PIF+i9ZGNQF1U
Q2HDH4UWJrvLtWvGCjkn972B1bFMwEKkzaIT8ONMVd5k+zsoR0YQRii3SpFENrTLpfwNL4CnOMhP
1kbRnPkTPGJr760dJEy6O6OW7Rye3qBD86y+sd81hD75gvQSuuBJWL5UgKVINaNSl4AnLrTcX1Qr
kQvLNrzVtIjOfZYQwmpWDG+secSZPi29kzV3DPYVRJg6xkBTnx3/npmUGqVIroe+xTlF64CMLMek
Zy4zrIDzmw3tGmMhqlf0UKebjVgh1AxGAE7AnJ9VAqLAFPovFocYFiu8m4ZG72as4U12wT4UClYM
p1i1nDEv9CNo7XBVb60dVL9HsBkZ6BE+SbG7jG9k7HUF5uSJivhNu9Gm8x6BGmpUl7jMsV5iI5qD
EwcdcYjHHJhhqZw+384oX145ytU1PktecolwK9fnT7TZ62uD53ktYTBugxFnSiXIOy8hG45sl3L5
Pi8U/F1xCYBjBxukw2BW06rwcRX6M/wqLTsKGGat1BZgTx9iVCS4lxIGEUVkfJLfjAuTc2V+UzmI
DlGByiDQwMOjlzX5Z61uJXHVKD1rWRO9UkwlH81aA52aXHhnqzKNOV4EIgXQjZFZMqZn5kvgiiPO
LPwx+0g6sZA2wOqSKmx7bo/oOvcI+mP3GhqFBggju/hjrgS5dQIZ807jXGAbfTw66mXZaLt2+YU5
XtmVsESIqgdC4rRbMT0Zr9p7cCMqiM9ijCQz1ghWFbExeGAgNMmUlceqC8Szf+93euMYUE68Eas2
6DOl5z09y4KsvjOAGt3qvWf7VbRftxd9QeSTCc+g20//nFLnzTUIojeQKonEts5Bzm5oZDsWTCc5
dxIROmMlkD53rh07tgl7MlH/5tzDdNGxCqmagFYPEscXXsHDLlhpitKAqgpzROxGkWblAxt32yr6
1pTfffI2LqdNAeHkpDm8V51tY/DeXTGSrJVuqN+pQh1zM7NS53XzI9MC+K6kFytEXYGbyofAFFQM
xe6sBkgyVnzrzE10PpcNuE51cLH5ZHIezdwqH62NoXFJbyA5V9skJ8x24uZcagFGqS70kTO6HTXj
3Gg7lHo90whoi2pBTd9EeZGh23TOpnsFx9VsxytdZxhtJErI7f6XrrAoKe4ytx2iLbbsIqzubDJ0
QRk16Oxpa1QKu7sZHhft+TwJCxQmJ4PPCvo6ec80yjQv+rqQxTnHiHRIv/Y3z0DMiH5nsly9egpQ
/b7tPVv7ZyBlN92HcjPq9ThBQYDrBNr0oaenwEw2CS+Et3jrz7dG4FDWW7YdeNAzWG8suBtt0MlB
rNI3utVBnYfR5Gce7ASljlYRqnYR9szBjzBNwpOv8/AShNH7/IRNjqEKDtCUy346GSe2BcAwqvIU
BdLCW0/33ru3h4JNDqjLN8tCBf0Bo4IbjnvbC/6XuuCL1cfKWIcLgWLRV+qcSrDY3gPe/6XKOclL
Io8LhznquwF4iAOrjGpdHEPD8gudPrepDJoU4I6mNUTi+7oLoNxgjVpUFCfjIYhxEStkBN0K1Y8M
5BAACpCP6wWrSgtv6+AmofxPNKVooMCwOEAFqnNi3pxzP+uBTcjV683ZugHJv5rWhoOFCW2oqWFo
98NeknOAOO/X1U5tAMNiuylVSIHf0/c237DsP9Dv9v40aLRt8epOfjnFxwGPWh1voG6mZEGw5KPL
Tvo95l+DgqhHAk9v2FsL5pSgnS+vhEXnkxVqIRqO9p8vvJzSKPWm6xSlQ1aTCrLSlP/XHXd1lBHg
WALtZKv16ok+IHPX+TlEqdh25LlDrut8/qyDFQQEQgGai/Dk53dOBy9Y5+QwF0FV0He1n9TiQsj/
cDkGtR+HMquaaMPz94cZGG20r/BPGf7Twz8sTa5Hr0fm9gYQ1QmH91wTh2RdoszwSGbAtLI0l4a1
WTpszr7O9CopkedElyG0JaYk/A6yrETK7EYR+Lg+UivfMtp/OBFuwH+5HPG7JrNsP/609o6lsg7/
jO1ja60gZ/EJOkjEnhD6domi7yWnc/xrljXXjZaByRsZbAHPOm2kkmi7dg4iGYOxO4vwkHD4xK/Z
xFwLtTlVpINGsx6rh7JFd6WJRXjTJDydAbz8Q3GELBxuFJgfAztLhrQNcLwSdl4Di+5ruzowXJ/+
Y2jRfEhstVyGprXe91Pvi70TnXkiAb9DxMO5Sj4py31HWEcuOXb1sOp+MmPnGvR+v/8/GkoPNI/O
PUhAF2GtryXXSRgTfdx5BmKTynLzVKmxf2zjp2xwvky7q7wR6sN3ZmxL3B/wYvvpTJoJx8TJqOxb
pTh05YmZ/r3dFrS5Iq1DnYX5iA/xZu3VFzpfimRitVh2OW4RYxgZIlS+lX1zdF8HBjvsDZWIIgVA
izAWWnn4i7Si5MFhft2Z5AOe0VuMGGyxI+SvajwCJgQQTFj+tmTpMf3WVxAtYpS4Pyg0DLkr13Ap
ZwiZ9LFuYm5waB08+YJlu3eLNnKPZ7iogqLxQJIuwyDIxzAqPaU4Ivo3apIM3HYwIexrDiCEv1Or
ui/D9BvcJSjuVinFXzebqhw65avIxMlI4kmoUUzIqmiGfuxmbnUExTTVNr3P6oczuXaXCzXytank
/M28ToS0N1TpTiJI9DBZd7kb4TCFsQkgGeQesnWCKpbtCYtYE/SXXpsxjZNOtS1S9dj8uFbd6fa9
C8VQc+Qxcn+PKNFbCVkaUoTvaGUllsIvIxkzZBL9PRJFDqJbdwPbJJU0zu3xJN4D5d753MWIgwg1
fDn3XycFEDbglhsPYnyQvJ1Tg7bcM4jXtQbkaJdLRL0nPb7P6Aq4NVionS9Ni94O9azERnS/eXEd
Pp2tgGwOueKD5ZjTANFzDYjQb9x+DXJ1hf8qnP07yW6GW4RICWaGK9BmBZedxfDFVqQD3faYk6Qv
leGAXwQZUFNhegbhM5S2wcx50yvSrNPTHp2/z7umuaJdpCUntuUWOrDZ/x0dwdX5c32xhkV1WKjQ
ViMijtsE4gsVyysf832N878fg2P77syXLPG0wuYRJWvnsDxWeWLPeqBkO124ZCTVOwuxzslLGNGf
lxQNoFFJabhSybu8OWCk7yMgpX+clQOuMUbRUt6xrSyVq3BR1ZgsyHtgFIgYxc6F3DTF57YO1Jum
23LeTCgV6gCHapngzWWVuZbrH7AhgaVSEbZpDsNRhBOAwn3HoD887stlaNK2pDSZE5N3f9LbujS+
e6BCHUEhCWO3FXw3s2IecbvB95IHcJNuCISrTtTak/LAVEnSMrVAJu0N0D4INAPjAs1T2b1nd+iE
e70e7orJRj+RWD6QS3xNsP5q60fX5lAXhdUIexZjaK9lNDQO+xH26vnb2d8ahnUmmv4dtT2b73H1
LhX+8UQktdkZIZgkY7WicK+MUT5CIhYM9uU0iHjYQZlhW3mToYPhJ6pNq/dLa0OJhZ/xf4Fj3PW8
hcn1lv+DhEkX/hJVpRdqYtnuNoMu/Kp2HwARzXEzj+BnbNNEfFmqpb/L3cg/TetKH9nf9g/gcJfU
ftaccbop/+2EC23LFJ2MdqnkxTjsufz5CDRECZv78JaEXp2uxEWgHicJIxGkcpVdGzXRc6zq216C
FVokOsIFC6fJdAJRsZNPmP1p8E8/REdmZmjlfrUiZBuTeUd9LIbwMRWBHQSSfXH5CENsJEpKo9hO
6D3sy2wcd/oCMJGZG5UCHfSBdOfPGBLrXlaK5kr9KSij5HaJYlNlRk8KjNxx0D16t1T9alg7RpSX
/gh2cbdTxXgxhzoWQAsDNkJuKq0v+DSyAnUpMjsK2JQpZo1gAJ5x8hSa8cJG1H1pWCtlwrq8nAZt
ymW+04h3TfqLfFyt63I00rtpGcuKKPo/iQ9f4zs71z923Pt/hPDIWWnpnUIwtpSIXuZxWhrbB0v3
K3gTQIHDYJu5aZdrZwNWfvkzWmDk2K306H/Jbmw7volxthoWu6C21p+4pSuwhNGQggta7gQus+Pr
rFR7pxm4H9RX67NIJclkxLudc3klIfvrXvQtn/brmE9rP23iK86PDgItOoFHVCGu7dEHxpmQsa6y
y4Xpp8aJY4E0lyDZGqzEKe9mZeKTJYvXWWZfP8mkseB6LOw+HaMawpT3jnX45dAm6CQxmXo30LxL
mZwGXh6ju1nmCsFVlTEi1d+u59rckoyQSpc8DJ7DPUjikeLcDhHpqQUPsTdIfhVfVYY78MbFfCzH
7tsFCYyF4BbxZ45uqerJM+GNVAH5UjKzNk/DdxnivPQSwwy6kP/N1+TWbc3welwy6j59sjgGmRuF
xzyMmSzUg2znxAUD3leuZBwcCMRd/EIjurZ6sHbzLHZ1M0UQ21x305jnRikUfCnF2CrexB6AM148
/MKsh6P4w75Vzf9rUBposcr2tp98S+b3Y8UJb76s9okq20eDLJDQcJm8EJZHHTwD93kULkTSkWkt
tLbDaocQ2Obnz3zPb1AFXq3jwM++oxhV7KMaesQrGXU2Z7InULyjSz2iHqH7XDTtCYCINStRIqKs
cD/RlLhoyvnLwVoHcGepxW7N2E7BkhxKIhGPyIYOLysjoQy/rRTGXQI7QtD5rATzk4W+iZVmhot3
BDqtNN2Y1CVydXW1nn77++JOrnVm82JfH4j+LVGuczQM0nHKneKaTPC0pw3DMf04MVzamFYmqbOb
uELI6dXsLJXlIUHoEOjtr453GWdnvbTAR48a15seoTSVuD585T9+GwSOFSYbadIeYz7nDuYN6JUS
e6YYUflc//RfiQKo9wlOeJsT5pI7ADg2gc1bPak0/IQ2DvNOca7n6kNxPcwhpBJosf4+ndRWmpyB
lOB3qqTFQFoaLrLPGYlueIP1Tmg5bUwOr/+udwSfCAI5Wpkhix7g4NdxUegEUU5hZoE/6fL7uL5K
LoWmvpx+Y+9QAy/pktFg6m3oHi4+onwFfKEU0SpkvRzgleLQLCSlH4HvFJJIf6gp3GUASNQdR8E8
bmvLyGy9ek9d+efW2Ptvurc+iFyYwPF2sh/d2Caq6yqaFTtnZGNNMj3K51Zaw6h/8EV+44tLNjy2
jexl1zQ68/mgqEBm5gxuDp5Ys8TTLJG4Q/Y3cd9xvEjMpEyNpBnLwXE3rcoZlihn/rjvloIwjahg
CxTYwgOS1+xtl2wZhtvYAuqpTsyElrRsqw2G0OdQIZtBuy0gWk3nM5KvQmmAH7Vd47SMC4oUhutU
N8Dvvv1NlxE6UUMQkxNCW6rxTRvu99QeHCvzfYHwbKP2mg/utQHAwVBX8OtnqmSc3dwZKqJz5rSS
vpI14Y1Wr2xw+OhPwfK6Swv5K0XrDsERmQPqezjEbfyfsFE1Ym2i/sYh2FFrIKCea+rYCSfWsPh6
TAQJdTQSZiSp/uH4i2OWAq+wi8FlNpwFnWe62TCFtJJhg1VTdgbmaxhlubNXRrZ8xD3ZcQPl0T/j
5z+GRW/19RzeTBWGcYSAzLc1afE11Me4MjWCi3S5idmEv9BQ7yoaj+3igzh4n4aB6+0hNcB1KLbX
rBk95OUKfM8NTkhQy3kCSMIW8EOLLytwjGNiyZt/mupdBgyVuJPZ7rCLX6XCamRdTXIkEutJQJYi
IO3vHlmUpbI1+5nBbMMd4vHaT/Dc0tC8ciAddOEdOkzEV7zu1AoyQ4m+m7XkWAPyBJY1oo8md/La
EAFpCG53lpNXZQKW04bD657gQwP2sQaXkap2qut5BSZ72/q8IEq28QEyqooj8zIy80eF3V+aF7Ff
CHlXvBkSJYWRm7FQDYS0x81M0HB/xPLKlJZp7aHy2F5CGOn5JNFKxQaOG8p0bwVFMMsjAQDsluuD
djkSlp38GgRY1OvSjDY0Rfnn+Q2JynZTG3LUoXtQPFWivEYiGgnDrC6CzRH2pwqTR+4FSsT2G8bu
GFjNVy3V53WSiCBplV52ssuLnYOMx1bRaeDvCxIcrPTZUxHEh+QAoyHjf3k/XZMm8tenGw9G6VVI
zixMBbfhyCpYdP9np1c4YXZS9Xg/K9YAtdKmywqLaPDgOfI1dtQ5s8/gtoWfYTBw0N0xYPM8CFs0
dF9I1nCp9HqBQmb84+rdx6LOAY00JJQXUwAoo5Whuicc+HebzTburFUbGWrLhxkPqN86AXluFsLu
fRyZ9Xo0N6BPF+LEmgQ6WQMx5p6X/g46mNpLH62Tag7EGzfNrUHmIsotnt8aUSDhvPgHns8y66CR
8REnLf4HO9JJdqqgDhXINL7kuHK5xogTavCosIvi0fn6ayatSPd/SVqQikDwatSTf0EDXQKbOQcI
EEW4+ZZS/WGmqumqvY3FqU9uja4v44C5Iv4ncWB91yVnrLSIEA1FOrVZOShBi8Oii2mVVGKx44eX
SsRp1g9jbRptl0a8T/n23XVei9nwgLnuOJysnOYVyUGz+B00wKvg0Pjv1skhxyC9CrzwPHTtZ4i2
ebyoCtudk8hYYj7yPo8uRlf3nCYE4F+lPY0Ft6K9cN+Y0Rx6araxTopzhVKcD3r5WaDnm2dEwiFs
fOWNfccYY9SoLoAvBdB7jF8dLgntUqM79jixBEN/31db5Dv4lEMRfgAW4FCedkO8taHrlJ0+G4xn
876qvYpjmZIiBrN5mDT/vi6N7pIkzPmk2yA02jIeP0r3/fwU+hy/jL8ni9HqPtD6QWF3Iz+HAntn
B1cfFpLfjIPtp8t8OiqRrs/gXz2yjI0be7D8CblCRbUX/3fiCX1AxCazop/ivvY8xMJ3+g4BroYO
a2epfmFQdJ9zSgl5JHoqVsVSllqEApEolOEL0s21I5+CBcdOr4qWb0S1bMFoaXkzmszTtCW1pMnt
VTlhPNzDBiZkBmJUlWmWX2Dz9i0p0QUzsZSRbap3LUivCSUWx3xDcq9zrlT07UxsASkuT2nxFgUX
AYAlYJfOsEMQOTrKt8DLTHLtSYPiKi2xKmymH8rNNvAUU8he+t/szQe08A4F4NQoXG6KFKHRn7oq
OkS1CauVv6yjZA4ZswIpKc9xIz0deLR60SuQRnkUISIIalLQrpaTEIfPmsMiniduvIE6xn5iUYwC
i7pbaSzhUbbNN+Ki/KevjwBCXRkQjT7rj6ojRm8iNinmE7EsYbr+alCtg+Sz1tUc5Al4LFyzb0uX
VA3wgY+hdcgoteRkJ64mEHb5SE+Wyo4u+od0GD+6oMjpZ2r7ruuk3sTDIC2sGpJELmzBXW/upww/
/EurN/FuMsoZHaJoICtiiICqnYHnGHRK5lIhtESvXCQ0gVZJ2Z9uPuaLm6tkqMAeGQoVIuCojgJQ
rfd724UUfD0lPIoYihOxqxt7XIUaF8LECVMczf5U6kROsLWNY0l7ILnJxIYmwVIpHDjjXvPhSGND
jtJ82Bz8P5cbVU/EPoxmxoZD5Zpy/kqS0RBuHDHibxEkGVe/rbHcr1jV2XaA3K2YzBcNW/UNrqhL
VGGESBSBKAvPGcM/5eWre+m7Xnl1NkrZpEW/K2eekGq7utRDG7ZlAUO2Bst70N2yU4FjxEHZwy/l
yN9B1/WcuXI1DaUFWcE3YqkSUegFiyX1PH54+NTwlHyok7JxgZxycbkBLGvi3I6dcda02gophFXZ
Nyybu79EK8/NfDvToxoADogeAjTVsxwsDcurb/d8XdyG2l0fGbXv/6vza4CB687xx56EYFNBjppz
Vlg8Eb6ELVCBVENWHuhJ2HtbZEW8dSEAxVwAO1PT/O66JpPwFoCMl+kxXf1pX1Nkq/P/sLSpWan4
Hy2s+VkY3+6S61q62Pch1SHvnqnupUeUyAaoCNxnA6gVaFF1XuoB8lDWGurQRkrdnRc3pdSA8lJ9
Rgk1g2cg2yrnGVOz7bmo0qJHHBJN8KkorAnjASj+wNG0o8ICOTULTj0aEhpJejfYdDYpnkhVuybU
tAnMda3CVrmWNbtvDXvdgwZrU6+fSRBJrJgI7/UqGN9BIxAMnTbB6FuytdCgWxkpUtF5W7cgdYxd
9Nub1eyTZ0MpCtuOXabK6BXscJ1F5HookJ0+7wMVK0wn18wrQFJas6vW4DycRo7blaezR5xLC9nC
n1nZWNh0sA5wFRctTKDE/7U0ejUVL4cKoTuaQN3vYoPrsQk1KDr4pwHRQPIutDGQT0LB5k4nYt+k
KTkpvYBqMcWO0C4/TTRJr+QP5KOr9/NflFnpbjlQgR76fYRb2C+MvVBF5qlb2wWLa5ldxtu++dsd
MuW5dsWtIiZXJQiCKb/4GpwOx3nm69mFTrbE4GlzQyRVOiTVeYc4TIB7KtNXFlDSfEqJkZwe43k1
lL+xjNPFIjYuEI+yQ2zyjCaRkg9IanZbhoThjmGqDrJ1QJ8BFTWbYNDU2kQiImzv1MgmYdsuGyFp
r05L4W30cp2jDK6hZk/uPh4V7MiBRMpENdzggKOF6EDHLi47FY8TNfkhw8MFwdpKbzdVBtLw4OVa
bXtbsgucxYZ3Rntb4Ni5eucqHR4TP7/nBMNbj5p4goTeLnvk0DQViu9UI8PKHVeO08lR6OhdlYS1
URLYlgl0wbyjZPznG7QTGWFi8Ipp8KmqzLH3FA98/QOLUf1MmJZRz8LkOyjcETuinyRmnPQe70nt
bbrrlDKWuVt7hNP5NIz7eKI0BmOP2djwdnFsavdbfQ31+DPMN4brDN6+F02KcTLMQZeDH7fedOw3
Ati6nlk6o1GG4KTx3QaBdQPqvAeWpwE/Zqb/YrHTuroDLED81D+OajQ898sD+HxfGgP6gy5UCOQp
ViXAWFRFyJwxE8pCLUz7l9kHe+Qv4FzTM4IMUm8jpQ2HAKfdTRz6ESqu7d7x4G6EQeiQp+TQbgi5
IulZRxhS723CQH9JCawUck/CvSKRBu5sXrnE2IUQY16hUQ3MI3wlTEpGDwUWhQb9r19daP/y8anT
Xtd/UHzmTbE9g+bR3CFc5KJR0EtvDM7hJ6oDUtTe3hLOHN6z6UaDU4oCABnp5LBJNnEyJRc22s1R
GyebZtc/1qUHmNfDp9cFNdNrn504kJ7IU+b5kTr6W99Xv3awBWGRbV/ZPaHkv5MKbYJTbVDtLbJD
wWP0lEgsAyKv37fd2YM4iNqTg7aZOwtfeoN/4KzWKL5WFYIgtC/YjRLQLQetMVRLuJbnO+GCRaSX
dQDDzFQHpFUvq9k6TnNRdJnhBykE2vBweb00bjvWoktQ6YeAd02/ExYeIqV/5r7OehD5OzAXaj1P
pPf7bMlKEelBgjFjhRHDdjU8e30gCRsOj34TDs2nnulyL2C7GFmutmgoX7A6Z5ERF9D+6/n5Uqcu
w5NyCFDQFTq4WWK477hAo4m2ENCWmycR0HxgG3nizArdo4rYK7RBafmLgne+EwKKnrDTYYyLLeyW
Wg/ixbZ5x0pfOytcVhtFz/mXPY8oEALgP+zuci/sOyXijPBiun2O9VmP/MFfqfbUMoStfJxYYKvA
Ryg1m+2BAxtFyYQ92/Xg55GVRbVJ9MWZXlZAYYNDXxfHTk+/f3kvPdQj45J+VpWx6Z6xlgh4Hrwo
y0YG2Fu7jo48sKfQQxAlowoBe7lKIrB5JEpJWFxq3ZCj0LrPvvadwLdTei58oMRFxq9/ZEdb+eNQ
lUHRFVrsOKROcKnK41X7pbifaLPkPtxc6Vr5+2htGvNdblhznmePYAFmIv8LHWnzTubISY5E8nqm
PqxWDpH5zC8vHwzCvSAc2wvb2cPEOBL0hT4Gvqbg8oSIsvKlIlR92pVjGWy/atRI1GikYytQ4CJO
g1phA1axu5B87f/jwMTTxYa8Qcw7QmWcsu97XLr4ThNVlijdF3J1AjVFYFkpvOnbzlu2TqNqLDpP
XGftefYqxqOpM+Adt0FY0ZKWAwWoOJzmgYtia7Qi5FHD3j0pZ5Wz43iKnK0zAaJJAYDk7EezGUe+
AsT8MR8v34u2kBGkg4UWDC/Ms99I2Dr343O0iSMTd8G/aQzw4kJCcFLmTEwiQOV5gErwKeochtCB
IzPuwIBwjphcz8RcqlbVScHLxHU2s9/CGk9hhfBM6o+B6DTRmC0fw3atofkLdiPBViDByBK3ys7R
arHEupgl1rj3wa+gyon6XnkDMR+705Xy9lGdjeKSiXiul0JBMguSW0YO1YeJaYNPn7TFfzv3QbBA
Fzwcg/wMY8UAd+c6Q9pNs/cMuRzY9Jrje9chlM+zHOPIn0H998KbaoLWEc14J4369rQt+vHFt+fE
6Ujm2pXWAmXuroHEn/cAeISdADYJPc8gAAQjBHZ9g1PjjJJfbEEHGZHLNw4cjYNo/Z7o8Kam8TH/
l6VXA1+5TmyxoM4Ra0VNuLEL5N1sIRJ9W2FcAxDKFWP0AJZkiiJ6bQ/pZi3gbTPMKe1d7aZu1sEC
FI+tvyJmeRDnSVZ/qJlsdOL1auMx3nwsVvcULEFN/fzPfXdD9Er/5/W+Mb0H/pJvlvnbTLd0M2mq
Z2vxlB8ay9UDFIuYIQoZ8IxEx7re1sc3TKlgffvr5x1FYVA9Nq4HFkC0NrcTceYDlQ/Pf/TvPgt2
DUl221T3ELM8FWQKXMmFRB22YXZmjqeRjvOHX9nY4ybHok9NKawqCBGGA9CWgqBvDrHFn71NaU+5
4FoQ9cKFBCK0eMOZaP85wNiI27e8QtHQq4DlCS0qZIy4dsFtDKT0CGd4s5XjMJ8I31m7bQt1MZc7
Xct2T/LQLeDc5QDNPpQKcVXmDW6olNSMu1P7XG7Xt0/hIc22HSziXj//V/ccfwRFSpHDWLYbteNs
ch+n+d30/XhnStXD8QS9OBXosOBQ6NyvKxZABtuPFjqLHeYRvgvI2m8LfB2/2hMQcACx6NSD4qzN
ErSYhlm8y2fMeqFHQgVPI5dk8vDjkQX4atfLJ6X+jkWu3FETkfjq5Vzh7TtjsrtCpL6lrXo2yGSo
hgGQgTP4+HWoshi5ndp2rA+dDhDTLx+9PFSGFdbPPY+fNhu9quBybG78URvHuPQBSjgXrH0KxrkT
fHgfFIZ69ZEDKjm09vAFpwefbS0CPDmLD7aAbYkAMA5G8ub11KqOAKc2piBwxwaaVmlYZpwY+Mga
V22FLy/hwDDRYf5tK6/5Nr1SmBipMLd5mV9l91i7IW6LxuyzKvzsw7SUGt4ZTQj66STSl42DvJOx
2rrJaBhuGHCQuBbYwrywJR4zDijZqmFX9lBtxhHEIRR6A/dOjUqDeKvS4ZpeBjWtaivhhcOC9Ros
28Ay6MbZujSeDpcuk+AoWT4dKS6pwOlu9X/5Z+ytUAm1OsHbjwe/s2D8Fdo2hvfQ9z04mfZe6vFR
gMWeMAmHUuW351mu1rCoWurajkMRzy25sI0EoPghct6xvaNlLaJhhiUTO2aipk/ChQ03rhI8gxmm
4u/HsUtkOvTRG7oVhYoNNsjWsStFd12P1A3kr/GmxoXn26mWDfFUsmsmpziKpdTb+9LGoQERW6Bu
sjMuJw4BYg/Pe1IDzOKT/Imuuc5vcYGxNzfNfplWwrYD8CxvosvIph6z1nKzIuHDlmKiJNspjK87
R06UWRjWcyMCsNCFBu+JoLmhc/6K0nLbs27o5K9AeR3ZyeKzDrEUtCndPwNtnQoJTgqyDS+DEqKK
7/gfwH2z+a7cf02HS0/tZ0K3HTkanhuc4H7MB4Ep7r3LmJsVZ6cx06VnTGj8hhH4IwtBXNEZl96x
4D7jrT5Dx32HJsSyiEBTkBJb2dLVWEXKL83vaXTzGdOsTkblXbhLMcTngnW38ZjXU5sbYxnjDKIG
rXKLhOVlpIhqX5txLmYcALo68Csxb4GeVs7qaFKbX+UJwE9i+EF5XROp5uhmCEPogN68FHfY830g
6JQyLRqAc7ukMgU3eFMqzMU4M+CCUuewcuehkADymHm/SoGX+Dak4xTJZdvtGJnUT3PtJ2/FfaBj
nDRybyBwXx9QxMnrX36dyB9oJb0ijQu77nE08S5zPeETC47DCcUbV+D4RoeVYfLyVv8P0JH2d5Q4
1xv40tqo7sCs4GPn8mF3HnmE0Yl1Gv+PWauXE9Cjykk/ylrpZrAxECz2FlpJdl+M7Jbwp1DVOmbk
7uwza48n8UsftoAs1lQPqKk6ALAlQsaf3bT0Aa6LnxrK+EEtnDMVvCC8VgHGNLNyHfZi/FjsTDkn
A0P+oxejz+DhsY28djOtcF22gLM9FONl3XJ4g1FPEwAc1T5KWBbXRNMfFx0+Xj3uMN+zFJP9X/EF
nc1LLygwfgro6hC4R679YUla2yhORMOL3DxdA22CH6XAgMAlm26BRDx2CFh7LoiAdp9ie3bdE8Ws
XyMHJF0p6xHtQWT7qJY1OJ669kw/0UpY+x0g/SL61gZX/A9fPHZqWPZxASXFCAe8zU47jeRJY+pq
JWaPAexs+TfBlVN9VwJCKvseJ4uhY7Fg79AwK5ZFf9lu68mgr3FbGnPAOYvby9I/mCd5Ow8Qf1ZE
lM47KrQBuD6hPkxq1aQaG84G4UZLfwCCGrA8cDRja4irAxqnDPCWAzVIaM+aahQ51j+DuwDMnR9P
PMAcdMxXnwwKb+eYFPU/9F9vvzPz/yGEQceU65hK4vLtz9LPKcLWTybbpbX3ntFD8+IEOgtEXY1A
laLDjLIeQwnKL+5WdSPduUvuysJnrxbW4x0KXvbCsrRQTHI6riLMx+h523ordZyMC8DawIg4H2uo
2MXAsCc0pL8nJuvnUXJQNE+VJcgIh6U9qAazH2Rqd9SUhL39kTL8ce1s2GidC3JibNnTSz2Jr0JG
e2be6kD23h8950atgMEIrv2N0NjoorU/NkDIrGwXpDT/+2vjQyLbKBPkkyRCaXxThvKJQAgdpDKw
xDRtOS/l3KP25yCEYpCEO46gdLbAcv+5Zy0JuvrNN7weVdIHhVseq0DWWoUIT4/pJtzYzU57SDp1
BQUWG+/B2Cj75zlBT6RK2Gq9oI2s0BcWkysWtV+vPx1hwJQ5HXuRQstVvzPlM9WjNpEyatWfMd83
zPwgwGU1bv4gfRtKb7eaZZazGf4W6LyEW4IDfiT9h3WaEZq+/ZjzaVJk1eVh1WaeesUXCDAPjToV
pr0v5aeWAp0zOJVbAIZFkwIBJ9U6ziWlfCzgMZ3bASUnA7KubMuobSH+k1cr/PysEoHRDnUatLlf
7N6662EMN+LiZirIEhI3FZ1yaQxD4HMEhohKUKMeM2MUq3BmvhwwH9pt4VB37WO8SyjgdFiZhBWk
tlpC4r3w4XCAhQYe0AWBYJ6zJ/zOQhx1U86BT4DpMM/I/xCE8YWKPFZm8jQ3WMORpDJeRDdmKcUF
dnceePgb1sH29sgi/nSge2/jxv2MQTMddjfwZB06SZSLj2AYiB2eCyap7TX/WoisvjymMdqKR8rg
+ztMCC59F2kz3ArNtLBfgZEWYsW9nQVjzT4AkdL7HnoU5gNq4w2p9Ma+wuQgKiZ9mR49x+LjLrP2
haX4hKAfHLVZMxfnzXZX5P79qYKjL1zBSAx51Iv9lnN7oH8SwXgqeq2+fjHMZDmsgjtKxUgaYKz+
aPs4CIgWm3A7nKrKWMTUB3phL4VaPSWOs4w9Vknxgt3OzuMYCoeeD05FwmUxKvJTgN1r4AXIGD1I
ZMbzcMP9F0X6jc20Ym4eQ8Z0BPfden5SSlGnTWi/5lNu8iOBtGuH0rghJnJcBu10h3Db81ollqLo
r8M2SR3xvytpN8cVcCtlKzLvZVQp6DYHIT5VFyXLBH82TK7O/YnqdAv0hECKzxPbTmAISvJ9uBOt
JeUSwaeo/KHWeHyOT4lu/IM6+kUAsKUFVSARuDcmqEIZHmzP2dEOwSCtwsemGXzmuE03A0aP9bno
9ylbMiTmHdWQo4p6MY48ikgfjhkYUMog3dhHVgWMphDpcrfEvDEtBnHEsiNHtef4G0tzxl8fXa87
jAWG+BVGrMog6dAhdVLkyYjcavN/DWyz+F4fxTrAwLShgG0/G6yuKX5J5WkFB/+KTvz/DzdqNAKM
rbokJmMxFjTFJYMQ17DBspGiERbeXtKau+Jl9CJ7yuO9RCCpvEf9Qnhauyh5+xLr2Fwf0AmYLVDZ
euR4z4cSiq8yDLo1pxLP/Sg9zdCQDYJYlFzAQpd3DZZJ+Y7WpfraviqluxL15pfE1AwSlSQzuDTs
qRKCcRsFzgfUU/X2ar8bTdBY2ScVcs9EJvYtYAbNIIHPE7tOKJHSbiJ19vRCN2Z76fP49LuSGlkl
MSV0sF1hNkDg3F97sDfmABIXs1sGbTDA8N0Vt+nWims+DvBqPZbJLlco9BiitsE3YFcGPo5UuKoE
MguAMHPVIxbYTNQ1VmOW4kPiSgn3Bgu8jCSuNvUxemrgk1NS4URFWTyiyNS7/eRzOOMqdbWHh30l
1i9XOJaCAg3l0oP/Glk9XCmFFWf4wZqlV7fX8hrpIw6+9+5kIGbwI0peBN4EuI9QgIyHhb4amICy
EHoHfqsYiTDzMJlWDA+pHu+5E7shzagMoy0kERyrS7NQ76UtN7+UGfnvrmXibMkONXoIqGMji5aE
wv8ExO1EiLOottUCkB1OLClDHokQvldoOT/dAOydVjHZMz+HculpX1FONhKTZk2k2qwA3UXnk4WK
bZqoWnA++B38IB0MPhWqyxb6Db93TnqC/gwcEQm+qMNgxJvH8MSu74zFCgyQqZSNx0BY1F/df3zk
1eae/FXDqCT16DEqE7Ze/k8laFma3f0wj51FY3obTjZE71hSn7daIswSjXzA98mKGs67EA7nWiO+
crPjpTTEaBAZjfv70AX3rV34DhzWVK7lTB8GWMrT7XjWc5tUsV2gRWC6T0cebSBgb6P2IKmA1pEp
b0Fus9WaB30XaU3CEuVoJ5sMavpIFL1Y6Za+0vuE2cv9deHJSVFES1dh2MYDpY1NJQ24FuSVUikW
kjBZHiX9PYmg0NIU3ou1js5JIX5zT4ig/68PQ6Q+9LhFocyIVYJdB+fwA2Zbczl6aVFs0q85uAwm
KcYNZUjA4zfTkaHoV3ZP/K4fKLO8yYUIDCQrpgUY9Z2Ij6XYrv5c71bdIokG++nFPSvqzEl/4Zfi
7AKmio5Wd4OuCO+dPXVZXgbvPojI7SxKmkuLpBGFflC9HL7iMcT/ZP8PnqhOwSLkkp7BNIPeyil1
MJza9GBjJ5cSgcUg74/Ej6wTIqj/Mn6cqFi/1Iy5g40TGnNfLzEe9NLmxgM2wQWEzDULXFjN7tSY
tHg4hxUNdYYFVkcFFKtf64wY7v+QRol4t1TGDYVC4KOc6TnF7YQUXzM1Gb4YtMDb8TkynYH0tmVd
lWxP4d0p9z+VNyh/WhpPpzntzATNpsagEAvSr6FJ9vC28Whq4WulVADznSSbZuc3QmP3mBlcmdaq
9MA9cW/O2OCm7sM9jxHYF80PkqSBMVQqJF1j7dIIMnT5e9GzG/J/SA/X2ceTiS8U0LlMcHaAdu/w
FXqnnKbSM831griwvVnHhDqlT3xft+MlvkgD8AZNY89IDMEmsEIMN0kje+cPZjTFTlpYhge53tLZ
67jjbWyg3a+AaVN2ZZ46re1Vl+Pww3EjRYZk+Kjp/u8ken6rkK51/6gPJepQZl/W1kO2fmLYpVRT
rDUahHRmBqkDVDehgpkLM3Fs6lbqzEYC5wYv2vMNgNdWgLqS5c7lYCO4geq0xonmWK4OSW500Ggz
Qb6a/OZi0Bp8DAjCKaZAoG4o5oqfgZUEPg8SS8uOBJPwiu/uPYKWUvadY3gplJUGt/zHLyFURrUM
iki247+pfQuM441AL6H6gQj4TdVkb46/Q63SarfNlodjYXNelay8OYfXV+GvJxSLx1KsMlLN4M23
sMh24PEaoE6ubBSsaycTgah599OPhG8bg+9uSLdHw3YDG6FI7WdkpuU06PD6brL9go/Khi9BmciL
rgNxJNIZEHL479Cl1jyJ+0pzIrcMKMA3/RJeNbu/S2itQVgPCPJA//yex6zTZZh8r3KEbin42MC/
IeSRBXsrtLMTpEg35Hdcovk9QtgwRsvMiq1qqcR1BLLuxocaIUKF2PVnZXqOCaGVxq7ZKI5qGaVd
liPtKAcCa6KWtGirVgvoRUY4LL9p04UdkPZVUw8izDu4SVDtDCaVWrzUhdicAKasTnj8KAcZ10dw
AtOdFT/+GfNciSCAbDHEOkyeP0DPOjrMF1Fa2CNYdnkIA/iPAjqJZ6VGq8XmWrrRUa6DGw4d12Xl
yY+An858yc9V9L12Kkr17zHlNy9uxnTghoMSmhjcPekdxL1zw4oTW9yF/heJXSm+CHx+XNSdkMPG
8diM3pNDS87X2Ji1vHdnHxe+6cU2Wp+olRInUSLanLyr6XC+jcsIITu2R7T2BUrwUDUR/Ragrf6I
92pDyRFWQY1Q+Q2KBlJEJY3OY31zHPj+8yj8o5ZhuE4fiEElUp8kIB0Ussm9CLpXbJ2wrPMFbbHG
MWrLmK1cuUWNNPnx+TBFSlomYQCSaR2HWWvGLt+ajdvBWbpU0SuN5sZZKyDOWnHfIvRHGwbt5NN7
1y6h+XiRoVp3xN0E4QKASM4oPLj1VPQIxx+J7W16X4PZlBOudjBYgvguBvIFP90/C+39FLNFFymL
dVv4uY0xbpVd2DXo4c31CNCsu3ERSIVVM52otL+xNIBuPofdtzELSYTLlmga6LbumLf86j3nlLDY
X6mWx5gQg7Xx3dQCuP1K1zd/KOmDBDGniX4sk4Rxi9qNyIBiPjIhOz0jJNK06GhxH7d29N83UR0w
x61808kwV8lJ2PSHuOh1xojUyumheHDUaGIJ6jTNIeSR7spnJ2YGi3N6793ieAoKrYcj4D3gQJe6
qLeIhA66tX1DPJ6nbS+DWYsGCF10RELghIib6kirrgvLayUKMPkjDdfHpFVUobxUPWpHvtPeddVH
/V15LwWquzCjGKklCTOsOluEgS6gaVW/d++9i6YxIq5PA3fbmQ6auUz9uGFrzb4AM6wWiFTDXrEH
hAghUrqI087y+hdX+hv69NxNp7HrvblwhT60JcREWpEgfNtqrP+FHKvrIv7SCukYqTd9pn+mWu1Q
kE7IJfunml+IDJn9z9pHSdFd6Kp8N2zFqXzgloif+tfEqmQjd7h53HEs6v/2GieQR3bif/4uMBJ4
6c1W7rizXqsci48J3rvSxyvUaXag67XwYMymMEU2n4sM2HKuLuEQjj+IwrT7H9Jyveto4efrIESM
7BCrFaFtrx4x5BY9j9Gkj8iDrj0zUXUtRWnlXgruIc+i7I0NkGWH5K06XcJm8Yfe8AwWFul1UMZw
rBu55PMhHbAXk2yECtlJ0h+5mw/EW3PyMylg54VS3CZL1F3uHdFy3SlTIn1dw3YUrW9CM/YSDZsQ
xA3elcVUN5Ir+HfyzF18LpkDI2idZ1roZHMxwgTSLBiiZjvpf3g8schpGNzr1ZtTMnrVQ08o35ow
+QMGJPXAWg3pKfH8r/uwQMCkj1fZIMP3NehvprQsPDHcqat5g1hPmHN/2eVZj+ETj16IW7ekFArA
CKUBZZOqAf9OQcj4LX1G57D+X6jFW6604CySMYCoUzHTP9NmqflLP1NRB+S9XuRvD79rYWq7VJXR
3crQkfm1S3fm64yMjjw2BDSGw77TA2CpfyG5uf0okXkh/4uTfCBxKd7MQCLTEqYVYdQsKDjTyZ0T
cq2IcXtZ5v6VLIoNsUhFkKppKtYa24TEBm0Z1omWr1IWjsJgkZN66FEJHyOMjyg6no6BY9wTPknY
qR+qcekQng6zmBhxdGq2XIa6j42i5WwbG00doHSuixTGgR8uEmaxLTPt6mnzjP1osfH8mIvOtwfa
mLAtNT/6Vfivn1sEATYT0SrjjRLaj5b2vuv5LQIDlv7k6JAqMzckY1jReA6xjjkBNRApe3mWitbz
hdm1/YqCI0OWSFNqMVx49ag0raNPrEr8EK+E8P77BhtGlbLSWI3O0+elLTtyDfAKUHOPwU3ryyPE
tSl1nZR3kC7dugv6VVmCSoHvEbgR+BuNagY+hq/HvVQzVwrirVr/d+S4k+zoCxP7Y15XOEQapjiG
VIa40iXekGOly/ip9UIxI+SRaiB+c7txYBwAXNXcDZBpO9u5tPm2TfaJzBCf03pxQFLQ5IZoQj1D
0p6tEBHKbGBLCMNOSxS0xds0LSNiyVElkMNeE7DSdK8jnYGCs9dk4lLQE34REboGj8t8bjyidt6R
1nhoHgMz//8FzQ1zhHueF2NNiYfZj7HtqobEM2AjHZJ6jnYBBItz7x4WQmET3YHkQxhlm0Uub8mQ
xLUvYSbhngCQRBkp0xyOB8TmzNkVmlKEQNWc3C2jXdDt9r2WpS2rvmDYfUSHsp64vuzYHVy3E9eW
vSHkcgcXVoLvoeHKkDBCmdhDqZpj5Oayi3B9NlJ6cLShnJoMgMpIYC8W82WuaFlkc6wKQOG8nMEy
7FwjeWg0cGIgiUNdlyNNxkJK+sfYY/PhbLx9ZNc3hEbOW1o3lk7kCwSR38+ajmYtZXcidkXU5r0s
enkfTsWEy3poK/WtCA3tcPNPGKZXXw4D3MmNMmHc6A6hpQ+eAP0T5TmEESQuzOrBf2wPAB206dvG
UhzPvRBUzDxgdQg9WHjI/HhJn2D4BcIVPjE97aVWvFHMBk1xlWz07DBC+HsJRyAgXrzQ9emLxHG3
5L7jzIG452gUgsBdmrvWH+4g+Mv6voJYtI13LnihmCJ6efCOnUyMT2MzFgdGACcvH0oWDTwhwFcB
DTatVarbP52yJq3/cz+6hPcUVw/YxIQ7DVfX7rCxuJbeGBIfmteWypY5swBhIO8eikTxpHqRXcjy
WCf++bGs/Ng1MQK1XQUnxjb6xbWBhCsLEMIzji50WPky+OV7a8ltKk3vZO/PqK218MV6SlbtoOe/
u4pGn7yTUjlfsoQyBTCYMkeGcrJ3GdFkYOnP8fXdfFexmge/vdUJVUD0TkqdIhrCbnU6I2qPz5Xx
Tdfyxar0XaOHLPKdAg9dqif4KnPUG6CvfjLwc4gaC6R/kp4H46NUzXFmmVUrUCRd9mqYfrL4gzge
3RNhosEXaqV674koBgcEPqntufu0Feb7yo3gESTsnjmKMaUyZVFgNzxRO9+SZuXQomDSfWGIB2s+
RByuTx7KKEc4pHTax37SCBjr2OwT8H2fJY64W+GG9TQwrqEKDrZ4rFEfuiL1ti7Sa98NDic4aNYf
kP5Ns8jEQAff0yP06oAnVM4EMho5s1btHgkl7WbsbcPPvLjEwEysmijKIiZatVaLAtj0ji+trfJj
1IOkqlVz6pE/vRZOGI/kAgypIPn8Hrg00l3QYaC6QO5JmDnZ/8KOefOjjrnCnEKDpmtApQe+VPJV
Bla5ZTBKeeQHjLsIlJ6D/aYZ27HrnfN1cwqvHD7xUC4uBF71vUEmwOaY0IxbueIsCs/BNja8M3Ow
5AqvDM3GCyiQPi4rC7wJAYxqao/nhAECNqomqqGjTshNaaYvkRYxXALH4cPXsUOUUiP7UhnPQbYW
nNJr7EcwVCggMjsLb2KEELBzCnvqkYorXfCDyCB/Cqlz9yfwnt5wlT2XdfPZlS81rlK6tkcGQg4j
DLJ38g/Z4kBJ1CR7p2/l7p110HJUfQDJPnALt2bFwbjAm6n9Ytd3Qc0bSu+yv2GTeGwR6NilNkB8
evV3dMasjsCmjEdG/R2r3sZdOdSk18M/pc/AXs9pyGY3SAwrO5NG3RoxC5b+TGVKsc8skvYQpIkv
jBBNWBMJTSQxW5XVzPrNjKmJOyCWx8vGdY/3xoQiSMfGFobQrpJK7lFILnh9S5on5YD6WyRpO3rN
vhmHJC8MtWOIrkBeUpss32rqr3NTXJRuNY4iDH7LhMdPug/d/xHZro6eNb4uzqDixIvhkhQmo+/h
4wNFG7HuIdbBluuUcC7KVf5YWgPN1jq017CpbSOPB2SnqE8LJIn06pMJB28l2TJGOXGb3QqAhiDu
XOI5HUxQoqUQToItnPCqPQmHmYY4FsRgS2FT1tZqWKvmrhzmv7aeb7JTxaqZvOLDUTYJzs4oz3KV
tSmHKl6AGbhQK3T9RYqpUXo5PPHQILL2rTsM4d2CTwnQbKDdOu9cqmvXTzBpJfzbRH7txxIuOeba
uOO11eAB1Oz1H/ZJni4X8OSdIhAwTt2z8xT5TuLHok+BChyYmTAe9aQuhXI76KuvLdA26h079/2A
SmNiIgtDNpehiN/H8Wc6H5DvYYxT2HXPIsID90UWD7O1gxvM5aD0JbTBqEXw6o905PsSeFMpatN0
SpTCH4Yom/LY2Mmb6061TcKbxHJJv1m8EjSdDv+WV98CozD8l03aqMFGYZ9DMtayHwfNj1Wzm6no
8F4+vA11xhrBLLW5aXfc3gO7yKJ/7aFBNN4/3w207fYKazJStCEjLEG232LTfowIBadHu9L1e4sW
fcpSW4UBODhYJPlZwx3IuQnJqPwDL0Qdr5o7WJys0Lphvsducp/sCM3ISeGo/g0BNbyGF+bV04TB
Pe6jEGBSJ/jkTtOnPvChGeh2K4TGrwDs+qltsOpZ19IinLhS1ufdVH//Z/ZnyxJ/BjcQ9DOPm5FV
4rzZMSyAffNBbwkc6iwKVO5SQhMxDcTZwfZSCt0D7/SDx5sV1H7AsBP6prQB4F1MhVzRmTJKZ9yl
LdB2kn0JB3ZwFYFqgq8dONSxGhJD7e00gFmEZZBkzb8kJuCx7NVtQG7bbLqefMOQ8dynFiEh0I+z
UODB+3uE8jUG151dIAyGpDddcpaYYESRQOk8FRJHFvp+hT9eQwbI/IbAcWO6AqUh7woJwTDvFQb2
486gB/AgXSSLEu4/MsBH6Cd3ri6dOXWOQMSKiejl6926rbLhkjyASr2At2LaoidhPPOzpZwrWs4a
kzT0cTgE9RlQj9sjU/QR3TenEhRgRDSitNaYo10oIF1b17ejjMeiCckMS7yFJH8i4U1bY9lo4hCX
jJyDb/nwkUZt7v2W0Z/lE/ke7S6058uB+C0OtbCU/3+Yjpc0TufgBB9mcCpjIa5W2ULu5AXLqDWY
4rmp15hbss7qT2PAS78Luz8sFV0qa/49anAwNfUyb/rgXXNpBpqi8UcMRWC5L3f05Xq3FsBkag82
BkvBxUHPljzmb6MFlXcLk+cSQeIPW16RRgmTr1/EySpWqiVkLPASdkn3ocNKcywRJ/vsZ2Ra4Waa
Ypk3s2t5oEKAi0Goynlrg9i1HzTHdC/wKOYd6i78ZUi239mCYpDEUUN7kHLOnolGpmetUYhaWGJn
r1e3gs5Vqr02/g5WpjtVuhX2l9JJuY+LNku1X779CoUYIhu7FjzmqaH7Oippcu+R/I9+qMMXEOaP
FmT2P9PRQ+ePTJabnieg7+J3QQgdlR+jiit81paiq7I2RJ+JycS5IqP7ZFnnFDCVwEsgZs48N0YT
gkV7KvuEoYklV1iX3lYYnNG8ioO6PU/076DetbR5fIeGrSW2ZOqwWkUqGbUFhaecFfqFdMWcEh+b
plmTrIF3sAFLAg+PT65PTLcVE4XG9w2CByOhC6eeXHuowM4qPaMsVayTP4NDEQyHG/rtL/vA/040
o2rM/ZOMekdVqZ++Pw2KQMmssXgHQKTik/rVQOVTGgGBMEmGQxHu7m3GoQmgTHebsH+q+66qOI87
i5ic+B6/Vrm/RtOA5vDDtec9YQ1yGBQzIBUeylv8smL4xMSi1s8uTeixxYPFNqnv6yArkITnTy/g
AroHIQvnYRHOeSSbb/3vOnavcqmSGlX4XOkV2irZfjB3kCUCrJg34kBojg8c5NaxkexU5rQkif1I
KsW75rHFwsBuEa9RA0R1YXkajMiqxxw6L6+tXe0pcjRVa6Su4Mm96CslBdDQ6zeBK/32yJV1NcnO
hanBlOUrxv9WmTbsjAQpn1vV4vK+T9IWRqRbz9K/djbkGDkMsMhgPTS8feqPW9K62Pc759Q1cud0
hBV3EF7r5IhX+SqC+bndy2PV/mAlfbnhhKMATWaTTbl6oB5OumxRyFqq20aYD0hwZqR+4Pjrb408
HR8JFcee05KLsi7VRbZBWvJ8v54V47Nj+H1jVcIAbxUMRrM4svL1MN/zrkdTLh9qR362hAXN1EBA
dJ6ly8Si7Ube783+S3J/EFi5Dp6Umo+h/aaFlJ6aqGxdLvi3SWfNDf9z624PJQwz3dj2e9agZ9bX
2RAPcVI4W45SDqdYiqkAOzJsz1Cw19xlVKn9tMlFLeCi/9cQn3yyCgpZ4D5hCZUlVu09Iih0w3Gt
o6sVjNIHXzx3iOOxoPuhN9+qq6Z5r3VaGlEFGch6JESaqHaAKHZs1oy81tcWn3E76pIvf8n4sSKu
B6tUwfkMTTWnRK6+ZR+KhN6h2smzQMlbO3zqRNBcUxzPOlgrmnGSeF0JTl1wmsYe2e5wdx9VcN+K
Ld1JZWJiuHXKMv/vkFpwQLyohPlv9RhU/3ZG5axUsivyWCs5lJACYMyRS6U8untPVd9Z2sITkW6h
a3xtDUpiD9WcP6XuyQISNb7+p+dnou1HuW0DIzCG7UkrkREwLeKKwJK3dEuM7d2BovSLOKbGYgCl
WEEmu3Nfka0wv4/giNgNWIF3UpPw6U99pKgbxbgWzrvZzniRIvsqcZLt07yqMuiLgLgXJsbcdxxV
muFFpq4wLLfNMnxJwaT5ekB9Cbc+vUcLFrFYDnimaECMX6TCxd6i2I5tMqT8gyTGdprcHon9lifk
zj3dlsCasHz2UIcfwV5CLOkk82sBaFEdUF/HsDsPcoH0ETunNOpkHHocx00KeCF3X3b6OoR4QvOi
3GLa8aJOf8FJFCgmEZliWxOh1HLUV3SDV9chpVt3duS/dZXTg3l4ewoqXBS9QM572e7BHyVW0B0D
FveHZdlQ7R4MNYLSn7ZJbVIeFBKhh59JpFTvq8g6fokRpxmBG5s+VHurIlvhxUhdbrOoQ2ElYH/g
FoDC7NrOJgQ7sqYruX+vJOX8KiHZAqoSga7LBZ44F8XdvRuBM4Tj3kSV5BR0i81dSA9oCmL1PDX5
1omj18OtyRXBqFBAIOa2FZE/GOLjnx9h3BSs2518Cy7BOMt6O2gHt5qkIick08sl2I2G7dibDfCT
y7dCXxve/JpEMNAJf367ws1R2ZAVY8YejnOuqqtO+d3n3i940qb16pccqpFL/d9g01kDP6POC2CT
HiEq4oa2PvEQ1OVtcOQZcOM/qYP48zs/I22yd6dVxHU98cjY+CwpQMYt7c8bJ44ti+7yfvxQBHrY
36xAtlTwd49LQTS19GGWN3dY4qRJSiFRPcoTOwMyy4LsYlkZJqbiOEwIVz0dhO+d5J5rzfnAKlq+
d48t2VvTcsz061YGOPksZ4p4K39kiFLQ9ylqhZTI0au8Jfld7oxJTht+qfp2dBHmP/KQmTQKli2B
LQb5GlBOusvR1L1euZepLJltGlUMdLdiKeqHpkz/9NrrTiTStRJaDljT6lMe1zleSY8zlRyMdAfd
3a5rXUEO5YvJ8CQwU/VNilRVzF38F6b3Q9ox3nHmYSeWN1ysfhd/R2mGu2CAvIQeukM5c4A0fzIp
xzvPJH7kNMNGKss/49udkjDNa9CLV25CsjfS21OoYwkDRKOjjWRfRUzYabpM3lgs/t4E1pIanPoe
YEQ32Kj0C0hnGjxGJByHG2lOpkN0x4J5mlhUxA7V23vRewBdgQ4DKpqYL+Ya2xb06FHdqv/HQbbd
WzXRcseX7CtZjR7d7dM4zlld9hHcQ2lj/UNIdRdKSZyq71O4MPIIaQksWGD2Wd+meLuVfQ/xLDda
qHAS/EqSlNO7awmF3nFEGe/uAtjZhlfFywZGGkAgPWX4uBu7AMSgYfHSsmYJZp5+RM0UYSYZMe2R
ea6h4GMC7HJqcBM5YFLpwKqmGWTXrMgvmv5KrEXCvEr/OqcjSPfpBJTaV8NO6vLAqzQKBmmRMrHr
LPdSkKd3SxnTbppI0+1NcvFSi5QmcEP3pD3Dzj9F13R3QYQje1qPQIn2fNA2EJKqcTjSv5hH+g1R
BCr8cuUWvjHLkmzWUE4cmrmCl8xLzdgo1yBldtKH22SnJzSzZx+JIYQ0qmIBAkfSxoqy+YbIMGub
Et1unfHnuGnZjS4GEdrYMswjBMm3Xw2SQSCepVVrkUZfutv3xLmR2/D6jkjxKeGIm5ixf+iIIrgS
IwXhr8EykWaAVeo3ZyWufsYRbk3c/pl542h3Ky62TXMdGlzNlKK2VLAZ5ThT/4VMI/AB9TRPZvFQ
bnzE7Jq9So+zHCK/TzoyyIFWjLasvgvJ0O36TPT04Ehf/yaVqKmdKDBYsSgGKY/k3jLQCnhWcFbK
Rm6mKEq9Du5aHSZQbb/9tzZPHely9+i9n3OUSID4fl4ekUNtj1T22j/KyqMSZN7paW215ErwrCCd
EXnnI0uYkXM92MwcVqQBIfmNK64DmbMLNe05LJ5gV8bLOXFNCM0vUTNhnjLXLy8bAAl25X/0ItLn
5OgcFu8Cxdw1muWddQysW30zi9mE/IBoBH27ykIMax09tfDXFNNJC7cMBVzrDU1z9f+sayWjRcxL
XXAzMX6MniIFl7PMn9j4PW6gQN0j3hpdcqoE+V9xgv2wCrPVW3tToFwTdJvSU/ej5VZq0B6GefyP
KzYHWu1qph6mlnvSG191blcVwrU0FiZMREbadiaQ3CMibqP3EjGpWv2MR+C0lsnAYBQQuGmgGbO+
e/2qEIjapGUlTrdOHML6eDCGe7FXKz+43dBUUCiNOto9c7gDGDrMtbtGOA3/xfaoQdLV3kFjCfyX
12tlMXs8AbLkrke7otqAYajI5lTUsbQu+z6DUpP1LXZAOOYJ+00VqbeqnxDqx+d2XQSYrUWF80PG
TIZagQrmozhZaJWqfs1C4IDhdeZH2CG7YXsKMpVWz3R7hJJrB7Hp66C+SGuzM6rTUCmEurfG3e4q
l8BZNqRRzgYRXgWvvuQp3Os0aPSjoxJG6qa/2EjqSnVKS0+32xh3vSJNWSJS2dvzVtQijcUMn85i
MxAahu/wwWpPw7YGoeVqB46Po1xy9pTnegwKZJKQX6xvzVl5+CE0cvoqFs8LwTwc477q50+/3JQi
RGv7aI9TqJ7sAP7uCF2amzmCWCjahwkTJiBhOiZ3P1X/1e4aMtSEHdJso3EE+xN2EwV8YUyP3HEW
PkbHii1mRGC+yq4OeWPwRx40xHpfQlXV5LapqriZKptL1G8FUILhUWU6fzWqg7/UuABGGKXoFJaF
P0oJaWb4fE69Pbig805oVILBTHjhUCEtfv+aeKzZ6QsbmMaLQdJ467cQEyh3M744sTLWPlnPrMGE
MGahHDiUy5QaJYM9mv/yQUcBmZMvHM0CVoKOgWsczPiqwgyknBGbIuAH6khvyVkueaqTfYttS/dD
XKynJylDaiVYXajxUDDl27p4rn3BSsvvbieAJsFZXM/G/e6hrGXAtoOwKMVIeCYUkKs9Qk1gMHm6
Kz5dGpptd2NKOT4ebsf1HK2G5m3M0Rtcda1nJyXpmIZRS7kyQgkhp+vdMCJ3CCCnSaRTz/hSOvqm
aCuUHtCaMso8h6w9cBdyA50+5LW49JDIp+FeHGVf/k7VtGOhiYMRr9rjVVRpQ3jQSqKTao83uwq+
iR5pmd58Dx0/B4fbNT84nV7Fr05JaxgMRjEtqoqTqfudYhapm2TMiJj/2J5OONkyMEXtcex6nLum
h87yxBJqUT8bYXU48M+c4ZEwPie4ndD+cNLRasuWQKV50BDO5DQnMKziv5Arz8BOGr/pWLoS5gHP
8FYVIx3WIgI+RdlYdsc4P5sn3dgUaC2TKps2NrX3rm1O2GPl7X24ZDjGEuQLyD6bI85Y/vmTO6Nq
rXxF+L0DS8woJhYXWeu2gfl3XwKmiofT1kemUDVA+i3iodmKtY1jc081H+HHOa/6fgfZxdY9IAdJ
q+cuNSMEGRyHfbh6EYYTCUYv2KNC/IEX1/QqZTfw0mtgbCT1dnwwC9tf4cTicp8dBWJx2okO2JiZ
WsihW5g4YLWpMu4QF34brVpHw8uZpl3A3yegnqaSHS477GYDbLuE2VkjDtVuuEiaYZkSQQYhKedF
1pdHvBVpTjQTdF3tTRhwArw2/+lAKE/k5ifXmR23Cwu+JlGqAjlz6EQlK/kxIEypoUMbthj5B9Z2
GNLfXL2TSXQrSjYVOkiACl7xEjtj0PFQL5i/HDpYj2SRv2QIlIgS55PXT+Uv+Q3F99nkbZDdrM9v
iYTX5h7niOsHWS3B3H1ui9QOpadH4HbFnuCjFut9j5oefNADzqZ8f7GRIHDqMbrO+XucNKtrZswJ
PuxPCxRSiUEKBR/uPv+Rh45IBExSa67AUZuskK7SN4xFKGCNC/fkoz2coFhUS8jaSK8m0LNpPDuY
i7k2m3jcbKTVKbMHT2VtxllRUY5nzwIGcpUz6gQsdR9i8AlNJe4yhWgTE0MW+7iCy49oZVDlKAba
hIMroN+aNfLAuVlddZXLfv2E8Ow7YH+dMdcEtG2CwLVu44eNt3dC0iFxWYvbtQ9TVV5dE5xdvkAM
7QKiDS/6NgGMGyeEvwCbBchS5GC8WnIgXqOzMAlYbRAgiibNmYNuED9nAlgjVUsF+4nWEfMcdOJP
IceQc0IbNjaIv+G4A1sakpCh4ge0aVRKu4xHpemDYBi5ELqBU5loWQFNiQoR6FX3AuIzuSowV2uN
yCYdYIMbYHZNqBLIZm8atnigy5CQEbre9ff0ZhjwmFx3Z9U1felIyQQ7xc0RPCTM09iXtS47vggL
ESpfFs93jS3WLZCAtg/oO/TzZWpVCQ69ahUEDVaaPi27uC7PK3kBCP3yF+2TcW7mVl3AIwwloTSz
swLfeZy32peYlbid2D0pmT3bAQItQn5wPWlsKo90KxCFWgEtFnM7nGE9+nB4+cGXKO+XAWbyQb+z
cYQYYkGlI+9tOKdvtUj1l+bVi7eGklIiswYk6dhSqXVe+g2KhSb1dMfwoA13+6dxp4KPrh/BpzWh
428lL41Jhi2byucPk6keG2AOqt7KY58FvrX6hf84hEk1z8WbLBg2x6j2B4GKFK7iK75OweqU3/jd
sMKcomfClumZbTJFS3G8LZohEEhea9yA/dLjWNkNRE9dWiv+sDOvneOlTg2tIcRuJ4awB58rRWqc
rkMDZWeKYWWr7ERS3yij3QaXP4E4wz9BVBp6uVwUYsTCsf+s8m+TkN4EPEmG6Yk2cg3kz+tKwSQe
wFwyCQQowW9WiSQveFMkos4wAow5H8tfkZVLDwmyyyD1yYaBcx/HdQr2/9uKEEEIMTPoOIEmxW54
a7GzMv8QVAPxG4x0czzSAcejacK74rcNn/tWnZB6bctKoY2UKdC2rOSwaHG9RUlJW3P1IBIiv14r
ni701oVBsRn21d9Gt6xz1M+uAPIayY8aGo0ZfxPES0bGpd+Yhdo6UP/kNOLEJ8ioikZRgRDHGWJx
9afAHzfRaWzuTmYouNuoi5fmbK77WlpHMxXWfv97oxpL16XHT1onqHKr0YA3vRPH8RmDfTNhReHB
VcKbpLJA4n/1kxorh+i1kJGMYpvgCccjR7aN89+xOoHc+8RaZVGRO78HvuEZjxlYUN0cm2p0qeUE
QmHLOBkZ+Dv4/oME/0A9lXlqb66roqyuX2o5Ko8XPTQSPoOWXnq9RO4VZ07vkhblJsyZkIZxzUpf
3Z6c0011nfb7GtvQQQtupdYtjtHb88lgn9/D7l01aLSC73LtLwtBeYUHybK0hIhfPixv3wFUZjz5
VJ8ItMF2q6f/bmJgCVDQhNk7S/9R84JzruN39suzY86dA/T8b0LSu4srEXJ6iso7V4XzP1WXU109
perEKv9f99rJ2syOuxIMQsSmGCQ7OEwxGE8U+EvDTK/CSYPDCxB1vJcb2a80ah172PLvKJTAm3AY
sWLKCjWGkLG/eockZ3iCsevDECo6FUGsJpC8aQ/t8l8jon8JHCDETSMckXkOUMuSCQ8M4ljg0eOK
0tjILQozZ232VrqcaoZuqivbmj6HwhWo2BiGb2JMZlkVpQXaznZ0KXxQbFsl6QkN/ZO+oAhRGweK
INiuGW//MbfkHHmkEOeaoVBh47gWt+bXwBnneYtpFpKnIL08ZLZybZ5ddVBvGz8SRMCPgeUNxFnx
CQFbwMEnjTI6gaMmoEuYvlM4osZ6hAHImvLHd2kjeMRCCI0L65FxcEMdPVHuLDzbTYRV8MDaVwYG
WvBsX5xa8O6CGFe+8NEn4pK8QWOqE4ZwkkjicEC3V3jKGeQW9GeWIW92OewlIy1SgR6DC51PZgYW
6KF0rnApGs/GfjQZWPkfyLYRVA938Z1NZPpaXlIPaWkYaLJ8P1QZO8fLbih3qDzWHl+2xUIKxeXx
TpEapnqggy+ys8HxrMtr4OnCtqUMldg5mL+rIPQVmFQ1B7GDIc7183TbrdQMsm5Xl/nqvqTrMIX/
z4RFMy0xlK25rShtTvfOrrDBEqatzFNemluQ+6LqVLEBUKfJNk+NluhE/MwQZBDXm8ALcZqxVMHW
4RywgXN6WmFt2bKBgxHZUL46HU16AdMxa+G4UvdLbu+v7L2uilAFfiELfQ4Yod3ged6uRv85IymW
sGsAyX6gm+EJemDfYavun0aGiw5oxdZRhm/MVa0Oe8gRTKkZ6UfBg3RBC/slErcJwYGTl8YVmCqU
iGPuVMpw6gblHBBKSPuwgCy/lgX1CgjiQeyB7CbKt+ADGMtYXNh5iQT19NG570gzDxsSu7lIIneJ
SSLL7UXjsVTM8ExHjOiO3zdlhCeIKUZLfEINa3IgKC4JYA/MJ4MY2stDFkPXi+GRYrT9PobkE/oK
V8fZdCxZM8DvUtMdBd++K6OlCxA8skNrhGUlFd8m6vyR02KB0T+qArUFqjob8mD4Y8e8/+3Sy+60
jrGDtMLRIKg9CXGBOscfdk5ZtdWnQlvWw7B1i1TRXAuT0j25XHOGWMkc+GYn37EnjhpM0vCJ3Fi3
ZSsE4a0QZIev4DL1B1l2wnWDALdJGowF8nBHyc4GMcb9ZRHZtM1z7Hocu39sV5iQkKYtpCEOI2rq
OuQejyMSSAX3/ZsxJjIF/2VUGfZjG+NkiMMkqNILROFMIyXB5mmfiyCV/ZM1iKARAmyKayICGJvY
RvCk1XqDANDiuwXBfpwn/QupAuvzp+R8BNsYQnvSDemUY67hA1zKbL/l+g6yd9MpyfRjSAiIfuzw
NyoLQ5rJp0MKBI9jl54V++hvXUuUT/65VsigbwmYy847q1vmcXv7ifxB3OUg9I8hvWWlH9EtD7ZU
CiGAavy4Br+jLzqoVhpFtvX5W1UoTi1Zr3Nnul0eab1vzRtDiRzxRj86yhw0jKvQ464XJp8TJxRK
/pjLT3mkW5jnNGj38aUtAJnJ6UGma/DL2kTyjRP2yLvRoLk/sCkWFM1A7TAdzJ1gSuqYf3o5fzXv
o/TsIT2dHnJRRU+qDhXBA6Gh7XIE+XXn+I7YpK/cmRHvy/mskhd0YHSE60GTFdXUrdcOYG9qcY4U
o428x1stqagPdRMRuPkNr9ZaAF6FZKDUFya3vtf9cbBO7Nbd5Dhdi7LJPI/e89Nvulm9bAPYfkfO
T/vXCeKSvctyXmSJbIpnOqvLnYro8azSH/x873Mc3oWwbvCtvJnyW00jcE8Y7ar5E3ppQfSAesxH
lKRmiwSgzM7PWV+2B4n/SnR4693qwf3lNUdoC3OAvBqLi6fE21F40hgBEd7/X/K1cZSMrTMszodd
1+w4x/pH3+Lren7sPNyAWFBZApFY92Vq4tX9JCYlfvrXiR+hBqCuIKqYGveNN+Br2rjPp9rCcVHp
yOOoz9qAwxR9BXe5DCUaNa1K4ZOsVw4BQyBUYZvCzKGRRP/SKUdeuHN2bd9ArCnUlFd11ZQlU5rm
5+W2CArkcb/vHe+YsSkF3OJGEbiFzi3ibM+hzZweqwKfi3cPofRjHcT8+h1W4UKTZu+KRs6Wigq6
gwDbpai2I43moBpnC3OGsi1gBijnsXQNlglBGsepX6z42P7FbfWNlUsnrKEivFNOJpJKFE9gC3l8
9stwZfSP10q6Ku6rMM5l1Q33tS1xXnYHzaNDUZOwAgepxq0E8FVdmU3iGmFS3Xjp+ns1xCqYZzr8
LyZI21sbPN9S0qFw2YffsilLjl0aghg0QU8cJG/LemuNjZsdC/yKmZUdrstU9Y6YeGEAgLSU123p
xcamChKa92Btyc7sH4psVQiqYvQUhUIf67DEQ+z30WX++2YGfED26+k+QI64roCGGmGKL0XsD81j
QgybZLJC6o6tbnfbU2BJrw/i33Wf9g5dL+s0Gopue8DbnODVz2Ga6xbdGba/5TjZ7VVU+aktwtzo
gB2alhSshwr6ljIAhSzP35kOMwVBWuwM1cy+l61ohTSbpqWDljIkc/yrKGGgVmwJUco7bgZ6vocW
SnSf9XTa6XaGRfiv9QQU+dvxeOZnpcTJxjSXqYRX1ztauBqr0lX23+nZcB1WWMx2wBCmvKdqhIz1
wm4angCcE9YL0Mvg8O68EfWOM1DPxbhXH1AO5yJmwQ14FQIwPhzhYzyt7OhBZQyX5Gmfs2rBRRQw
CyP2/FaVus87EKd+hP4h933kLdNuaeebeNP3ham9o1SZqAGHLU7CQeXt/gXkB+mj8IX3owgprJED
q5G/8q39mzbi7Z5I7Cg4uQGn3F7SXDM9DgPQScMNqCV72xGUlBS5C/f/nn+8GKxceKf3z78UBBwC
c2jvxdcd9C3Q5LekdMddWWwPgfPUW/M7q+kx0UhY04G/9oTEgpZpgE4YpC9HeZDmF77G5/ofZajT
8eUumAsheqBPic3S1hvlzKMoIIVv3ZSEYuB3H9zpZWSEeJjXPf7dtCPm2mvf73keIPG269VphP+N
LNjXkZ0/c6sGv0qAh5TcbPTCH7eFoRFYrg11Ip/2S3QmBGQ8yIhyAOfgVttAjYA5WNTP7fvJ2ReC
Y50YpPb/vN0PSkWiHjPOTokmcxVZf/44GbMRbhfq8dTzaxP5dLW1BJhHI5IpvUo/DUW8Stg0EJz9
vXbFluMj3M5meUHUabZSsUQQ9AUrly0Kc4BIA7t+hLXlN0TADrj33I4sOpK32K1DaBXdHKcLG5Tb
Y+TPIU7prW+mjHKIctuBzCnsYf/WKORuesZmGAfOdYDZxGj30KV7eb8PKyb9R5N8ELT8ejPJyGEX
5uX5zTuo7/ciUIUZiYHB5IFlHSehvcojlYF3u1k7E6eoRbjw6v//PCghzCB4PQ2YzFylrdp/r2O8
p7iIfKNQzffkuSh0QONc/OoMlADVGloTaGvhKxSXXN9AxFAoT4a84BEqPg3T6ciTcejxzO1ESOtM
g6V+gFwuQbVrSZ7sJcxSxuZOEGOlHOYtgHxfBcc2K/zv1qZwzQFnh+WEBiYLIVabdOYGJzYcksb2
kAMX4kGqQItxyztodjZR9dvrALSAduvkYAT+9lCeHORW9CmDFZfHoRU9/lPmFAlLxXsi8IQE2twA
Yx0m97rq6zOqGQcYw7mQ6D/D7dFYHIFte2oThWUZt42Xn4bymqnId4B4sE9eV0TJWJC8BWQ9NWFy
PkPxqeCn1RtICXsybOKO6tNDnuUnCPb+bumjilMbYPFLj4vPHKvpsFAz8GIzGAzGpioadaBXJKNg
U/NgNfb/79jJiGhGqPizdhWRL28XvyhNhbpJ0fzS8h8K9kEIInwOcHdmp7B19RPWDMaNX3gmC4h7
ZWfeAtJi/d5rYaM6ZSocBBf6f/J8ZxLs6DCDWFO5vVq2foY+hXZGIXemOKZBwdxVgW1BLniG+nAY
2BrORNXaBb8AIqJwxPMTaGmtZVGVR09b4M0o1AIJTmF6MfXuvdouJfC2LjxPcfPor+MDa/iq3SRh
/S+aSV5utEqh8NwKQSBp88n+ZgD0zLKHHJn0fMVenDoglP5hhKChieq7VdM2mZAAPyDLJAAYu/aZ
Bnr13ul9DBt/KtGz+Km8jwDoR1HYm1NRZ8d28LQ4ZxvWxXno28NsC4LKF4Jg9DrllnIt+dK3U7C6
y0xtf78n4uKfIPgFaYc4KCQqVxThSunyoE+ua+GnsW/jm81ipNYb6WNGeadhE+5RCDfenkYWiJ8g
Hz1kEtU8OPrVACMO/sJ2wP7Erc4TEnyoY6wIuf3rzsojY9N7WikiTszigN5xlG5fhOgfacQbK4QF
i4ag9mn0d1n07xyyVKRQCmSDMdpQzOuOWUIVsmeWvORrgWA8zN8S1QMZNStChLciyYNGnqMjJ4kI
xdh19lgZvaZleDtBXDoINKAy/GF5O041eUqKbIamD9tmdg+DMugwfGPZTbio4tZP7TSIBbpnPs20
jQeaZZ2+3VBGquV9xEt+IMefcQLkxzlK56YOyEl456QRLczSFqju61wrK8yihbiWNLqvOoM2zsut
Qjz4Vm/Q1OS67/1y2NLFFcSC6pqasNQDAmS+Q67pArWV541IGdLDa4jLc8NrirZNL8SYqELUiH+I
SWg53WhEB5XCFRSylxuhkJNNTv7HEHjPOzg+/WlE0j+usSzAob/DbmHpD8cPtWb3BZlDA0VCaoj0
ul4uWINrx8XQejkYePP+zv+hmNNEP+mmwUrp38SuPDZ4YCht8VUHBjFmScICMZOfd/Jb1EfLqyHT
QrZiMFFsARDh7Ap659UuqrOylNfvAzDWtBBQkPqtqJk3fHAzM0Kn9bS+QTNTq5+cFLRoZZUTmo2/
f5QVBRiUb4p6i1ejp5/pqLKsCELuzM2idJnod3hBqdK10lEkO07PifI7am8K1XOVJuNQxUu5IF6a
F6mpSXcJP1AG1eD3Y+QQVl7qwpjDEdSMV079P4CPKLn/T6Vphhvn02aHVz3C2U5PrGS5z2mHqaMa
VRp3U0yeRQnx0/iWF5GFtdEAQSFChS44ZhO3Hv11FDSSw/UrWd8IB3MzIKRYgDzaNB7/do+wYT5s
w3EGsV+9YsNd7bqAp4fwMCX5WW/lCRYAOQUAlIAhhWl4dTs3nqayeHtGeO6uwYmSQzCodm6FB66s
AQfaED2km7d3QonDdNn81+7docXazisJ+X54wDDf6fjS+ys2BDLBCuYldo14z48CTXMkWUJ92I/1
5hpLgOOGXCv5nm80ZsLHLdTMWUo7z6UQaWctl/CXNCg1wnshwCVicBPDvW53MMQMUV7VI4MbhVQi
KPdHuHFFOkU/Sbu2IZ2WYMTGbEeBHqHVBJV0yzzClMb+6h0m2EGJC0bIGNUrcUjnRmKc0ixb6oXB
oyvM37LTZU1jjpiw+/dFgcXLAC6e+2TSP9C9NyyIKZBvWAq6PeS/T5bjnj8Fwv8T1ldezr+6hJzT
WSJdE7+FkileyxaQHqhJ4+HJOt9/XVb98L/8fIpIWXWQE1wlxLQ4UJeACc+XF5YD651aj+7KI7KU
c9k9pcwEEOSVwo+76k4+6m14zhpsUgVEuGG2gJ6rmHI2zEjb4Xyipt3lMa8jdpv6yWYn3rCreCoL
gCmPGR7MfxFLYchng8Ns5fnK/ecxkSkZpAwiOwV7x9H++ba7w7mhkm6VzPQecoX2RIQaBSvMjsl4
iDdPdF5nI32OPjXY+iPz8G+7JRKrwROmZpR+fjGQ2/nTte2AdGR/nHxYKQy59Gz7y/z4Jd/e/oHt
+80tWkfmwTuYXKukMX+35kpD8HJOwKtUWJ77uYULMeAgxtlktZoRNihJIROGIZxvm/ur0UCoY9TB
NcePI9TnKSSmKEvj/IOJAt4g0I49F8LaSYRkyLG/acrYA3B6m8jzi/fvI8SL/87zCkHzZ9j9ytO4
Qpa8R0nNYmMuyqOpDbIHitTIMtveir602YQdZC8bAaRi9q6P4O2lR3UAjoeM54xEWbjblJD9o8Wb
WGXtqz8k/oJib25dGYO4hWt2yIbl/2CTvyjhtkp2wErhOjNUhumIuYNK3XAWrzA1ZIiczxjxyW9J
ltfAYW9CNkgcnLtRchiwyrLHF+8Pvnvrm1L7y3OBkHHaC8W4hVewfRZVjXlk/nJ8UwLWPA9s1zWx
ewOhdybVJZ+7r8tUWDl6XOdsxLnPAOMbJYiOM1dvfFeDkN/9F62TEc8n7SYQHcIL1N65X9gd0N/2
vOgD/nGpFHKt7TTrkZk57mXaNg+PHRtVJbe35mZsg4Ao5L3xOsNccj8RgKQMhXCoYtjhcPnpDVu/
KBe6Xs++D/mAgavhWDwfbBlGvEXw6SF0EVi3LeVGNDhv1LNaATTTgEmYcapHIMM4OfljyQ2Pt3zs
b8wkAvyH7GK8ZrRYLbB7tTdmbvBRDQhLPFhsLVlJq+9TzhCHwE9jUsygpa+DahDbkFAzAevQMJoU
iNTtkccmp9guQ3hY2AZDTlYVIrfZo75CTm1qroFBDhtDOb71Vxjhr59/biL1dk72K40cciTQSWtq
1hh77GaPCBVkP/pNAX65k/dhSvJau91Nc5pumzdha+7/AhLgnnaxnPQlbzWdk1BhdD8A28fAnHtl
jnXaPoYG38Rxh+IP3QD1JcADbC30tLR10LTn//v5+ntYD13QtGBSgOh2jAMgh8F9z2sTZC1IQXmb
U/1zkuVX6hnxifZ5kx//7lVekRtmd4m+EZgNsfEUKeSeFdbCj81HGWJxADQ7Wi61sIfDzJHbuF8w
xZ0BWq+EFQZMe663RgkskhMJ7oHt3KHabL8twWJQyZLE8oxsGwuj165j2h3MwfpHcecl3Uei+sEj
i+blqWMakrpr8gc6h6mqkZj4d0xMuRs+a2Vu4hBrZdfdBiKclNTOK/9YE0jF62TNaL739hIfw+T3
SZsVJVTXmKcMrK2e1Qia8Hn02VRHoDLGzeO/ATYAI8Px8u6QgjCQCpOpblp38V0FL+56VjsFaVdn
EBLI5z1fSNiAbcYavB9jyiyd+pSTZcLe0KOUXbbLe94/Wm7CRy2vUE6QsJp9cIa/IcTHgKWsP0Mg
YlKq1XmVeUgJZDOGA4zweYnUEf/7TrtRxSdWGZP4JGjN4pcCrkUHBeP+19jy9WI0rS72MFQ7HeJM
XKv12ussdDWcQUdWTZWkdFzfnEchfFP03eGYHyNlbQwXeYnQoWW2YIdRjXQHryuCMqbH5bB/cmUT
PrpA+/xGe6xQ38/PZbW8RLIrruah7jrfVLdmEn6jQQngfUrjMhdbUVHJVv0i9QU04NbaEv2T4AGw
ubqwwujXM09wImWgFNDIU/JkdlcbjkCyysttOdOh70c9wFplg+FaRznqEhuVDNNpYsfLKCqNxkQW
fpOOnoHistBzf7fWYcjQ4oNeJ55KAWptxq8dIImiwTUytqokDAE992lDLii159Ub2J9cDLuf7Iu6
GuDF4D7fgx6TqRT4UiZnDq/ws6TzUD4Zaey5dOUlQUvtXrgTeyikVJ6IRYje9KfZ+SjzlHH6xp7N
x6SA8XSLUuk3ziGIxLis2CYsDPsgd7gDpTl8DZG/AmC0qY37A0V2bNyunNNyZUhwLl9TaO6L3Xbl
FlhW18o02v0YhfnecCn0Irj4zSBo+gFiwooo2Mr7sJpscLhWLJh/lmQJ+DpHIzYSFCMuAv2fAMmP
Hz6MWmawrP4ab9z4vuXr9ApRGItPImb1CX2AhmExAgRmi21+H9AJvRl0DtVZt0s+xGfiTdB73V2i
8RhT64KFmcTMkvSSxuyVaoZMbkkc1eMa7r4BKR5KBJwkKYIRjlmzsgA9TUcGl96/kB99C5IZjjzd
eLQUr4hlPuwK7xE8N13uRxqepPAGqQ5IPxVDU0ZhBnslPDIanghjZPy9hWecutHFnTSVBcQmeT1U
s687a7qDkpQENV43nV2+qMGD+YaJCReq9IQHTBGfgUDfSfx2AaPlz8ecwYLYqgmkEU6wm24VECNB
7n3Xai925aKa2eH41KpTj5O3tVVuc3OYa7bCdsupr8UR9WN/UfyneKVmpkQCS0bpGWPa7cG2b/Qm
ZP8nawwijVk74DuAOXA+FmOhJE70pCauJoblUi7L5hvDfGtgV8JZ9k49sUYpiBzKZdOdi2yjqH1x
QPxyftC0JvGSpqsIAzT1aNQLR2fY7GZP4N7OK1e/yIDxB1/b1K0boJhq/iiAQidKkZOZlj8Xgphh
Yof5zWFqJEHn8cDCF5W88xSQ7P8qTk5gBMcBZiLro4q3RFZMSA5UKAZs0jU/IqODe70qIjRMrgSP
DS/QA5yNaqW62ZRUcfef1RxFD7BObc4tbD2eN6TgNAgZ9Mbw8KCL4uGYCNjY95MjLlwFHT92U5HM
W9vgU8S7VB9nUXl05LKHPbgcNboyD88SRByXttVIDBkTAxPV4MX1mz4F2xOOlKJ6krExNkMUpLqf
DswvbWsIOWtgqYSGrs3HVQU+6Aajla8tAKux5Y43OA5O6QMMK6fuPKMd1EYsKn9FsuJVQC1I3E3E
GsCJnYcejTvqeBOzQte5xpjHYPZx0/CWO0lwodWE4aw8jfzHhZ3C2CJu1VOWQw3GngDpJEAhSbwr
/bWZx+bWx99WHSPiBsQ07XS2DzCXuc4EWIAmkk1BE7L1U9uGkxKWtMsZOAA1JYkqG2N81Oy0hyY6
xkfamS0c5zbuJK01G8bssP/+yAyk+Mmp8xlKY4iL1CcrMpROwUCTCfcn2hwcmgxGr4SltgFOd1qG
4f8Zno7WpHwsHtO2TRYoGYDQPTBcoN1rerwPKGEn4UzPgRYspGp6FCCHYHNwW6pMMlS2DHH+fppL
pKi4TME2UT8Ed8jNyJbZe8p9RPRaOsO3mTXfuZXES+sc1MPgO2KelQIuXHu36WZQ0n0n8/wD0tNO
byMFNeJ3sEIsDmBEewH6pz2NgC+ZlZOq1R8bfEPMLHYmB24zcp0rH4x75HJH1Kx7qoYNrP9kXWL9
HaMt5gvsaQnkSdckBrRAQD6PINHw0b73Swn0W0qEu18K7/lWIY9lDqlHYBtn69NUQzkQOs46XjlY
aaYLr5HMG43RdkVZKe3iocpP7872Z38LTHgNBx03A48sNQtaa6cztYBef4ey9rg8uKtgL6LgR/M2
f8rAj7mcIwBTW8+gA5mwQTzyd4B4IMuXuwmehfzQoQq7wnKHPHHZfaqoEqxaSmPfhm5+6vzjmG4i
0rMvBDT2oVT+4H3EC6dda1rREMugtRNglmLFzLLZvRIkXLE1YskGf8BsJ5wpJHu6Ly0Y/G5crCcy
sd9awSTjQ/n9ZLRni8tfsXfVtBgdesv+e5NigVa+GLQMvchW47YwqTJw+3Xj9NrYejcxNaYpxhGS
gLxLTOwxOUMtMQT52n9JdOcvGjrUXnFU+bqCGxDPDdRkstew0shQuJfea0axgBZ/M0C/8/ASI8p8
XlOWndZpRGpweu/dpM68JyUnzyydsCQB0QfSCnbccQuGpkBcfpj9Ee9RRv2pvR3fJG4niGc8bTAW
6YsuBgf0Z3fAw9PlDIkN5qJMg46Eetvo7IZ51dZCDDbFtqljfmhm8Jf0kKtUA9g8oI5naxE4wHCU
H0R91CB3TSPSfER8eahDwM+Y916ya2CUPrLareQpNODk6VBLPJlzxwNK4yzqEm73f2lwma0pwM4B
NO2CremQgKGgaB0KRF8X0G+MQiwUcQuSLoWcYkv8YXZY9V61Fj5hrCqfdmCp7R6wZNFsvGBp1Muo
FIuydTjN0T686kHt5v22G74AD7bkeX1HcRhPRV5NJxCTmbrvhT4MMO+gnZgTRt6N9htKCD7wa2uC
qx1nQr6XDQhSXXY7fpAVE8vkLe81IC+dSKWE/1//RdvD9/K5+ATQ/0t1AYbR8mr8RWbVwB1lKwE0
HlKSrgc/mOifxvcrhX955nly3vw3QqNFvlVh0b6ECwgNsZ889BFigve+IxsuCq/plKy6rh+l163S
9lZeVq5Veb5p0FOKJi7v8a+ZgHjrazzsdn1NOk+UEGXGQ1MTOztZEHjkDmO+6pjVATvv/a+xfUKo
Dh47gQDBZ/8LV6hIE8z0ajCPpwwbuuR6NEWNaCAGt0kvKjGdVZ0+9XU9ZcImL323ic9m9TfumINS
iMYJ3WRzw9weFKYGrxsN2SE6MPyo1SPCkBpWau3JGFP4BrfRFrYY7fl2CCz3T1N3a4j8vN5roUFJ
qrdTXzD0lUlzh3i7AHu3wK4GblfFsimta+LFaorQo7i32XhQ356Eg8GF1BwHuwBrusf1uao6+FL9
+P9CxyRwK53bm7nUoBRRLM9JTrcly5N3fxgwuxY1Qly1/xgDYIKM8wZklJNW5LbbY+rezgOKAfSB
AMXtEzoqNyDBwh2Fbo6UjTpbP6JilOe6rHz+zAdFG066cMdzIMn3IaAURLaPKmIiDaFlXgkFMfu7
MM3Y61qnlNDxhfb5pLP+mUtcpShYuwZbhMlI/rS7mdbRMKuhfxaOvM83CuSjSQXPwfI+SMSOPTek
roI6gNcABWwbjRLnoIuDJ3WBfbGNRftEKDqvd7Uzp/oS6UTSup3NoPg2OGaYePAF2htrV6Hi+AvI
pTH+5+XtAM3jdeKdBYSiyV9SO+wlxCchdc+rIHW9RHZeRmPRdUfXY7OwPm2V4IYD3e7w/RS12rQR
9DhDjTGw/1jnU6zSV+VV+/ZeTSPaNCm5T3dhJhe2s3/TKRYVWqkgOjqbvdBnWlEG+PdF8mVSn1b2
XxCbEI8EYklGtUp9CsyqpJzrxE23jiZwtHYWrISzEYKjVfSC3uxieMT/9DxPC53aKIQsbIbdoUJV
MHJLTKtzu4z4AL3fqj4ESZWdiZ/blbZt7gT22DP/zSFo3EhEspT3zRCSi5QZikf2Bynq245P/McY
c6xlFk9RlIs2ninnWAqChNjvlfK1Mk0CBHLtFB20snhtDOl3mAsNjZQLfogc+Qp42V7cJ5mcbcZ2
2PTfcqs2DMtyyEsOIMnSd5C0C3Fcb9aA/e6Upm9w/DvPTf1gXyYryX1hcSoCEeimLOFLyu8sc1IH
OAaWmwxoLJXftAGeehN4sh1BKu4SN0PEKfgqwmT3eud3GW1Ta1JC2xirvrDHICJ7YsSw0Q2auhcg
QuLksK9YoEi3QQpoHbno4qWIRsX0G6zHPJPDGpBuWltftK9/lj3clancpA8MO8FJcobeH4TASyJk
anei8vdXQ+J8vsmS5/zubnzPMZsS5XWJo6V9vdILL5djUZ5IiI972n/ryOZnbKKF54lJyYnJqs1e
V1MPd+v26ovNbvLiyRU5v0R+IwkHBdLG6FojY1oqEHPpQ3uiH1nenBfDY15/KQOhBXldvGMH7Q6J
NwvekgypeAQgY5pJl7E6fzUZ45OLAYf6slm2xlwaJR6d8BV55lJpn46SxWx2DEexrweuMVKmmraI
WAWGuaaJ643xD9iDVUvROHx1DMyyywBDnrBXjEYxDdC6Ixa8q1BSzOYsoDC6v4D1V8/PIEHqgrjs
xqDVz+icxhewOaN8xu7yYyoh3yXMhLkdtSy1tBI1HK0gwRgo6E9ik4UWfj8Cz13x1P3CRFhJA7EH
wzSS4TtbCYJYg42B4ZDEa2zN2feTkIypEj7Mo4eks4I5JIi7geFfkYWhbM/3xQlckpqNINDtv2F/
IJQ9+aQ4ZuiMxQ70taJwEJ5Q/dYFnnrs7cjWVi2c38LJ6Q8CIpvmaMiNz1lGnGl39tKvWI0MjoKH
dAlsUuTcQrw7nWTJhyV166sNk6kY8qGg/LXFj1W3mjK/QfnyXl4EO3IcC8UUifOGvb+vr1CGA9yB
KhaaXxDaJhgy97Xm75zEu7c4gu4MC4BQTjm/Jhi40mEQX+Ri9jvVXMZR9fPBCmBP83K5mQ3Wed/k
iWWqdq5CIw8X2pcIdXaq1eP7RJOQNKux8iEoRD68/EyZ+f/pDrISUOqdDQqq93bv/rIzd1SG9M9a
fDkT7IHsyqzBf/IoJzJ7kzHHQRsQGm+pt2ZYFkhXs8xCjNfZpOn/SWhokjh8/jt4tRov/E5fAhaS
WBK6DolE66kdt2TgGb4SrYeIBHLBkP/saFWk8z2CyzZ3pvGorqkFYY58preubZUBxH/vJWW4DVJ1
oLHT43SWzHYpIXDVAwnTEaAtNUFUkuLwNVanL58Wm5VIIcKjrXTm8ex+L6v5RgRNEOoHbFTYhsPl
YkH1lImeI9CKh5whmiZJfHdumykFcmw0oUg10fDsE9k15Oz6u4PidXELkEVQ4cATb/H6R4QuqiIM
7sy+nbrbf4RHHh0M7nKyslEiVWSlA9j61EBgx9pGepbzvpxFE+fx3Xxf7Ms9QoCwOfqbJnzijKZu
CtXp9aDjNxiOmVoNTMGWxr1OTdZxT1ZLxY7IRhWQHG6vhhE4DGhiUiNcra8I0b4rG4x0XE1VDa3W
6JZspfSfGzE4OoaPtt9srpHdMApOVSZboCE5qn/xQecf2SYK6isV9q2pJQ2H4JG3B6fBGgc4vh7m
LbO4Px46n8i1Hhly/A80qURZyRnoGwX4HOZuvclWjjjLcp45jqI9Yc0T14kNwm3v0snizVNd4j/s
T1USevnjI9vW53bi3FO5bI9UkgbeIhvyB9glS9Y5w3nmF/2AqFAZUDEVogpBl23ieRpl7fcAAyS0
WOpAmzIho9mPtIRFZU+GQkm0gycQibcho2lcKggrK7tKFQK0tig3fMm9Jz7vRbsoYu9z/IA5c7ZH
qM7RuiGkaSrB9JT7y9jUa/ThZpNNVZPALYizZUUqLkYSp4E9ndASg5uBJdHfz3JJS80B7sKMGpec
mIwm9blT0U8ybzaVoLfwTm/gRjFNg841qNTaSYAUlo6qxLf01gdqLsylffluB6ZmnTgHOsqhJcHE
9fKyoJDQkruNEGJ3ubJhRFdY7/jUo0+9Pivls3SxbeTtNj+/BD90TDrRNTVuAl3BGDh/ZSCDE5BQ
ueFxvDpByxRN8VWQC/MW6YdoRNjFYQg6H9OaHxdlGBNAknL3IoDefzvjTBKDIvyxjGfvdTGZ09QH
U6ncj+gSXMKpPTI+iCTE9OrCnrwwSPRSA7WnHWfV+Zgt9GXBrDQaAcBP68VTy0MA5I9crwKPYcaO
9KPnaQRg4H5mCfI+p7Kru15o0lCSjGMLIhOpV/vJjlv4Xb0OEdtfvTxvnR9k6aT9Azpoj2abx84j
PbeTDccAaVwY726vMEOfE/VdkgjgMrHv8pDolhmPavya+nHhpMUKw+MsRfp2Tt4wDjGqFUvZm7bS
PC56bxii+kGfWbVUAvJm6k430aNu+kcey9mpoRpdCrXq8mmz/7KleyFsMxCj0tx/Hli1xEX/pAck
APANLts71xeS/jyo9gIrD2QLAh+PDNU1jpy1uvsf20H+TKQbVOmF/7MsIfshZeH1xgZX2RN4YNsQ
RjGrER3WiCrP+bIWwzlSRV4aeQ3ATrnHxoJEs1Ht0/wFHpVxa6N5K1X6LifhelVbFzGcGx1A+D6G
JJJ5GwrwEpM7enKeCJxWob3w+UGHBAr5NAryGs9zNocy4tN5slXVZJAbh8qQkWftzBxHuDBsPmyx
C3MEi0HLOsFsQiCdXFHZEw2eMbzt29f7n97OA/s5Ho89kDzMgxelQxMvreUdEq06gEOwm3OxtqwO
Zl8ZjL4n8HSmmD8jHuQcByEV9aQxCFKoIQXDbuAYBp2sDwAhDtx1lp534wL4ijm7kkJ3ET9lBxge
+tL3d9MMMPMfN8L1uKc1letJwouqBz5ZVUcrqFLoC+rGZGpCcffT6iUfFtfj8dmuavGFV+MCSzzm
o6mJ7k4asuFagx0Hf2CNp2lIvo8vxJFYrnZuF9LTSgsy82wYDN2jSeBVrxjrxVngg1r+kLdaVw7m
Ubb1NTREiRCNvLbkHMRMUfi1bUurDhES7tj5bxW8xPd46kIhZBk+eGitFs9Dr69jCPpw3DcTGDHd
BizDR9kHgKMiFr9ysiOzRrbTm3Gs1D4VF/L0F3SVeY2UqWhbNP04ES49Lug9il2SbSGYdYA/UE5E
5HvD3tPSxeb9+KbypIP5xwXKvjYl74MUX0+5EQ/bgxGLqBPUNwYzYv4P9gZx9poTm7irOwsVxYaT
uLE1Ix7VVHet0cUf3/WRhIz3vG6+HPSkpwq0QD3AuBbBnNjhh8OBlEZCsXugzlxOLdpoSLwhMT5c
9xgacUWeEagkeD5pPqjAywarAyPHFwWyTSmE+eDyald+75662qiaiOw4swZuJx9OkLGm1UpkIQPI
oW7RWhLlePI0ojbCCDtZKTl96uZEBVlnoephHuDlrxId+m2HGWhwohp4mkSG6hHtCtKLlLRGVfzo
ui0MKX6OfBJlWQPMrWoR8CbqJygYLt5IXcoTmO4l7baHxsaAw4AltnlXl8iivaCWz46+WUyK14Zt
82FCfEA/gkaafMPFgrXd7RXnU7q8osHdCTo0Ls1a8VOqSJnKKEi+Qw2Il5Z/VRjrgpUIKeUcxcPR
djDyNbLhClYIzeJ3Xa5tP5mx/7Po0hywnlI0PfzGpehu+iDkVgJB1kpv/L1L2ZrefZ+J83Ava5bv
4kaypjHV2Bs0zYZmJQ+9rVLdd/8uLjkVE2ItOXQpUWgZ90nuA2yUJbmH1y5663F2NHEXtyKWoT9/
eZei/1xUEii4kkJ/yVnHDnSX4Ml8gU4h28caXbUhejqwnyRzNb42lJyRhN0sVyqx2ojzQodNTgvS
D0cEdhxoDRQxQ5LeB42LD6yEs/DDZyTwx2JDsyLArfwGnAOx8JPovKFjUS07o+nZPqGgfbjQFI7/
+vFucRKeG8+zxrG3rwAUNjCzsky/k8tRJbOPFqlGKKOFooNvl2j8V/FfFMJOOIhVy3cJ+dI9MRtU
1uhC1aqY8l0yp11SfhMO+kj41bbOZ/Yp6lwDJvtLN0vAkvca/vWhZtQazcuDEaUs2yrFfWAYmzKr
CCdVUoTTaLBkqckJo04vxscpssMQmTXzsqy8PfXDuBkX2YzcQ78EFfjFXaKUcAB7jfQ0RvT1u7DX
5faxVjbTiu7vKPY8Zo2nQulLz5ljjQPUK9GKfFz23oWEdJZ1klaUlwpchDfOCobWZXwx0LF1UGui
RH4S+o+zJCoORN3GZFSFEy+c79ow4yXK88Tnw70W4DTmdSsGn/n/Eer664s0UUVtI33sj/rUZiH9
vxSgiLtjJBKTtRorf/2YzQheedKz1Jv4H+6bvVHzekKvvqBw6O6/mStRVHlaAeCvYokM9i32oxgB
+0vqZrJFyl3WBsToPjN4ZImrX3JOraceM/Sjv/5whLV+vp5bDZxNZbogqsW3pbBJU5kzCDwlPwnl
SGMqMOZWbw48VVqxUUNTwYIHWB7aHEc9xfPwhCfl5YyVuie89ZD9MYO4+oDG9V9XirglCkVDHjO9
pH46YIk+aDcCKLGU75LgncAE3dMyODuWf/XQTG62TMFjLljhLD8dO8SRYH167eeTRVLZ8m0YArhW
8IaPSKHP5VorPpD5UEDPh6p2LYOHHdx+mJv1gru53seDJAKyJ/oF4MON1OQpCgKRXLazd+ufTA83
wdTMkT7wythvaqZf7zpYFwn6IuFZCs7vksd3/N7S+rP9USUoXl8PC7OeXL/oBRQarH7eb0BIDscz
iO1tAjutSeEf0Isv8YpUMab5dlDhMVVrOm1O3ffDbQ+QIvseLjTP0+5CxJZox+uRynAKwA1myLGK
BJnD/attlcrbcDErd6nh3JbznsYPrHPiJuE1lJYbflUdDG5zQ/TJTXMyKxI/2kQuX6amyIHaEHVe
s8MhJ/DQWCPDkqJre8/ryFViTbZ2h/3g4i9VWG564NT9p7ZPMvOusxAD+NSc6bpFsAgGJ9xkaf4M
D5P6Nxm7xuhr54fVkM5EpgRkgDfP0a7SQroM8ohx38OG1wObAgqwd1Fr+OTlGYE18hs5K0sE1bcp
M9C9si4RMXpj0SUzIKIYRYnqmlSZhlSJW/K5NSorfCJCBkqXQKtzMCpQIn7UowwKcN+mf/H0oa+y
Uy8SuarTggQgWyftcMtKsDHXzNaa6mdSG4G03iOUr0EWKE8w1FxyUaH8hiYhstHRZkG9J18OeG9H
D+XLroZ31PU+6qBO5b57wiNSV3/KIEPVp4QK+zepTxDVMaX0OKY5Gfjlh863Ztg/nIpMuE/gBN7m
`protect end_protected


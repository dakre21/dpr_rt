`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xa4gS6Qygv9YL88jzuMwNWswbRbOWc1dWV4F8EiQpYBiAQ7/N1F9T63QMmo0ZTFPtxfTsrMkVEZi
FE8FgzYLBw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oQ1sV+yn3W0auajcdR1vM3Cn8FL+JdkS0BVxqUZmygvdJRLEI2YnvRQ7X8nd+HOys6FuXeEB2KgC
H9oU1r2LOyLUW6BzuKCMatheNWfa6f5cI6prqxHjdVMeefHKClgSwbmrmuexpr0yBtZznD6MifBT
6kFg/LWySlIeKqROR48=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vf1nHQvGKyz1PRR8v/QKdiu1N5wfIwsHhJkh8KvUdcb84Mk+G/wK5QCI/TT82HD+GUoDUrgSdJ0G
1kAWOewbFD3YhRb3TKAnxMJMbRFXeo0pK8ptx5q7CpFllg+Kch1SOk8ot3sCr143YfUsy1AX5pQV
/I2Mg1tGj4xyz0AKtvMJTisabrDCauem4W/MnQAzvTA3RfpgXYMOqBB4oiAkEiZZK0n5sPvxu527
Nqi5sd4TW+Yc1d7FMBT6pDbGipyua4epwMXaBdXIg+KHKvV5ToUU5xrCxLELCyJ+jKeMaDI8wNai
A7S7eT3oW/0DuB7A1oy8ZsyK4wJP9FWNUjFFbw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KDyf8IWfSHQopdnS4IN+wFx/CVezVPQBXeOld/FGLuZyFQuxYTh1QnGArRPSFpOMHIfFgxcwyGoT
7zqU2L++z/Ig7DpNMbHjcKypukzq1xfMHCX71fpa+Qm30la37/pDBdGiCgJ1vPF3Dhb+l4whaKNw
JtzxgwZDy+47Y6Cpk8ClwqTsOfiFWhCTY5EwQekWNeZW5fTmg3gmS5JQzxNYYlLdVqO+nva5qso5
XYTLE5daJhBNTD7xjAYdZmR0q3vazpvnNxGgL5MMmrJP2/A+TR0DMsMqbWU4mib5HrDssm6m+u4N
kChpHD4fsv+S43LBLPnJTx0htYZ5GYR2XzXzpA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hd23RPm891CVWP9FxOzpidoPIVBu2VR+S46gpO/uGhDMitrCE9XO+JaI8PjzymvZaaGMsMOJeHPu
efzx1XrjrobGw+ggRnLDY20PdJ6UTW9+g8cUeX3Y7OTc3s6rb2pJ9y7Mk2CJGuMvMUaaN3apZ8cP
+zVemEP+oikm6nHHm3N3vqRQaoy0irEHsgbLTR2r+a+7P2CtOd0tlotPjuE4abnvwlTqCkfXRCxG
6HNGblDqeG3ed6vNEfd5pO/bpBqzr6D3IB4wZFfy/9FwmevPnWEQOdcARw47bF7OnYdHDv2Hvy1G
tsGQUCNMSlzskkjwKrWE452hLCpKl2Dk0Bjq5g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pnxcs996xjQBH34VxtXMCZhQj7UaTZWkmAnr7NXuav0DridpcN8OiguSlu1Bl9TbW518iEBPQYt8
brIPawdUoT9Q+2uptCLv75NWrLvmDXMliQ0FfGyCkqeTZBSKM9iM/Fry6He7xgyRFxSOyQmqBDxX
b4joeqPtIb1cVcIsZnk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A4LzLlvZdcbUdjoX/flZtFK/S7vDJpuHxvB+OT31syK+hajoL8qgSEHCzJAOfpgUNh2jnyjzn2d6
ZTpAVJNVpPjNzJBaBW9fYZmYI+IkmcU8IHiecQNcZL3P5q8kEUcxZhgGo2xSci6OiXrNs3BMcqZR
yPQwYdVxCczB92j6rrkjDwcim4UA+hFSpQ7VIagomI7u307RPLoHrio+B1co+DbuXQdXcoA0pWtZ
3bRcYGQJJ1uwtNchh2tvqEGJKNAoZR/M8Tn4X6O6pbU0nUyc1kMyxL3tgqbWwup3EJY82C/vMT0y
IxlIpMGmOTSehY4ruhsvraDp4aU9OfXqMP8kuQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 883216)
`protect data_block
eeabDO7HhHiD3DuVSXQc1S78LdHOCyYsDdFoh9/7KqViQhMvXzmgjZkO9rb0oTMK+yAaVY0OHuai
WZtjGMi6RbukNssPM06Dr6jNnlJiriFO37MiixIg7qDG1ffjzFdCbr394WpTQ+hqpYRLoNw52SHF
FNncZOw2Gr82H34rprpLVBJUXFD2oEPyjORQxKZNOgD4YpSd6BLFanfk8ZUBCufWl7vTXeC0IpBk
NjGd79RDmZkJySyqwXkcw7qslFYZCVReX97T6WHwwZsRblw5LwHAJHpkNhJVZ+5ROTuJRhH6VZsv
SJmqMOpL737BSAC5hAv6NK3Qo2xNcQkySHHItUSgvEpIXqfeKt5pC8Yty4RHpbJm1wFu5fqpI5MF
CFf3M2eaWH2LZtRaEI6wYU6r7PF9Q3Sx5yt5y5alf8/hwfoXgHteIEi+4FK3fdsT9jWtFBByWQBS
m9yk3xBXAhOkVSRybthrF4biNOPjwaDPEXrC3AKueEjilZJyl7bQUiWBlZnCAPICysiJWQnJ99bA
E0xIxyzBoyE1gCHLI2LfCMr9N1L/E0QIHcQb8lZu/K5pRRlob+fFFYq2smp9GiiII9v9ZJASqImw
ffWXoKs+pvzr3v5MB9lBTkz8CmlOvS/7h2ggIfkn7SY8HvfX7tuJVTxbpRdhMJDvvh0u4l9fALdN
oYIEiABE6UStjqMHT3JSU9fchYpZwYTtvb7ZQ9L+IYmFyysgUYwaVZTpKUeZ5JF6B0+uDE6pDYUx
w5yHzz2ARC7Zqw8RFRvzo5PgagPIyWUhjqw17Rq+svmI9E7dGz84GHFkMtk+Bxgq41x2pkFvyPWM
Pxfm0x6scSwgbgP79RZSKD5+iNO+Cyf4C5RIvaVjGXfLOzxqyk+bWi8HhCVhoNnm7MZF8upFn/Be
MSYX/Uum/Vfj9acKakUndvpx1zDkj1iv3+Y3dFyYEE7kQLSRNV+LlgzkhBhUhHHnFhMDDnyuSbwI
PIQdB4gY0ZfqcmZKRHJzxelJXzxfsGaHx9wAdzP9Dq1ud8GRrDBMsSInnfzuYKvoanshr4AtuZz8
Ad2qjmiQ5fErK6CekzOSRpfv4mh/RMd6yZ9Tzdf6E/3H2JkW8IPDvMLGhedwOPw/U0Y5M86NeXe5
IvMBmc93BqhJ2Eh+w+VU2VtheySm6WEboLwjL0AnpbugNA1YP7s0jv+nL4+wSy7JrjV5XLOeiyKy
es31OX5V79x711KNkNf+7AaMn2sS1L6HqXK/cqW6e/3bm2OiogSlu68avRc9OJE3f/uvqvKyfqgv
oFo3t4d7kh+C1mJqhXkGMiNzvq0RMoJqzfUpyXXZnfCPrqPHKaYacUzAmlQSOV76jfpAH9fYeMGz
YM1Xq5pU68Ocbw2oOuJi2oY12GZyYJWOJCdbP25HMzDg630StTAzZxc76ROzkqIH+KsLMjh18Ifx
jk6+xpJq6SFms916IlmgznvvEffGFl07CQ09xyk8AW6lyq6C9WEwUjsiG2rv8QAXC+1UOW57/2t0
a8KL8UxagDnr4fPzQ2htGdO0DrND4E6Eirtsb+MHApUX4JfJnKqTPstbGdfiKmH+qzIpsCYVY5jZ
4ZaHwLW3eIx5XB7Oz8e52IOoU8UYXYOt3EDXofDl0r+aehHCJUcG4d0D8GHzrqzxj7tMsUr39h+P
TCGr1CgvHPrtkoohlpeytRlhV/Ee1dBBibu2aRf3q2YYenuT17w7k6ejE0YxnOkm9OJck8v2N/AF
1pBlIeE8h7C2Q3FHZJlMLYoy2tbYUTQcjtStvJ1gtcowNMgdMYD9T/sdRCfp8PHfAYFVOtJDiIlT
6wK+cZPuUcLLPaXTV14PBgv2VakZeyzY8aoZbKnOkGesrIoJOsR4DEUslYdR5l/xCN+ngDwIBIdJ
SHejuy7mz91k3rZbGT0nDESwrkKBq0L4obXE4mJEcI6gVLdb8FSoi6WkaM+H5opUfLTNCy+aaYSH
xN16YJDbB0Q2kif+Lovo9QagK+P9W282ODDqGfBwRyq4A5Unt0udfhslvVQYqkCk71xW8DV5aQxS
gzLJzwCGT4H7fJJWL5hW7XVaPoKHZ+pT6j60JDG63O7EeS3sQTSRFtzrNzOuDBesFA9wiO1U7K+7
BXMFTNAXRyO3S6iZsfJo+834J9+q7uP/AN+OZqvyzufUpqXAkHGGhn+OHsYJdwVPnSaxjF0oV8k5
19IDHTZlHe2hoI6vBL3rtlmdPfj1K5WzNkP3fM93AGb/3dth+Pc/PCZNqo3Uuwae3ZWpfmlodqL9
xCBhjequAg4+ZWNw1bDuRZiKU/EEQcA24tpw9itEMDRy0qn96oqE78/ttAQOsAbJZ0TR5q0HVAEy
k7PFvPkwK6tlxvePkLAQ+gY5h9gAvEKQuVtMzYs42lyD93v1dQ/eLLOQP4T2lJx+jIucCUsyIa2K
uGH3tavuCkV+u+p1lkiYyxAN3lnJCdN0X5udexFaxvAMJ+z4fJEZ1r8yO/9GF/sw+tk6mIHNd9nv
SVN6thbChqgql8fkWjBXD7NV9GHhdqb6yH7QFvWvnDepwkAP+Foaz/UV1f7K5vWgh3bllkz1TEzH
3lV0oHbtLz4YFecNh0yaEqh1BaZjithLVcvdpBIIefoaFPApZg6DoUZEmZNV0hvnuHVwgyiiQakN
p5m07uEbM2ZaYJmxmuGeqSaZ5b5kaYCP0+bqvrERRwkGERt5x/y3zEoVJlYrn2+2jSz+02ZAJF00
Iq5ixnOdFcLsXW1YwIXOw1M4JUMKyWVNmpjzx33TG2H7gZV3bioSsR5WMyfxFSr/X0z1PhbOTgpl
6diANQSUTmt5e4wy2EN1oxAyiu0NNCB/zrZYS56uFFSgtBC2Oj73eikUEqdQ1h8doaLHGKoC1vkx
O3n9ZqOQwdjutEIO8AMRMuaM2K22UVH4idEJT1JjHDBLazRXtJn0O3JN3LYrZRkYlkKUFaBH2HeA
eaene67Q3xZi1UkeAA+VPGGgkD0aa3ezYHotgnJDsmCm5RSkQav+5cAKDsbUxtatUeCndrNeeIDd
dJZKjJgh9eolGTBJWuqmm//J5kVL6wSLyMbCvH0rWAl2jk2qY8CWGOepD8LmL0XBU2Ou81yIh84S
7u6lOHdziMOOzu/RXjXM8CfpRagSlyrGA7U/QgtDtlNMu/HkLqvLG/PsJ88Ayr37NZCgl8CA/Eup
F2HAHWGfn1icjTV/2CCwLh3CVCTjnxCqSHBLSLHePRxf9bCjLUcElML79mnrd9XH95moO+sHF20Z
Dmt9PdDw1miqIAtXDvKcKPndhh0fIr1XXubHHvBymD0kXPi8+eY8W3BbDbi+L0OKQ71TTYGHmM1Z
lBYvpXjwHoHNIrzSX1PzYQksePqF9eDVf5rTYDTXJCdZ1UGerqsOddfjdkefGWeaFOtoDokAca3X
E6uD3B3jmz+cEuf39AJVNzbW7SSCCJQoX2Ww/bXUjDVtnlAt27DqVMB6Ot+YrRL212G9FzYMYrrG
nKMGCJ4Z9wbHBzPfNltVJQZGfd1ocK9sAkp1KpLYsFzt9SE32oWRRqf+oohux2DR0KQbVYZtpu6t
psuse9sYnkFta7cuTRrBul4Qt67MTmTIfyGrb3FGRAOjHPvc5NZ0sGufqj/eduncP+7tKjHuivVA
3+Y8vqD/jAXlSSd9tCkjhLdjTju8LSbRoifDUDYtzj3yDrcpcx7gGdWMclapahNZI5jrZO9aU+C8
TkOp1bBBnxB7RS+fz8im4/mp50IkUUTxE+VjCvJU7DRPyGtUbtnegcaQWQCs+Pei891X4uQg/GhT
JQM0ROW9tlWI38sc58asrW6E74riO+AKASrzXNddZ1E7inud5kxPjVgr0hbXSFNBh4odpm4ZGp6H
CbYklkKbGyGwiW44J5Q6UsOGZruzdAMprrhxMhiU2j7n9nUv+bPHbjOykym3tm9qTuhTSkogQJP2
W2R5MutyeVq0nQHhhd8TZLpONLvUrYzxKVe0jjCWFljS76dmrtfhiSQroHWrC7842pMFsrLjyUQi
Le8qMq8fmlLnU/5ynDPWpofMOLTOq/dvwP2jp8mokWtYw7tiEZ8SbTvVYX+50TZhwWgbIHSfuUom
rcz6gzU7VFhPp8YWVk5UkyeJzOPI3oapwgBAb9YUxCcsiwERkKDcJKBiLTmY0uc4n95tgNd8Xuv3
ctQNcMRxnQOEbo7jeDtfahUPGbf6QA3XW6dFm7O5Qd4WoAJEPoBEUYPPcgc3eUYOjZHf8Bd75eKK
IEfFegbVI6nlHj+yjaFBDV2x0muIMhwPI4LEjsu3CMfPBENrDTBYq1Obl0OblSVMLIlqKxT274hm
keC35Nb77KQ+DQ2cp/G7HRzhylYE2zkX1NzzQWfj8JdrBXRQR8u+aNvCcJHJKI+yhxOYP0qR3Uci
bYDxmBlrH0e5BVqVih1v8mNgvL23SmYf1Hvi/sRvrzwggYfeA+NUgcywqxBQwtgxgoJNvPt+w//9
g97t2CMnLXqY9Fe4haSMCFZhUJUJXQlqu1uXehr/ZiGhZgYmSoKij7GqSoDWBfBYNeX8BvQyGWvk
V2c+ztSrC/lPEIG009eDtp8Yy1AW0rC94C30hQYl7plFjJuXJRivXN2butELVOCklON1xoiJF27P
LsjxT9YATIj41NMo9En16uueFL0mvXNaFz65OdhtxQur4mr90/PL20NtvcFEI1dhb9kpJMOP6Bcd
BQhiUy5Y25AiIH8qUgHBXfMcmAitUSXmCp7gLyZNGwVpMFVYB4AGKsILJv1CIEzRzdFWkL6PrRjY
MOEalp5bpLk8XKs/AJWUceFvRo4Zvixcm/YDTGEfKsPBRlCtOoqnLmM0ndIvS4flOufxep1gvmFG
6tkHrQHJ4FvdHXRrvqqIa7QNmEmypJLj3Pc/XZ/+vzVVVsM2GEAFJJ9R0sOvjMgVvEYSE16A7D6z
g1IOEkIHm2h1ah40IKaFh430q3szhAQL6rh5n9eS3ra6IgnKxNSONFRuFeQxLJz+WrgPDxduzle7
2t30aSM5KpvIy0SkuEZgvyTky4rqzuQ4eZuKurU7Dt03O6cmO2PCesgIR02vYSgyS9d1iWYb6pSn
qtJQZlQ1ptVSg8RwWG//j56b4WywLUVFOmO9GtMtPu21z6sXVLapCnW6NsHHEJmGQhJF/xWdeuvb
0mczPHZTj/QUy1OxZUkpZX3vmi40dEzO1cIU5C1yI5mNFJyQf/dJnYbeSV9zABriI4N61aiaKtSx
qcOrfLP36Heu/aM2mEJf5zL3sgQ+jKU/UsdezRJMGH9Uh6tgw45A2cIh8DclqgaDbV22m2z+FuhZ
rP5NibMKzywjBcq1chjntwLd2CaijqxpClnd3MoGZPw8YKuXGdYPv7yCOtnabZK4dJcojga3FzNI
fd7wDe6IYy9kqDrrqliDjpfUyQeykn4IS7HRZSg1HoB5/V/SiP9wwI7AZas+qwmoVIMh9hisz5JC
XOFFrwUEUlMas+TkKXMEGdDAIWP0UCJ7ic+K8xWu/WSBNMUKPVeVEfrpvNv+3QWMbolGVuPqf/hf
jVwh/HCAGDrl/jK84NJt4I3s3FagDGP9MYzx4VnBAzgiv2fMWiZi74G3AXenRqJFbHmQ9RPU7gTL
K8l8Pq0ARl/l26uWh1c0D/WHqgTkR/VI1CFm4HbJwPC7NXPV/kXljPUeIoWpqTRQyXAyMoaBFJyC
wwmi0l032xb9ktbafWLWXE5B9OHTgwLDfmTNKKDYWVJagLiGEkfTF/QK/3cG0lmNAS/DI1d/ANXk
T+672eeKdTAZKGBX/GI58BGxIHlebSGT1fx0SWWj7Nql7++6wVDPXSVTjK4C+PGl0unzFdrSrE3W
odO0pYlgSFLcRh2ek15rmRSsuIEQehUpTG72SQE5bB6o1uU1ny6vAEKK8qjBiAzgRFljXr7G/hPQ
Yk3WzaxjCYw7BP7edKNA3S/ZMU51pNnK23eFp0Z2Alksa4+ld8qMNXhcNBw50mDYlyQH7yAceHEg
+h4axLC0nbz3JHvDYwQWqlEdXohhXn/4g9o8n7PTHDIXE4ZxyGV55apo12B6G1WAiyVps3NLPFS5
Dqj7NwkRJ8ejNM6dKJy3DCrFql/8WCBU+73SRaEdWcITAKg2RgWjoKkOcNQ1aXRiGV0ybkmG3ct4
90eacZl5T0E90qbnK3vFM6uie6a1sz+vGZp825xd0dOSxDa4SHpT3RkXFBSQtmHbkw7D1ZElf+UW
p6W2/ebjvkFxu/E9XjdmpHu5o0C3LsRvURb4lLLadBLX8nh7u4JPINnpesnZbHF5G3FvD5RZPP3s
vl1KWgPXNTHY9BuJ7IZCagEEHg2bE26ViaVgiH6r9FtRLE2mIHQ5ui4Bph+KpaBkcKnSr7TJpfn0
NsO5a1jKQaIAXBx0Z47bkOsUIOpQoI/F8byHjOtSIEEA9PdqJYeIVY4USZA4+vKi5H0cZ2l1q8mm
slzvSPL3Z0Wo65relRj8D7qFmptLvD75mK6ZyibA9sPLaTK1RD+Jj5H5lWVWqutYQ5jY/+jmc39+
9FG+JI0RaZchMwmpudUmfG7RhTQVeoON9aWEOHXB7suw8XnVC0OFk9UBpZ1nncmhasdIwELy6vAV
Zs/RsDk+LICyxAabMDrzS344NKDjTCVKbTI9Y+lzX0cs30qoLBc+Ind6t1aViKDPfrHYGavxvrLN
PhY3oigKNSX2Dd+rKx7+Xe8OR000A+lIX4bSZ95CcUryzVa/xnaAKR/8yr4EPQ6xZ0vQvvGnGuFs
0SjazfhYAgMD/GPiPSpOx9HDpqezGinCYidy5Jz2dG2Ykwig4oX+9WHHKx0p/dGjZjIwKwC8AcNa
mKMMce+iorRUP8Lrlq37i+V0+yLS7UebPoWk+LCvBnkFCNtLxzAASwZfJp60edtI+z3BUoZJs3nN
dwwsIU9ZKbn70JXkSvzEF70/46/O946CDe3h3nniLEiQPpN2/jF/iplHLae92xYv+1wogetiX02O
9/PRkNpGvSJ6RoVc0PteHhxRftzROZpen8wMpetQBavSnM1CAZG2P1MtMQb1rWl93gUnWoI+aDjI
2NbI+4t49zEp/cX29/yviw+JDnKi8SeWMVec3IJNgGEwSRuWPkXyI4R1IeV7YeCfS1V6MefU9rzy
4i8ar3U/PwmTlGLq9BIeG8qFHKpT3WOyaSBw5pp2eRJNfzvfX002Bk91h2fsVbCUhs77ga+nhOnt
jz0NBhy/GN0J3h4AfM5HhF4StB0MfaPJzkBtEo94nAs4ltafR4JI1UKornBM2tMbtuHKz4yAjXIg
Hfx133Qv54U0+I1fhAZwL3npEqHv1tzRhUqY0e3kIE6/yI389TPk8vRZmD/gUYknNdWu2wRXs1f2
FoSNRrLA4I/M7+K7q4Ha5nUtcFxI3/M00vSU0jLL3Jz+L8dDfqzly/osV4H1ZhM3SYw/IfpysxBC
K/mAJuiypvNPX/ionHcD6+s/f5pHbfp99DdVAOm9FdfxdYEOer4M399fk/UQSU88Ba0oizz8qA/8
o5SoT1yPScLBy7A1m4qsuOWafJEwAOpjzqj6DuofVj4jx43XtltPZ/4jNp2A/eRcNanh6+7OMJmi
OObRnX1G1BxOmYyyuAaLFfEOADWcP1QvmtgZeWD3kICYW45hsT0iO6Bff8MDqi6u1AY7tHsH2Rn6
LeH/JE4c0AYXA8mYaqBcO9BzPtOR2Jujx2ThJlUShODqJfLSFrO+Q/CDWfc0y8QhObmaQP4/XExg
EwIzBD584XL1mDHEJbCkY4TTMZiVK+DNE8hbtofC9Gb5GGM97vAncP50m3WYtEjm4VAo+3Ffc/o7
Hi9/Dyt3Kv9Jc11WchdPcO7SCVcb8yVZIzyHVmwXJiYN7zLAPhDvB4U94UmJIk1jg9MksiP+2mOw
waqt/03R9K5gPdPM0sKkg6VNK5y0IZIU8Ofaj+dhxYu74p5c3QGPi259cy3czah900gjzqiT8DxJ
OC65ykx2Wt85L3ygq2ZhdTC7b0M95Wy0rrfzex5IfJfGbrLNyDG2PW7bX6ghPfPCeT5PspooKrVu
8jP5Y8S+20u0x0m26s4wivKL4s85IDX288CYMLgyb2gxoOIh3L4p9zrDqx9v1YnuEpEcae/9I0IZ
8dxRhK0vObX3sRqX396W8A6g2rdgr9isr3gfDs8eZOpdeJsFZr1tTOUTsA/+FJV8vDY80FPtvZLg
Nwx6kbSTyvn+mKYKJ2bD7ZW6JXCKkzGr2rcxf+sit1FgqSEsLYNxXUEDNDZCBto2eGM249n3l8nY
k+nasmqLokHcBen/lr8EI6hfbx9wAl7eyUuZjzoyrmQyK9RexSABGEGmAagBs9wAe5wqLCpJCFBQ
diLatQOwDV10p6q8e+n1XrOoqnc0A9Vkgg0eabhiXqxcXfN+MAmyVoO0gfVxDVAv6QY/xjKBDpMr
pcU5XLP53ZDDXd2vQFJen9VbziPTFryyoolqkrfIxj9B7axM1GOgUPPGaNMZY0V7auvEuwZTPoXk
izUZ9w3HXh4y0qO8ir86RQGlwsxTwr4bpf4IKM1Yo6dGKhQITxKFIZLBI4LeFqZUI54Hyknzr06o
QX/zOUW5yFTwAWcKyv7se2FQad2haRfmYFRV+nnPISGtQN+c5+UTR2UYR0JxawkO1sQ73nTOlI21
T1105uQhXo2cVh5X8F44gvslyoFpzOowApl7oM/D3VJNHaXKpsTbfYq9KcTgGofe12HnOJoW32Fy
mFF/V5pQdnQ3ARQdialr4OiJmLHCjAXcxkINaf1inLS1/USyiHpFU4pNg/gjy+eZjXzwWRf1Ka/o
Fj92kjsDxGeSNiMRkORfPltVtLeQ0H0l2TzPdcyypNLRdHcnWlKVzWoWsx+QVpISN9LEkr8N8s8Y
i3iTwoVegMYA3jue3CELM1qlSfQmUrkqrJIbuHg33eWZaw305s7GgXbPQeTNnhYavMyn9Gq4X/A4
Drsm2t9Hl/3HiXEBshVQ6d1xn7cYle5CJ6Mq2V4GRjo8ad8pxiI53P1YIiyP1rlUbmeey+fAtPgV
3uTU89U4U1Tb71+qCjQVZXKMSr9S57nQ1OtFB56Ucox3lZJZAjl41O4WeIVbN+orsLnhcm1/RvD0
3Biqsz0nCedqNEP6akRf7NFvNI83pC6h1CuyPjKDelz68OT20Ho4dqsTnFuDiHPPTGeiuuQgKVBw
x4OQMNOpf0jFr6cR1OJ2axQutRef2/YMkjViOUrDEvSafahUi7f6sbYlsi8bJ0UeDTULIWdN4iUD
5QGApZYOeiVvP2IYnVX+fUHgsKxfAaEgQvmqHOi9Jd1xFLM79z2kjNGHx+wAe2PTLK2LqSOPzQth
GA/HCifptogTct5u5v0jXbPaJNFt4hIyy6LFNP4gyTcZarspkfQ9pVfC5+Xln6XhK+fa3e0NnHUF
gPVCc8yuv3EibkaoIbm/bib0Yn8dLuzPm6vZwYOeIOQvVHvaWaXnCRQGqPrbid3nINPPEVteXYoh
HgogvTUIF8F6xS5CdeSzpgy5HM1vEfMhMf7iXwSIL6ZIbCuQFmyBNmWJoi27gTIEKFkBtrVn8lgk
qr51xSwS5LZHU+CAz0X/z7Oxhziuwa9ePASzpihCI8e6eX1y51is5+BHFRx9D7mOcitVqTDCkaYf
i7Q4yva15KENREC/ibT0C/dg9evwUcG1THc2V0G1IkrGRosrnNKXpicIqKJqrIEaTxy45hpqM8j+
n8Revx/JDW4Ow/Mt+U8G9U7lLaHQ833VIPbklkiWpKx01uiVzBbAJiEzevUS2GCSV19Q/ntvIScT
jxKb5M0Bc4RVXjUOi3Hp51nMhhKDZDdnLUg+2RxRvHeQlihYtY/7ZvTIsOft5x7Q9EYcR6x3M5o5
ECA4p4NLvqYnPSUmIF+Yj0kXiRK/Y7YdvZnPB0Z3F4FQUJRsenRE4hfF6Csf+2Is41ZOeANI3bJT
qR/YWgM5ubvDbSh2gOuzrAc63UPhzGLPdm+peLbtoj2ckR9ZLUOEzFGXhMsw2e7eoTl1cOXqiAz4
lQ2YB1oY4tml12Oa0ef/o1pWi24kNZ4VgKS7mlXhhTbvl2yQ4dHVK7pFv8/ddW7zwYrQrs5gcRx0
Qceml8V9cy23o+I4T9f7OJFOak/uhhiA/PCfSqdtmV7cp0diXqEeB0uZcme4gELrlBkZP9ncxVd0
AY/1COlQQERJRdbMEW49S+OvD2R+wot46MeLtF4FukYMDUXl2lxpHUREDf9WZTxYuCUS7eTmijko
criUJ1cWNSgrPa6HIU2HVuVM+CgBm0nIOJOIiqaZU6Sd2C/Nz8dgARRtmHEOSTUKSb/e6g0Ew9D9
18DfCvQ7jsfdmfFY+/bMjbDQ3m0KnwCo0vJuIWYjeKMhAywI/JaWkFo99R1mvCNi+E6ADmBQLsau
aGBsgdcFxkr6Xosd1//2c2NZlSkZxitM/h+CHIWnefms1EanyZaxAaj38LH3TDowPaQhYGzQELnd
Ni/4SBursEjN7vFkK1CXUp1Ehu/uN2/aWkXpAcmi4Io0ApbivBTikE+IlArLT2GaUgzr6bIbo267
+KCPD8E+Paa4BBrcm6H1LL9rabdppkeAKYqIT6/ORO7AInD6RkWUdauPK//cHElyVeUiisL6lygf
mSe45WxWy3aWsVZsBghyvbh2cCF9u28HhauwSberhCKW6e4DD6h/GT9G9wvBmGc1aBDEbk3slQak
168+dHyf9AnavBqMPUrresA+89VMVLgCr0aQwgtGc8ykmLzBam7uS2nq5hvlydaEDdspqEMQbHjR
BcpHL2IUZI7tdbVdngCfnNzCudG7y/it0GyTw4PCEqNKtv6lIplO4wlBs6nWuYv7txngmbOJvInw
OUEvOd3hP0U0K2lu9205vIz9QrAEOMFE8Kbai/Kw1SB9NplcARsKAs0ZKLYl9QKT/jS/SoYhINsF
ofIw505bA3oPpTVTV5N+tMeu/Udhs+TfWdI7offHYK/r+HzWoGaiXXI4wc6oXzRRC3IgaOjkPSFL
K1PWdbkgTZRwBNizyT/xXJLxeQQDNQXNUm/qFDrqh7IvCB9ovVZZwc0w/OQyurk6ZsMYVIef4PZY
24HNilirSAuBS7Fr/Qo/wE8NGSf9TKDp2cJohe8ieMe/gKV0ha+gzYmpKufkmxeRkNC7h4V8Vdhi
BrmsAKvPD7Wi7lvBM4lRCLJuTUpX/wmm041zkeG89jdFG/+Q9elE0xrcU7BqoUCvnZi3gfxog/Ea
1U8Vef9c+HuIt8G81dRaygTRGxNBaqfPVRgEZ0LpKSwcyiLPylzpGeOsBkaUXGcRzQrrmmjtuY4x
PLV3MrAuCdtPsKN3GwSOp22k2qU/rvU0qIWGa1UQmh/R2aCXGLLtO5X5GYgzCjOW4gxR0y3v+Y46
bmTeZXdUBuQHt1WXqh7LRStTBtbzZdNTJT08YIDVXKS91oxPm52Esv63WvQuURmpUIQq6PPmqLB+
mxv7m5N8+KaVGnpP/ELgOcNgfWk7gw2sYkVdvCuKY3svv9yKwyEOiDgAkbTA4hRAzUss4mnxWoxI
3BpamCG3sJhHs2dMWjSlL2ncEBaEJPcHy643CtR0Rezc9w6hbDveo6pl9Dgnpl5+DPeXms/nF8P1
8QotnGzAMmeeivyRFhzsgNzQP04qwdFARi2109bvz/XY37KcVucNaIIB06yM9M7QQINHmUcqCvn+
QNm6hRA+NTSemJXtWtJn0o9mn42+j2mJFyGF55pICB58CB7HoWLhdCKVcv0YB7p7eAaiL79PD9rd
QTzecJ34pn0fUa3S5TwtcLjVHn+jCXMdYTFo8YRr5G8ubpNCPV4KRFQGxOtmpK393n3o0kLChB5O
Wp4b/2BECA9MdccKAz0IbCe+oMDRh+ecH9WeKNxT1kgdCrCeXLxER9KuG2hINfaSVzH7qe/1GVfl
5HFQPzqw6WQzqtGmnpAczruAxlmZntSAaH76zmA+8nbDmMna3Xm6cDsyoCyaO5vgx0mZ3n+nDH3Q
hGv8nGk0hUuT2+gpSE9sKyZZOw3zUAZkKhfWKkffqBBnAMnLc/LJcksEH18USg96OVkDI/zuvYja
UfEC+zqlQQw42qACOeTmOLW4bHKTr3aaRQo1MIMAuqP02ZE+DhH767f8iuJTpASik7Ay/vDe+o5b
5PSaObgu8SoTCixWxveEfFc1O8VFWMPostSp9ARdDIi9diQtChahHO99uB2aQwY1zz8RjVqoETAg
6iW3PrHsv90AQIbTXPYvseZi0ncyId7/HNtWdvl8xiETv071KV8O96KAKQ+5aqhoiclzrbZdUrm7
3wiopifF7Ixhp1BvrY3KY5AKOX8pZoTohzRJd4Tc3R6Bc8u3OwkkFgL7fXFX7iTe5JgVjbiBZ+G2
JxrVR9imLzIO+S06BiLSnZT6CNcb5IfgDikQwOMT3R6QoToChJq0607Iq7qvzr1H+NkSfnzvAWOr
FOKIXi2Bwd0yoJ/inqqwxjJc1ByzDE+IRhFa6oa2MBN+RmA9v1sC2k9MDH0i1zU52epllwiRLqN4
Hq3Lijxez4rYgQvMrpKGi/z4NViVKgVQ2NF7mtDlOcs+H1Fb2ZX2emE1rbzY5yiW3awGIdtuZeKj
itUG3rNjG1sgIrKy9jQjQbdhRWLicNAGaWdEqstZ1xjg80Apmw3FgZML+EGvVJA6XmEyC+e9PDmI
r3FVW87RET/lDkVSuD16/ZgeKgXIOM+PBdz75NB8erbO/Yx4qg6SYuz3PQeqHQlmjTALXZT/T5Sl
xEAqNeR/UEjHCswETs9CIGcPRfM5sCvItQ2zyMKr8ryjqUR6ffnnfXCyor8IKD5DVMjJfY6Qq6PR
pjSfHOdSxzeLQcZtPJy9dGBrXftczVQJfwEzD+dKzrKv2s/9GnE+Ubn4ajqOUSMrKyrtodp8uHRp
iVtzhxUhu9dK8Qb4c9Gk4qpBpu2z6b0pch5lOREhSOG0uTCr/STb9YZdZvItmZ2hfOz59A7fgBPl
JFFWssAHkiYhm4TjnYCRVi+KQg8Tj45CltUX71e1/SKgpB9IyFXR5rg0spuv/cj+G2Guxy7OKbue
xPp9BmYX77LS8KvVXj3PpkcXDrN5rDE00noCKcYpH0oQdN9KvYg13X/fMcLH2/82JAhWhH6kMqP/
dSHiiHs8ytx6P8mgO4GP2+fhSgYNHnglzERrBXufBOSdD/Jqoy3NyxC0+VnpCCsz9+wAS4YfEomK
CkKYs3JBM8mVrHHZarjCGIbEWDRKkzsRQzmchvGk0hzoaaKRzedg2yElT0xwJCFZ959d31Vy2s8G
dwqTqEx9q3YHlozQ+pr0SmQMpjijTToWJgGsEdInYugOLaOgtGqisZaHl8OmULtQzR/TanQyqT+2
racodtJcd5XUPQbugHap9qfV7oyDWSApLFFSUCgdBChy+9RHl4jO8DN9fI0ETIcGUGgCaKkffne4
NjkB3rCLwdkNMyeOCfXjMA3z61ADZNAjCI0IcjD2I6oTlTY7E7vfZJbOIctY0OoTe32wbfAD/5am
bKuciCx1Y5gfzx5up/2hZ8hnP0iHDPA4Sz93M16Qk50eSd1hLeB/hQXNzxWvPhnk3x4bIL9sn6jL
gFhS/RskMRjGdnbdUjKU6TLD5Y9WOs8PieXMYBsof2XKzhc0t7LUukIJcStxmH2b01vmsmCP5ND+
izWPqJdX5ZE57KNmefrDxzsH6Puh0wEEl3PCxfShjOP3X+x/LzaxPwEPoP5bqz9ldlXhIPfdvhCu
EqZEjFKdhZUxaqqsTv10+x5GljrozMkMuZYKPAUZfqkthozf6eeMQvgDxdDdLT59uPEs/Zpl07A+
ZvefD2piREOuI61ebXXqfwwxKa6WtfyKmjq0AwJ2tYOY2d0sHB5GNoRzqOhMQCVtqSuwTkUDPCAz
ZxQRIbJzOnxDePvHo2zwwcK68nph0Vv9n2w88EBozA2TeRyZsuqHhZPGTgfnP7nxsTmUhUvltrPA
xpeJcOkV/j1JJU7nuTGu7Ono0MpLaFTwFTdGWjw5ZWFB2qV0e6L0LRM3QYeWhxUCyk/I3cLkb3Oq
P4yuiK+BuZycfPJtBoRHJpwDzUIQ7zjO6K2DBS3f2ppKXe9v8RuinMp6YPKsSF8EUkxKP9S9rSKC
yOaJJyKLsx2HU250XQ/Q0Vzv4MeEddOiYw6oOirgEmqOMO69MjB+mJqH2JIGbUgsP13uLlsWgoG2
bNTqSdoFi9lumgi5VVor34YLZhLaWQWaJKSCIbV6QjFJgwZPcSZ0i1a9y7UxslBU1tRr4QzTvzVp
0VF8YM+HYX9i0/YOpOQ+f2BJKhJzsmGg9I/eB4B25IH9MItgD4aumJ3C4GIMqfzHfxmIygQeIvq2
+RGoG+ph4Ls6+V1Z2gMnR2QocFoAHTgJIfW1xyi+Kud/KoPby26cq+JossIdqsuVC1JUwr9KuEgd
RSJnG4wydBLDt7ZeXuOeEglkakqlUguSs3FAhleFBpnXizSjBiWOQ+F8By/MAWqeNc1qoB7dVg/h
mjpwHO+xsu0FoMEsd17rOv8Kcbtg58UNr6lIyY9uuuhGzv072/7umJ0hzE3nkxHXREP2MiS1Fsxg
/uhaIdkKMo/GkuCN6Gn/kzFSvJsz1bmCCJH0h05/OB0FVX5A7QECI9njOahRtE5ScUveZMMmBxce
4x5B9M+Tu7BgTKxwg7vDgTM8M14rGA9xDfWf6X3GOlgpoRXfr+jaTs1LfXlJOtTfQDh+m3IGBBkA
1KHgWx0ODZRhYQyZz1tQdwGtkZQqVpXOQU0Ci8vUiAqC1jq/9JQYlU07Vm1A9L2+EdFl6G68LSS8
8VJWmKTWn/lY6btaLZLaU/96eb0H4yRtF5VlcJ1gDgil4yv0yn+v5wWVqJb7TcPCsP3iNhRixY7v
cExisuDYutW9YY+CDr/HpyLZEqtD9AG5TFHTYXJfbq5KpBtShOEIk7txIJQRuICwm7qUubTe5ZLU
yG/QqMFZN9emnM3y+sQozq6H1jM7Ler3yq80dUwJ6r5dam9q/gClWTcc17/xO8kOO5X3qCL0gBD5
l6iawRRK13VPf3hoZMtw7QIfvLj1oaMfMRLQ8FYEnqJ9edCeFe7YZ07rmAeUK1vgR9lU8Q22JnNA
cbn6AoKeYjzidcb1Px2jT0d7PEOa8E0kDpUbbLKgtMrg5iSl/Q77wkLs0Gn3JPZ/19hOg5cueqSs
FPD+RvpBTdnx+8bvsb/ALiI7uYY5ah6d41HMJKZ9ZSdigg1yWbfjyZNBC4OpH67Ih7kuCu3YUzoY
+FaDk9iZ+YEY5ao/9zvrn1AOgRgmJGvwPskuSwfMze1GtTJIMbhL6o+JiogoxQjgsay06/VsaBjj
osw8rWuYbRrfjLgwi85Ko8Hz+9ln/MnbbYC1dVFWyFUVqM2w/jFsverNSsCY/BtHoyM5lphGsfvU
XUdtZrkiocaOB84BOxW6874Ee/K0oZuUEzKQeLmgrXqEvftqIlq0GFLh4fxWnJ05U63MIlgCwVjm
yRz5zZuX33CAVIBcOhrM4uTlRCW1CHgkClSuxPN2ryogsZbLqSZvdGJ2ZctrpZF8dU2e8sXyNc5t
tYVWYG0gLQDq/5yy7jKX3oth9+zgvhZNkxmq6EB3B2UdjGyMzBOrp3I8ZjXsU6dW12ATL1l+3yMY
hsXcTbJC/l57PyqgaofnUa//IpydLkbti2gTtIk3su2gdIqphrYdlrr82VFxWdZhM/IoNmqUm1tS
zit56AkYE0gGwAv+I5o7LFWmqQcMjsznbzSsFFrTxFrjPcVELyT8DdFyfpNy6Ox6iZ4xJUq5boh9
vSzZ5d1IurlhwqgioANP4HSpzYhk8hLgB8/cfBsqtErjzUhutUc7f03FhrJa2bLFd+fP3d8rTkeJ
q/CQF3KPMIxrisgw4d5UP4veIDtXEEgX11B5ZruJNmrE1I6PTE/qXNkHuidDpj8ps4iiqHYdfWUK
UgD/YRdCV9vtOAcJFF7jHdQg6esZHVFQW2ULvPv7YM9iMnIz7KcLr2fitZdrDdZmS3UONypq08Hh
vE+G4SxgkWxznKGrn+MpzqBz9O1H4ni7UUuAo64uO6XP5gzrlpglNa5qF7EYji1PAXyFGGHlxnsJ
pQ6oZi6S46OSB4V0b1h8qeIKZG9aG8HfNn5McEnVlss7Oh92JzkcxUyGbg9n9QkZf5p1nvWO9e77
TgD+rXmIpORKOvBx8k11dIKW/SgsQeBXxcvBh9ztHkSkVdwsRvSg4XXAITVgZv4q59+vrngleUWt
HT2t/hxviM/0S+ucr0TaMe9aK8kc/OtyZ811oLpzTQ8aywciQCTlzh5Lm3rgGM4KIu/uRXsWpLqB
bylQbxzQC0pW7ET6yb7N90SaRHRIF6FR/jNEnuo7yS5JaWTTkh+h++SIFINjooiGWG1Bppn1Kg2Z
7o3prlVMMgT4qiHooawCK9TGe9j0ubuIvaONdItT7VUkVsuLwMMIaF8GOyU3oqB5WZ3HzXNkGgfy
E/28SJqNLlHeLODn4l/A2BN98aMuZoFjXXu5SMGvGlpfTHGJrNl0JT6XM7dZgpui8ssudWzj0ayg
z1UGHvqV7OCbgq4OZcwuXinbRlXEIwEFHHDG9uoYWa+Z41pMqqr3xTWrBeINQSbkPkkCHywRGB8l
wuan4uNIWONg9cVeqK4lAoSBrF7ooFefLeye5NEG5MCYblMMOLFUniG7RYlThBSfGTNr2apzRYHf
nweTUfU6caM92+fwQipLJfztoKoPeWSMVImBR/UvlnOsRnqZIm0VEOUwahzOPE1ReiWf5RPbS5qQ
ukjFhi2oJdIFREc0STY5iGlJMfUkZERUGRTO0bY1/zt+LEZinvWzT1nULIWKqFPzmRAhDPpufmZB
6rvFfc3bJFJkilgP4ZVroXHeGW+LC80utVr7ljBKB+7DaxuSxcKbBO9A22q5vjKC2x/46MVOdLwm
t5uBPkXXV6dKT8wTHDNiECgtUIrADninwH0pJACdXnLlYV0C/mvTN2G5G14AFg0Jy0F3GDMuFKPn
oyj7PypCgMeqyhJ7CuB0tkT0dlY9SGyCS27yglI5gcsXiM6YtHZhCnmcbvDlVPh5xdukVyLgimfQ
fyj1bnW9QhmB5srog8AadQwUpT0cJIkj4UfMvnb/BDdCUmaYIyEN1lJLEVBwyJqQds5oZhYMbyDJ
MS+U3y+3x2Az7lMzrWLcgFsR0x6VZleydQH2x7dDiSkaOrnm7Y9CQexN4EfEqu7RlL/+WiozK7KU
8W7VF90gbQ+gNVOyTMvU83HsnlLOMMtdl4I06maqNAWXqLR0f7gc+uob6BOCRpCuWcii+5G/c0Wm
37sEa9/GnK4e+tjZBjTUK4Iu5A3lXVe3PjolCHQ9hXnFIc3L93kCNVvY6MPatDEwv1hyFqkCVNCT
kBDjzKF5+zk0J+Vf3qPy58i0Ai8DHVKw88Bc2W/g3x8iQ5cco0Biei0petohEfL8vErGD2pHQ4Ak
Pk5cM3XuUHifKD1IsJ6KafgkwLI2OK8yfk4D5LYQ8HJVQ3nMHizKdBrGLya3oegF8fLBPkBen6+K
rnaTTprOVWclxdGi5q8HlDP03AILLEQVHT9eACRnzJM14HtbaLbtOHpHS8ZALa0St0kMReK/ISzj
HRKDHOpvAfBaP7ExkiehBeZKMLc+ef29hXZPJJXLHipGV4qHkvWs9E5H3qIICL1Nee5E0m81zAA3
KtySj8qedDEPGR8bVueaVApD4zv7+KmkNW3PAFIYKn6fxs1/S9kz3S3kqrbVtMGeSnY9frbWqwAi
ALcPkWbg+oSF3v0Znnx9PoKu1xD+bgFwKomj2a7v22hHUt8QIE8ZhF8n68aj923fKLce7WOJE3Gn
+MMUOxAYVnGPZr9ChylpZOXePDUJ3gE/T8q9wyfqUmtiJ4uXX1vXNyM+CP16reByScoOPY61g1uc
72T82E6bEkYoe/clEfStTiFXAbwQChJYYCJ7sJ7Z2IUTZQ/QzGrt4FWXuznIrUBmc8zpnNU3gAL/
m2V7GqHra5wAWhrvQMkT5eaBfQsRAiPFm+XU6gCx6joaO5cljJ7VnmU635S1L9LTVsb1ISno7u6v
vSFcnrfJNV+T08kMg9qgS65fkU1fPic62ZUmMqwL9FdWHfb7cA6/uT6DxJGddsqSafcgj08iDpm0
xic8j//1kLD0830DZTqfQmDpLqwhMPINGOcpmZh2K11YRhM8sOESq3dICKfE9uxw2cM81kxhGZeQ
TtxENMzBx+R5kWtMeRiUNUAEFSbwWWLHcmOlRZbdtzeX9Lmd6QsWoGTzMEfroVJE2X9dWlq4Q4vV
WB2LZA1Qw/fIr94oJJHT64JRNL4SkTD3okfLAxDiIhDDlyLlvOoyVujKkBTL1hwObesdMgJ6/eaZ
AxEScLhOP3LQERKaDcrHLW/iCosCeCYvGdIxaZrOKwiXmiXeN494DU0ra4KKAqSPBwXqCX7D2ufh
WUhhKjCJoWzxMFCrSlFuDE9PBfUc0GZrnS7JUPSUlwEJWdZA4oYYVndJI2ewAggynlG7PkC5QPAb
NfF4uLtudAX6sTTCU18WkLPho/tyyf5RRz2gSPCUvr6cVSXHkIF2/dK+iLR1gZaMH8CfNDhQQlYp
0Ev7fSfLARsM6x0yeYkdd2RAPA6fXxUvaE73yajIrDKNg1oy+huzpPbGHE7RP5OTkgS3E/xrpUCc
NNEJyapc90SZ/bK5ZWxAwvw/AAp3TwC6nKDZOe5W1q71RuPYhibq2KUY9IUtXwU9idfyj+KMLMxr
UpXsX4XboAZa7HXSCFfQ3VghfdydnFIPow4VUQysXFqH10XRdaxy8zEkqBkYUpdbelktRvIbZWNM
D0bh1q3F0cDE3Dsb/jMw6G6O0ylG61KjkjPonu16fZDD2ENtjLiEy8209Ute+PVHsPosBwpWuEcj
/oQ2mrL1g9TOKm6b4wLPijD/42oNdx2uGCNqo5OJT+d2///HGhZJEP+57WQmBJ8szycsR6C8kqHG
FPS0/dRgZoHuDnKmC4zUfHpzfrUDBVSeDFGl67yKO0G20Pd3WOEki5tGh92Qbi+vImpcVWJ9JX1E
u6TfK0wBPrLnNBtxDbhtR7IbEeN4wxS8XVBWzTgGqsTPyzr2m6is37icU0cbsXcEApdhUhBYggU1
dHoqGN6o+Lfh029Kr2nB+0AkGSVwIHmDQuiVipopJ6QLBug1Rv+Sul12d+CbZd/JAFeKIKwi0TPe
G3yOZ6yX4xpBD7TcpYxmrLNVoV5K5Dy3bGsxxv4VAjDui3u/iAEk19Leo8rzqk/gBOk6yHc2oylB
oq8w73+XPyvJuCrRakRgeUobj15a35S9tZ6IDGYHzewbKTGOsVfSYooVkIrgrgduN559UOuxcZkA
pfYghDm925xf5o38WhXMNS+4QyHb8xpkXrBK2hc5PZn9lUx/N/IB0cW8Ex4I0TliEjuoqtTo6cno
uHIG+iDtGw3UvtB44CThwjQ7gx9jzMsuKPN1wckxKld0QLJ6FmFyF1jJaDYfKw4QR5A0lp6+/7GT
NSSdQfY10erhgyc0Ji/XiB2hnCmnpWKr04JzyafHHHmW7/9BvjW0sz9KGBVCESQSHIvhY3xbXe48
nNVhjKfUhJIMO4411MpG1SdduzRoAGqLWN6NHGOkLorLdYAe7pWpvP0DJLYV5kQjF24QuJKMVBid
/ioSMU5F70aJDR5+N6nqvKWX3J1FjpC5083JObmK9nvL2FZB7Yev9qv0A+F7JwDoHPRHqB7sF+ZD
ZYDJa2PD9j3OMsajyPI7SVlgEIIbQFbqzeFbjmLFb1frwxf/e22+LVfRS49WakAxr18Rp/YMXzUT
/LiXgDrj2zv10VixZOuyyRO2fdjcs7Xnovv49/gN5YU1ViD7ZnSt+8Tm7sccTp10Nyn3jBCaOzfV
cRwEl6EsAbE68uJG/bilui9NoJPDBK1YdB870vOa2793ToXRq7X2kKWL6ENkWxjZRETQjomk6uto
zNOvIWvNwuNwf/uLBpoRHqvZW5Xs+31C/e/xnk/M+DZ1l6gDSI/IVhvevDXo7NrchTFmo+6Ca66p
KeuZx+BiHi99EfEnGzrJze/AmhYRLFyVFVaHfuWTCsqoakXKRzs45cMub7DLQI0PInq4UQzMYXfb
gGFDBiSJxbchOxjVk65/pjHidNcEgKg7F54aVhqmDG9czTMCYaTCHgqc/L6UaJduIY30E3VTqYbD
RbKAVdqlWk6xRmpnpqqvY/Ye4SOFu1BAVQTe8RpucyMbmi/O31Sv3O9ixkSDzFBpOoNS93V3DG54
StHAU8mEmtIH8IIELNMw96tnIz5WPHjEubV1R1HrWlOlY/y5n7AOgH77yYksG4HUZFhFiNfxlzVY
IYZyiO/VpK6Euv52EdIe5BxxVs4UmlVeP9XJ9Kz0sdxXbcOhbtJHmr0ZZ8i+/ARMmV9KlcHqHkAB
bEa4R/Cuq1eaphthnF6ugNQq26mh+B8T0mfdv46E3vEUdCV6UdbbMQvQBjY4e4vtYyUjhX+x4r6A
338eqGzK8CdrEl/LIfOZLICyVsNJNnQ8b9HGAHEIrrMiBm3o6AKuhDCghAngUZKquj4N8tlR1bzj
9/6jVDXgqRO0MIPJ6oFSjw5PUIR2gAcHZqMDCQ0W14xqozdLF22zaZRNcsVKWAmsMrQ0S/nWiRBe
ZdE9nAJeKOG42usmchhV8KmcZvHo6L/axGTf/Tv8HmoLcNYlKxA0yzq0KIt4t5gImMHcj32F4q4i
GVFnQThRIGo6gdFGAf8XaJqV+5A3pmxYjyy8TmJkrnR7Bt4fckf775lOKgAAW+8/fCyo81wcA0AC
mZorIJ4CGKEEjD7OuJHtzFbswW1YXGZD4IMfS2eQKZU+OBz3J5R/1N2Cd6Sj2Y5DZAdPcj63ryGX
x4BSpMI0tY/t1eQ0KjPV6kbfhKVJ5wn7m1IdHMxPaNwH4Rt6GmWCRgAT1l3056uGWRzs3czrS9T5
5Twd7Jj2FeoRAKvGUpFeZrwogoGRvcc7PP9KgVtf3lfJKSMxz3etwYFCNl+0sNgqYYfaIAnl81ug
1H+ERlsUuSpy3vBNk6nkiTLADiYrHyAjq4mK6CrNfBtCDm1wsZrBZ3VEo1oJLLQGurhXcPP295FO
VReZeCsGl25WaZ04J+Xmgv0Tsyq4U8MwOfrSVZ9TfD3IlI3aAx74ko4mzsiWz6Hzt0qoPe0BkcIe
aX6noBHFH7Fhm2TkxTkNKrk2VQUIJkH7j/ODLck43RUtYT6XXGt1x2FX+AK5gC24kGMqT7UuKumG
Jaq5waH7pBi+FyABiKda/GsT+DBexlLyQk2R31VrRdH1fnBse9OHH91RA8Rsveh3CKsWp/NRCW6v
HIFyQET3di2T/s0rABvNVgaspXX4YmDeJ/uhIIaJTXKpCY4F684DiFiKgswTUDQMHoNEEI4S1iin
ia9JBPBsaQ9uYPgmlCzwypiWbaMXGSNnzid3xKWR96PRnsCnxaPm6zssPTUCOCRtflu6J9hfAGgP
5VXhBuesKbEkh7GsQwRFkti4UMB6vnRIEXC9yquYpZKMZMszsnjwpqp0rOZMBCJhR1tH3VtUr2yJ
CtFzsLKzK58i4HjzPkTAzxzw//OCvfCgu9JjNYSW7IPBBYzyJMFlwsNZNPBG/KG7ju33SCFqR96a
RUBhd7U0eLqVfX84CDx+znBkok4o8gAO1qNWMFxJ3tLvJaJvadrRECsbfo8PcxdZRJzESPw1X65e
AuwE9HXaLiypzQMQiS/IvmFQADCrOTR5bnjjO6Xt1xyFUxY4hFQHSJYberbp6dSPopByYm6kGyZc
aNIyHwEgwGJDc0/WOZLAqR6ED20TOFRAMZnOrDpBgGrTAv3R6Xdf2FeDW9H3gWCCKskA8bl6cZdY
4uUwoXQXaBiZnPY2dZs5oHoU84q8f9Kc/JfLi5a3bzcMJu3ftZvhsGbKUkc9TFaW785os9IX2tR1
O/HiuJx84nowVZqXrdMaKVojboZsUay56+Bot9m1fb5SW+tIfMdKtPVLL5Ck7ebHTJML+zlP6mJf
Vzs1BpeFqHXz6nRAdEMZU5c+hAcn3M7QzFmtzByR4CjyalEKhGbX6ZdnoxHytpe/9ydjOeGbicMI
DrcUZfkhcGMj3QcgnQcQvega3gtdnor9lX3mJgCA9rWpY5uR4OXazfWOiQrpsTGgmXwFVanRenC+
W1tB+uCk3tPagzRgc6ltfs6TNqLardcL6hj8RIcGCH/XmyKBQzcX5GyoVsYB3c/VSyqbYCBJthfh
pa9B/du8HcqThAaVVgoysbNSXgDPPlkJyjeuC9xniGOdDM2W0qWqktIGTVNMn2qFwpB5K3reCaLD
/e83HbUPycvo1wOB9mWdTecTOm95RwjAfqiVGExx78aSQePSI/03rj+HfUHOPIKOQnwcLCtLMLYT
fgYI94nmeI2NAKHY7PukyEjweOwZ1N/DAiHw5HWwBhtCOFt0L/BWBPSmA7xUCs/rFw8gYhkVkOx/
i5YYaf1qdQtqTN9xy1azekACfy+egUvc1zXLDOnzlEVh8cfae8s54gU7WvTPKJsuiJqrvvJY59Jo
KN3cVstRHIERkusq2e2CeZph94lr5ek8iYF/U0X7S1XOa8BWGMxk5R/Ne2+NG0JA+FZCy00ni1jW
nPKYzaojMIcIDiffDZ/YRDYcYTMb6lWCBGXWB76c1tV30BPqknsBgFX6LXTWxmSebBC/xK/xs+Or
bqF8Ylx4rsbSxTqRM6rS6pHoCyBLt0N0BGToE/FR1LWAmNVysFkDNyunY5kL3Yde6BG5xxRW+OoU
KUv8D0rLd/+x65PU82S2y4KZMPlZdXAzY3Z7l8LronOcboN9rmva+y/4Bq5W8iIL87f8T1YM23Qh
LnFrj/kXO3tULWndr30eiRy1shSY3LHFD9c3mWJMzHpso8Wyy1mEZxkMPBgDTu50ps67H9o1aEaU
xbKgvX10OlNUcQCNyq2O3KWssj05Ss+9oKDXpYyvO+e32vCi5eoB8IPUjLKRBUn55YqpPHziVIcJ
Z31YKdtuV7rxSqla/xMj2bV5WzjWYepilt6Z/ikvgzDc0gZwkBZrexjEHjX5vQ3nkecrEYm7Nypo
QlZ8UAqNAmn3YSTo1VRqK9vzNlC3N22QbAym/76sBv3fN+4Pfo9lHwMUhkguKo29HHfXhNfT7AQ3
Di7+arfW3GtppGap9E3jBs1K6yPCUfkE2l5GhiFeJ8lFa+J9NE7PqUwizkG/jOHBFIz7btQcY0Gi
k2jtAc+mVCAaw600i62wn4GleK1HN2Yr8jYcfSql9LAKpqp3mHASa51bFOD8wM+2hckVwj0H9iQo
lmRPUUMfaKAoL631p/MUYcJpJXFjWKlDFHFqODBKCae5OkWgdnN+42qCUGu14xXdWL6Fv2pZTh0y
G7L/1opiu7gV62z4aAEYFbwcMXuvur/SDS7F/9SmpB54mkkjF+hSZVcJA/EsNs55KxxeN5ZzFFUa
QB8qFDJATqpOm8RLj74GomjaWhj71ngRRzDSf7cyNe5l5yz59lUxNzpSjp+W96e4bXREYZlbqWWd
aBjbMN2PVOmvmDuUF7yxxpDuzNghbKosE2CnoFyPOooWdWnXJxom9xEaMaYT0rnWJzW9XDslBNee
awP6fV7ELnhsUIwke9uSS6YlC1d9hAcnn9J+3r1EKR45FkK+7rshM87gQIsl8eCb/EE8FPJK75GS
GN4UhLSa7a4Ruea4u8MKZVEaDhrPbujaxNleJ7fFGc3SFLsj1ph8mhTXjRrVJHa0xIzAoG113CcI
JtkFQwWbowP1GaY1QaTroHY0DIwUSJ5rmrLmJvudJxqd46m3NNA9RvuRcBoQBKDDxRWM08LD9Gb2
zUbRXa3Uv19ShoIkUY+Dj3uggjZvc5aDVyHiKj7+jvMr1Xk4vPtgXpH35m4fpF9EWQ3sJLgKb6wM
vTF6I0T0FzcDuGGSQhBqGSs4LQOLeXkKEkjagZeGxX7XYTQ/Vs/kvAmeyknUqoh83YRZeF2gAQOu
NgfDP6wLdhDzwMfhXEICEZsTqiGERCORsNotetCMLYaSpIDUd+/F8odWp40hFCQJfmhU2rHWyS6j
pTmEcqn95etUjZHzy3jTI/tqTZolGnov0/pMqGvP9LeQk33uKyqZOmVQBVlg+WfwUOBU6nm0EMvP
xWz86G6d5j0xe7hyT1QXHnhOgoHVhGOw5xFTOe1KSj6fbtqadGbuP7+OcV1Lz5FkUkVnOq791yJ6
SoTEY11VH6dEEDOJtuYcMvp4UagVI4hMSERS+0kgaLug+fRR8IJT+ROiejWTaaeWo/4g9zuBtGMZ
P8KlasEu/0CZOUl0bounlpxEFz6VVmT8H2Dk6lhHxt5quk7NdnxSH2hMZR/BaH98v2Pqex3Xr4M+
FgA0uBasFS57hWvJwFttH6wcjSKOYKIUNktqFmJ2WHnDxTYSa/LNEsEjJKrKuME/mtSHNIMhssAj
QrnM+NjcyWpAyV2LdWQ3OxBJYaKBjj5Iai4rCNCPipe5/N+2nCNdjp8AKCml7RXuWwmqeqEvqw9X
K6yenXV7KwdyWl+dWbRGLZKzomZz+R43SkCNYKyKRfQOrBJy9s3Kls6kpkZWS913jsYIvSLZBOm0
T51SqAe3j1s1Y5lXcvwWIQQNFOvXuxveoczOT8kUzKhONOvCPe5pbKRKkCftBLML1au/4Kr/+e9Q
89YsDe6zwmlQXExXR1V11FFT0N1+sE+J3UNKZPnPu2zqxwikimku8QC+5z528ITzgJomB45nV4qN
R+iL3OYodSgrNcPbUe1Wl1XeY4IbIzKBU70i0YYXlxUNR/UXUdjKlEaphUlozB+iteEgLgXL/Y7A
PUBKlX86pZY4+gXEvzqzqZv1wko9/+NdPe3D4Kti2kow2CrO8qThKp4i5rOiUpvifEe9zNabqcFN
jme5/4ZuaVqKr6fnEUqAo4zs/dh4XH8RlPwZC0cFMCRzWrcNlD+TL7wBwkQYCY6h0Nok03TS31wF
UvVOD+LBsI872cVtVGgRdUbrW2D6rqE9m3SF2pLGTLvUlv7JNiao/XaWvdMPyqX55IW2rW8Xgkwr
Zhy5bzxeQ7UafG8/Vi2Gil1EKRK13EWLb+UjlEFqAcxHU97vOISkWUAXpsuNRClRHx3W70ht1sQb
42V3H9yis4RcpizO9Eet4qAC24xNEnF9jnHHHEKfsBXK19HA/i50NQITxhfX7e/PuXgr1O6hPlfT
KhmZ0z2ZwpRPUDAhZ6gLEoFWXuX3AablhpZK2+uFmlMt5AyOgzt9YCBoGfaDKjzq93CZmIc9syJh
8wkAz6AM1oJ8bZFgacvYB7l4BZSkEy1sa8hdm6wGGeCro2QGNwJJT9COJUlorIv1JF/NKlYxUKdZ
Q9oFXm4zqiAwLSemUwwg6mc7q/ccxC7MDqoicQB4acUfeeydXjBFSD4YQlDzHjqsCa9q/JA+JHJA
pQwjx20gi/94ReZWmbT7YAF8SNDJRFyCie547Gw3FEqELssDX6xd2G7n612w8lA4odSD/kBLAM7Z
K/2u58DY5K5x3yJd6us5dzEPGCtT+T/4kIuKgLE5e0J4nC/H1fmrQCWrHvSfH0CX8VpD1o0e4Z49
Qz2P9UbuP+v1vPojhxnSMIdO+oc+h37PDgL4ez6ZZzJEcGE3bvwayPYNIUAfyQoZ5wUxVlPwWlhQ
XctVfPL5S9rPDv9f9mp+BbeMXz+LUuJZUMBzCDSbgY+u0av9EfjKFXU43G+PTXMVWr4tqcE8Mwvn
awxkWpUQPINbzVR5XDVILynISuMTgr1qZET04Z13uK7zIlde5nN9r0JEJ4kCUSDELugowYQ5LBYU
1eiyJdnyPPIvKoGG9hdMlDFl9GveWHZWasj/SwDeBOyggJkPHbPDaLAlR/n+n6rboEDkF3bvmKzT
KKZSnuhGGjoWQcAuaPqKahEvM8dzs1+Kfs+TX2bzBj5/b/Aq84ODfBQK667P/ejuWjK2bmq57mUP
3jj+F9PRIxYCh29z9jlCMO7xn/UPKiKb7ol3crfRunJo3Aa57WKRBDWAIo+tC3Om2I0huMHExqns
bqxEgRFH657JUo4DGvdTTxn8kHTeVizssUl6Semnj/0FJ9diXWlLlYgXINnogxW1fgCnm7/9kctv
Q2S9k2q/kEV6878ko3feG8KVEN172CSaT3/vDGQiKs3tKIuLmgfmTQLnoh2AE9ajpckVHZRSJXia
b6QTCa9GHygS6ElNAkmaY8pIOnpwkRwT9hwQLc1Xahfztia2eUlDFwyM1QTF0YMRO0+7KJnOskr9
q/uTYV7gT1+xoJoV6S6Rl/OJHPBTv2GTRlmcAPnPmcImUP1Z2/KeWkhBxnfEHaGQCd5PWTM0jxCY
lMdlxVn/FLzKOLUXc5iY42WGpVQqiqAfdyNZJhaky4ZnBK3pe+aWdwp9oOE7VNjqdguHRDL3n8BT
gzX5zbCZOxOKjzD7ZhZVNL6+MmkbAYGGslMsY22N2JteV+bSqiCA053AkSRxj41KJcvvkjUBn9lX
2YuO8Ie4nI+VAoT4qVpo+fwVmoH6Zd9UtE0d4mVfU4MDs7tpFFE/rq9gU1QOS/5Jrrl6Y/cINzXu
6bhXMUvnTqV1gDG4E+Sa1f+RzZhFMon97mGpL3tsss0fsiwSB0QFve5piO6KdVOfX1herDSLE00U
1Ld+cdQvfW1JPz2oT7SZ5tfsHoe7pT35UE3f9bl7iJPikg8iyDfdd/d6l2uifiPl3agzSwvQoaae
cxT9VjbFGBQ41anvT1QDXwhJCpIMmxrLQil68zoMioZFywsfnnE5cxLNNxHJ7UudY3IseDYZ5QDF
Y3huaOEg/nvvb5JkZoOpSzqxZOFsuxrM5EjocrgEp6Vhgtw1lPjd9Cs31+eUtIy7dfZtTSB8xobJ
ptE3N4FaekP17tq6AKNpsWJqiJfX8Ft7A2i5b60EHPuWMhde0HgWnIOAZq6o79RVfLikgdAvoTpq
0x8R5/ZZK31t0KCdce4ZfN6ecCFO5698MzfCfAqGca0n+vElYg+OBpg6PO3UgVdusRkI3xpLbLVS
MUYM7ml55T9wUmdsgHXEasZicA9TDcFaIbWI7DVDsj0u9SiGdhYmHXv/yTQzaWUyT5kMMz4bc9KY
yw3BucGc+0bfbCRU90vQFwJxbTaMyd7PR4PX+EXZFnV2hVjJUw1KAPVqFHH/EVDnFu7M1zMlJ+Ap
ge8DvBjL74gDczp++JzcpzmPTRyy2hqR7nrZkRSTS8+IfhL18wcvEEp67WKD04fyuyoFvEaKgCKd
Pe38KSg1kOrg/2DmHo9K5MLYB8HFwzMzL2zyErn9aCrSOTTb9YVrf4V70i+UkfRbgJkJ4XhSdhve
VX0ywGIghEIGdtjcyFt08R/LUHQSosoyzYpj3uToDpxagRA5UrAiZ5nI7ugSyqLZqbt8OxLgrNvP
QOClsygN3ZSeSKIeB+YngOlbHmb6hmoBLtH6HAVccdDiJAMfrM6gCdT4nwkJyeKedfC1frRqD0AJ
Cpzb66oNbSabUeyGbfnsPsKKXqwJlF3ATTNKYRyXa/IGnR7fY2Ah0HGQQdzjW9ltXGB8OJJxjs1R
aHFB1E7wNZX9yICbK5YvVCvq0w34WSAxxlEfvr3P4cxLuZN+dCJG6XSo0LjUhepO+TU/HtL9tfyG
6pmEFbdizUK7I0vp7v7De6HcOc9cEVYcSJATYmiYac89UxfmjuPbCHrX2lPtAFhFAK64YJAI8HDg
tJM4c2IJr7oZC4fKDiMXkcJ7lijVGpPbOJUMyjo4uHICUBUsnCqp2V288YLL3+aJRtE1VONj+lIy
818FgVesSRIiytr+UQVDfL7KOpZkuKpmyL5ueU7R9xRjnwPXJkGa7gp3fDX1vru4nqTmA0p0K46h
aUjgsX6XxitvMpceCwHtL8rxWAKeHVaOLYS9x5n+wCJRBbQHosWv2omLcolbnf/VL6wmgcPruIdI
L46aXZ1UtNmTQ6qxcoo440nAYJEv6tAxQaz89a2fAZNACZUrHhLNLLKh3NFQrOrwUKaYxFeIGxQV
b2sF/562TFbCPc8YrFdlrWV0tYBWLQtCp8eyWKZ0N8anmXz28Ms+jKxQVPjFRQm+Pd9wM/qNB3ET
dLvhqctvECmsnMfX3m0ikrupPPhKDp/+8zxsuPEjWrygj6HwXUkpAip4nqm2PQjk+99EhwO5WGWb
9VLghv17aXXa7FLVWQrAP3iVDbQdcenGbkBCx870gVvlG9RQZT06pp2TmCgSOgb7CNRnvx8RXgc9
Fb5svbwhbCGBv9ZrdweBgEAbb2uccvLjlS0/3Rnk4cE+ZYASWr93AVd68VVofvn4krIny6NKU1oI
t3GQk1vbtfFnotq50/iTfAztQIe15I/M/ztQFksibdzWaYsesKPjpTf0G5mRfVnOzg0mPBoP4tKn
0OVz6vREvJ8UZTFesYHfmRc0zbXDEN+m8iSlWwuHMA8QSd2kpdHgSwYydUwoNzmZt70isr7W1c8q
oKTtNhfylPe3HyPuFfM7oEU9gVZniazqSVD6hRnugbFDdI7Tw55FUdkGH5kSruhwOVfi+j1H8onW
azPMLqc/r633VGYa8+ZR/xDeHjWuckMLlmSbHR3r5xxXae8ll65ey5Wyt4+PAJX9lihdaxmyk64P
PzqSwNKMNjU7MLr+Se1wt3oCLT+/C/St//1ba5iE9zDvVTLbtxX0d4jH/+iiWzyLnSP4yyG4JIhV
ItOApLrjhein1PVMQ1Ww4bTqgVc3tYhXe9BCUw5SoA75FolabFNN7DCmtg/VB+Jk0iL2sQfCRTu8
BjOGWub2o7Fpga2aAaojpJBGOqgW0doUu3fVado4FHmToXCHF1/AZJ+EShtOnpyoyXGEgc5Kk/xt
TDyT5XyzEuzB4FG3ZorI9Lb4wv5N3DCaXYNpLsW4L2DKWXDlorBU0qRYZ4fw3PtzvGsD6sqXU4m4
EenT4RlX55WT78rdvuJXm6OFQBul/mMaDBCEDnwcpSVjtdOEXQdy3F/TdyMX5OP9Q85/SR/dHPOX
X2WvkVL0d1okam3Of6iQwavlITuta3RiB40y1cMkW0uVwZhnqPWbwXw4+sSDPrj2MLZxpiKvnx1g
uiz6/3R3H1JTq6wXhLa+fzGicoTHcedD008GS/FpCEJYz+ZLPgi2uctcqmP6SI+QitGV8ZJ0wVs9
BvVuAV3kDNz2sUl4zVySX0iHOtLdKm+drMq8GKDpo+IXetWdO9lBAorkTfQe0ZLfgGSlFtI8SVkK
5qoqrA07Geiv5kq1uVhL9jfYVu08fNhTmqTdaiCgsG2r7cFDGtcdLo0wa7o3lHc0YONIjDblE6cv
rPULgKZRpPjwsmb5V5t7mBn+mcMM/JFE9k7wpgUBbpCVc18YArb1LXY4BrNFSnqVTcBdFQ+9SzQU
LbYKlDWIaCeL6XR4rnRDCKYu6QNm3Fh9xTr8AwV77AxOG1UCD8mzAogVfk2tOF3Y85NtH+lm1PAo
R7519LvgL6rSa5J5wr17dHISPHW6pvjmGy0AeO2a4VrK0Tfydbfqmm4gAm/g/yz2ZumhV9yZ0Lfy
1ulSkZ/U4eiQOKEeO+rxZYzw0kJYRVW+2DSvuIyLCqwScAwjye4nPRK3ybS8yHZu3Pz9namlcALh
+csT8xQZxP1rOXRjHCLsY4J9+vJcqx472eB3P0ZScEBDrG7kDYSPMYIMHj0gOZRbHumzOoGDMCTT
P/tHTDibfBSHrD2+8pvA84iinBfkP06Kqx3tFl0k4YatxP4yvFNZ2DjPgwMxJ8DhQ6csv1UgQ7H6
rie2TtkmvxgyiR6LJAyFnlRavIl9wMEA/9aKmobZTk+pgDwlZ7jbH623WoZrLuwhqwuBarjQxytn
lXXAV6prE0X25mDmXC8u22U9m8E8fhVVTJvZlSRF8xOdP/wAdEIhrk0r//E3PdYaAURjxhJikCea
uumhdex0Il8qeTeK5DgUG1y6nKA0MU3mL/eVfprkBtImunWeSwDdh7XW8CGoiuADsG25k+3VNpUK
S1uECIbqDuiREVox6CPGjy6eUwbbwuzsxmjBZCFGQAwOYBUtoyW8kq3nxsiG9KYdFnZMRat4I3yR
XIKh1YlMKe1aPimtszD6vGTMO8HJBcm/Gl+NUhYO4mDnh7HRlM8s+UYSByE5hOlej/+tmH7Imh6X
GssjNBCwhVIBC8NJc3z5ut8SNQ50BlLp73Z15n+RqbvDnU/3mmMjYeBBbdScwXf01Luh1JOOygfB
ws2TBNXlAokfwmiVOnAbPldyHOOBMxQFNWPgMdKHtr40a+YjSzukffmAWn0CnMg7zfT8SuqL+ZnZ
TvuZI/NTHE9UXQSYW9NuiIjHbyRc70Z7TsZluFFca4cHdcFdc9anPyi46tI2uZW2WEvCaFWr2aGq
4L5Oo5M65KyPTWjZsNyBtvntmiLdYZ5W0N1pWoHgQvl5/Ca5wrlitzyDYtyNsmCb9S5xKlrmxJEx
ATdteZM/pYMTq2LP9Q9QvRofgsouChHff5WUzIOLaqNhjSqyxbCuivqstOQ9GLMCS7QwKAko7i+Y
qzTBxnqaPRUaa6w8Nv5gHNRL5s6eoDvCwvnM03A4BRf+tIHefGzm8B++4V35J//eDgQqJZNqjg25
gebEDj5lgEdTfDu/E6iVyzg3tCuWGt0cfiQMtlQE2RciPZzsOgwZFmtzYqyC7hQZ2Kt25I4F0lX6
w6Aiz4nAqPGbVvZzajUArP0IdNyawOO9wqTXvNZaLVmS5H8oflzH7ZWNDekXNYhExDKvrSPAtOKE
mAzKg0ux20+4a3vWq3yJdl1euNW7eBZwtyNp0hR8M+HDX/QoYpE0iQM3gikkrhT5q+aBelpw/Unx
Ihbb8vVnFpRr+/xt9+Vdi8aBxQuX97GDJOu6+DDnYlgUqsFc/psS3tjMLWN8foBDoi61mCGy+tEq
dZHE1u0zaaM1FoRZgTV9HXCNm2jFQTwstCVmvVQZoExEckprLRLvA5ncbhw2KwQrPEMKE0Rwe/oY
GOBok2LScZqhQWqFWh+i3h1MWCZg+jM0r+wWVXmexG0bSMo5j67PEPf1IPkb3T7IDF+tqZhc51T5
jAWUnC95cTvrB3+AdmFaeXwVVO+LAZhIdItf3e8oa/DpdZK+rD5oh8tsu1hnEZRIAeGUK8yCGzj9
4jChXxT7Cm+4QSJDhkgUYnuPO0hOct1PrCnrpbmTBGQLSBOW71z/jAA5HcSIPvqwxqIdgg6aCW8C
IadLnH4hDetwNRp6k2NodrmBnelgXM6SK+cW7XWysU44fWRDpKvj1q44a5R3+JuoZg1/vMVky9rg
r+nWuP/A7wSrNI8z47V9MP588+nBGghE8CVdgpEN1HC9iIi2GJXhwvNUx63pmQh18Tf1QHRm2sCg
rCLhDGaCaD09M2jjJa1pfRqnG50z2Cz7Dylae/XaerXIvrtP+IcXOCWboEbMQY9Aps0dzmdbf3YZ
NGRtz9T/IgfY+s/hVPL+i9XOcPHqbYq14xtN8s7WAxxRrr9vbMI7gwcXIpkYE8YTF3yacMqdycuz
V0A0BcjERjX0gwwVyCyA9icKXhp1UiBIKQthhBp0IfkjcpMZpoE5QmEvVXpgBZgXi9IBbUsiwRx3
KS8sqBXwxEOn4rAXwsIrOmKkOXUsUsjaKnfKMAZSAlUOLqd4RLKKjAdN/EhlsPX5JKvqlVDGIRta
m9Fw3N/j4/ykSyN0axc1JG1oPsyv4PW2SXQAu87Y3aw5gr3vD4sS7iSIqHBiKRsEmhX2RSAcAVXN
v+j6sYOdteWFq5id7pWRykbqcA+GiMtY15kdn662YVudGRUkofdSy1N9/m/cml/Ecd8B35LuNGXg
kY15U453mmwvSLlAh8BZ01lyFEhw1iPKjWP69pcMyC12Dd/c+kzT6FgOjEsP3/QIIOT5NHq7085v
jTfZ8waczwddxowMk+gdlFaWHtw7rkiUKmQgg05nF5PLQfBrqEJ7ovNoRfJlw0hYPTl77uvM/bAz
cw2484/T+AasioUMqAcQMGcRKJV/h1FD1elmvo9hVS0tHSWLdjF2tGx4rzdsxajZyQ2URZMNpYiU
nJ/w6AB0zuehAOOYo4+KIN2fmClwDhWScP0+xXgAVX4tdeyuYIQZX8NdQGAP0GBPAiTGilZ8ZaN9
wlmoTR8wfM4wfVuegxOqFxrLfIEEImA58A8LiI0v4Y3PGUcNvxbahfJoZC0a1fiY0ICrZz+CBY1U
hHm54TkznnIwmggTZQQYhLJQOCaXwagDdAmzZXzH+6m4I42wIqKxPcAl2z4E1e4L9i/NKglHJJz4
dDV6304DINV06H/vGFT+x2ZYIz4UUW6Q2R8h1sX7RmAP7mrLpcfsX9gxMviW5ldhWN4jgxCXXDMN
2aO0cU8/vVRTucESpmY6hg30NPbv0I5Ui3Lk2Aet7NVZYQ+xbR+QGYYkDodktxwTXqaNbANrc6Bp
U98Le6FGmUIr+FMXhpINadaOe4eeJZUJBSwiTxqCisave9dLkr4VjJq220FrLVGsoZ4qVkEMDPEV
9h8BcMM+mbJs/DJZl5VPfH+nXJvoddDmBk5m6nG3IKnEo3qePt1rVMCUqCJ2IJ0IlvvAnhO3RgHd
h2RKwGbz1p3zdsRL9N8Sbz4BqNvld9/lDqIlfby3L4uVEJXOsyYSvZ7L1ulwuAsSWYut3gQyuqSF
wnuVXDYXCu5KFhXvzjynYmfnywUZNrcAEVq++eGyt/QYdwpHdAr+cZFuidKdYmh0AEv+LpyZjTD7
HX/KaeCaPRdXoPdsnX8CIGXOG4/JHbJ/8NnEZifFWk7yYsbgbSkbeuocn3TTaHSe41J2mu2qtmu3
wkDp+TwF2yQa6PeLDTnTLDHHcWJi0/YJg8sNsfxZRxcdLPWDqZCVPOTZmQU83CVKPGyDKJw1igfR
4S9qs8fldL7M2Z1ydARWKFtVKwZH5dh1v12srIdOxHGe08/SjNUBNlRCveTUPbydgjolHfpms5GT
kr7iSy82y1SeE7CDyuGykemJ9T1DK4PgNTiDC3LcuSVvbpZe0Cctn2SbLVPc3YaL0Bq/vYfSrlmw
RDFSp81iv9tWMAR9JPO6ZpDyMoS6CcPyCQ/VG9IkYTx+cg+HqboD3ZE9r/OvHIQNWyLR4zQ9xShW
9rbtQL66TWohKfC95SJqsv4EbIfJHKK61ISa/pFGkjB2C4z0h+plIGNZB1i7R3rSM+/VwiiVcoTc
Wcrr0+da2atqKKQEj3RcRurBoTxePLE8wefmziyNeu79Fd+LDfe8TVDRw5cAg7b9emh9ER7BJCbz
utLOmomv6W0cE5yGUn678AbJerWrpJdxxtuxPiLt8Gd8LVN/fA3o+KbY94YV/xOtEn1n2MHCnNN8
2LgTt7YlPHOmePSS0AqJDEEhNbd5Lo3OuPSct0+2DVRg3rLpCRDko1rsk/d9PgL3V/GzdHmT8doX
h3/vWGY++SnqAwh3VJGZTeBvR1tcDZitPg5u/3f985FiZmbhBSQl+DXvdYZ/kLZpF31IGjIOuvnO
fNJYuZWl2cdJJhByKJDZU1/XWkb+U88qq6s+KjroG48r4IwD9mjG++5hh9mVoUPPtyCzDV/cXRFQ
WPZRn0EsHmSrH6TL8nXBAyyKnSpCQtR5g2nDCWl6kCnwlnh+rdz4wwAeKXsIs/aC8EXI7wWrw8TQ
WKgVNVdlWe87zxsEAYpo3/BfTOes1tkkZ7MyBk3dyRmdu6Hjxs/J3Frp48BWaDdL2F7spgGbZpNl
rdb4P1IeMPmviZDw6Gvspz6ojhUlMfn/tAvtW/wJmETeoTi7X3gqaGScnuOXABOO2NqouIysENYj
q1VczWjOpcJ6c+9lXWmBDDGvxBK8Jt89B7P/s8l8qWHbLv2OkBKQfoENlxAi70XZwCAzQRYL/k6y
Dr1fMZN6QSu5pSuMKI3M0ENSDOmGe3+mqHhwJ5qv9E+TKhZgffYP1HVW240nuO6W5GOtIa93/otA
Hz7mTNHYD6MGX/40pLTaa2C4kohy1Acz6RsfQLSrCJuPrB63UnLX5OiilYp/AUhk0HDpOiQ1qff4
Sg4QAdfNkjcRzaWX88XUXvFhSjer0Y59Ntr/j8N642Do6DIAE0NI87VxlBSXbRFt4KnmtGXy2DHf
9VG4oVNYSG4cs/scMnBU2ySpoIuEPRFfif3Ikk9vDWuBvJU/zPSSziZZOampfga7hAGCmattKVH3
U+LmdIfGBt66UjrFT3PuKCBL8gAZeXuJG/IRrLsQ1M+2sE1hU8xEycc6emq1jE0bPXq7uG0A3cMe
k8OOFLHO0Y8kinA5RuE/gqQZk+WqVJdy+dDY40vsso35rI8fPYpPi0LnxFOUJaQnHOe95uie/k4l
dTzEcSTOqGdxFbbg3HZXo6iTRxID+KV5sgVxn5Q3vQbG4gISroRa8dugKq7Uir/BU8F40C7CDvhQ
bzYI4myxFADARVVvwY/n4KTZvrDZA/RV8bRQA8Pk48INK/Onikl6Rm9OMxY7gzBFQiro4GYS/HfB
FHNa0am/++1nZDN9bSR0ylwlXfa5pwbnGzUN0pfdIgj2cq+56PmI47XDl6KsqFvJGs7HxXL9MpFi
bEYaQZuP8I0NTGbcH3HB23oLW703x7Xz23ZqrklIHL18QQcUlTzNuiOjNMK6RlZ21GilcAfaCnfi
akcM9gI4KEoHBIidjPeIsC5D/iRyoN1qKnGQkEVSrwDfQGPbBvzpGcflsTWK+hrP1nRehGbem80a
+NC6tovSHWm2gia0x7pNtTG1W5Kb/E90P4bXNBliCQod/LTlM5KiKH1502oVs0+k4w+o3L0I6KWH
sV7+d6cSFr3srPBRNmEEHDENxSgWMthI4gMkGoMmMk9SU0nZsR4qjORTPnqVO1fsaGJKla4LaVXr
ku+Ex+1YkwgBEZmOWqdusD2HfLyPqPg52FxhevjU7e1kqvbONkltJ0LbqRmma1UFeE4NmQz1ozuJ
Tc0rBDNB3JNqisWdYWTI647vWl5hWBbrytxWuqctI08VtjKuyWw2x1HUVmO8pslx9QSTCE64blUT
hI6meUxASGZcVgNcR2Ihhx3w07sdJWC4b/8vCPNbwlV1RiP5lVSPuzCDtWsRBU8i95dIBK5OrtUN
knceQ14a6S68O43rCSmyUQ/46Jc+PM4lEsyttkKNPzhueWXLXuezwM28xzVlYFJ3Awz2UcnkB/rf
EmxavGtQYtF9vBmI+aDPEKEK4XpybMYjrcqD3rA1mmwyAtR/WkOkgfp/1g8VmBiyYQVUAPEuwoM+
bi+GvydKgnNDllIKeeCaIDv8CRhEmB//XUcQHL8ls9XsrT+8T8P53HfnmFO4wJFsbPPsjxv3PIYf
CfQ/AjAnjyEC4knoWxk9Gjv7d25mPYnSPQYRc3kjIYDUIpG0oORV7A+Wfu/S74MbRS6TTmM9DmbM
OnJibycMv6+x1PXMIj0EX7oGHpWroL5sN8gcEINtog6ElSjZvCje7SQXBAaG+hDmD2wKaKtV0a2I
+8pCmP6vTs+7Oo0z5IbsnVrsAO2cnaoDGf97S6UfMCl+XjhHcXfRKq9bQ1tFzjrVUfjKcitu7DZH
FmVzWFHpjRKCAl6uV0vN1wKq1mmGdkSi/VtSqwUz0V+3M9Ae3veUHZAk/9OkSoHvYnzoMX6c1cJK
kseIaz8FhC1pGmhEJNCjIxmiVs0ljtJ9KRbe/3aFWr2KwXEpduwS3Uk0/nTy96Lc5NSubT6waE6i
53Pb1TnZEL0ScmMmJpXFPgd6TJRmlZ7Bo6S2UQJM66zwW/Ce8J2kHapni451wCSluiK/IfvEdyte
cx0zENbH8jhKFKrZIuVAjVWvYcBdoBwH3g7MQA+f89OSsuRi9Dgas5jGSsxVbfHytEcxWcF71HR3
eoK2Pyv75gT178l4p6dZbhyTJi6Ng3v99v/1D4CurmGv/T/Q8NgyBf8BN3CtIfCcCEWKvILog8DR
aig+tZpxX2rZMTmQPC+HCJMBjLsz4bdQWhyn8702BJrMQCDnpaBu8f8KOfikjP6JrKt2RogILpzx
4Tbqj6zxYLOxtuyjdJEPQ7IbjQ/5Hotmhr4kfJaTE6L/KJ1p6GVxF6oVIyEwu/6zeOhnB5whFz7h
fFW3Tl7gM+LnsWWk9skiznQL8R5W3RGuNYL1bTHQa8eA085pLTNbPdXfXMtF03V5afy1NSP2qQqz
FM8DF8pqnvXHyNXBk2Hn3Sjk0qMm5QNK7jMp+5X9zYKWuaDypF/KtJzIttTRQAdNp5lkF00LiyIw
DY0Hv55ux8AJ6cRgUGW1VrNI3ytuXRYTWpofYrj6U15Nl3kPBVIo9IX2TV+wped3ox9/nIgoB4Ar
bsXYuaI6m1Ya0Jk08sBng+2/Du1/cRpwr1Jiym5J2GpMI5oKo0QYzl2BxuUuEjBWi7j57/N4J67w
4J/HhpbBkBzvBV9thqsnKlNhuJwCoHT28E0q/hkQKVEe68EkVvg0AVnNVJAmvzwepZdAKo4hB2nU
TyhNNHIRX4bgwi2y+1piKWae6BGPUO63blzrzUSa3xaIKManVWt5xODKIH0g3zYZqnlZXkmkfPSw
nOxMoXxcW4dad91iPixkdfC79i6j9cX8EgiVEzoR/HaHw/6LEV2e+Sl5fpbbZ9ieJUsJ4STpL2wL
SDMtZ2HCQHuQTM+vEMzbkTdh1Bc1gtnZbsbdeAPOE/ouKBf9eDZEdBtlVe6esVSzoRK8AJPlB4/n
ZVN12qM45QdE8HRNIWJ18icGih6sycR61U5DHhY20xCoa3l3Zjd4MuvV6JydvRPzdXQJkMh4MYUb
Tfp5eQEZ+0CfutMadFXpwuRCZpk0JWhUjTw2xe9wz1ygSbezUfUaN/WpeBWhfJk9n0RdQXbXm1dW
uiHrytkwMt0tPepBGkrn1nzygvEEh/KCLCjea/K7qcboJtcIa5hkc5SWFqIZaOMCoypMuUrvH5lT
xpmwu/K3FJuu6hPqchTd1pSVX8Sxn3gbYF4jLqJYBZtSVGlZJx4bfA4OFmGq9H1P6WeebOAtK3It
V6cUfRrEZMgy4mW4eJ7OoWHucm4pofE8sXZqJeLeihU9ITX6xYqQC2aUR6sKHeTzv5tKiW/Nk2Ql
tu3eU8Z8ZqQ74sUIH6lzqYk/TcqJOVOtPPSxCMaz2TDmSUS3CbUuDeSo7ufrz8ucZ4c7G8PpaBAk
DCNW49euysphmgsBdrpsR4LfwcihwRZVZmHoiingxJxvPCNa8Q2RcCERr22/3iOpp4G8TPbu+zeP
oCvBYjrx3QRpwoKAbsKt4xG7fL86RbxaVe50FBpTCT/4MBrkpnUVW9HibKzmtSIkI5g4NL+crX7Q
uHfYcqDsP9uJLioTt1B+p40Cj8KZ8mgjlXGeQxyOfDRYAsnk9rsAXvk3s1U0P7lRdz7rq79Zg/c1
JTeFCAnc7EYF4IMzs3GK8jGq7J20DucZrmnQdm0bvNwgfsLhnY74C1TL7ml4/olL9WfQDmPXp1IF
5+shZrhUet03dWG2nry+M9YgozGC6+FyJs6JAeDTgZnx5LmaKTs5vltY6qBMmFQaUpGhp8e+bIVk
MYJocUQfpKDebybX+eKKQWc8nbXaPBPMp1fAgG4tRV2X+SgpLQkFHVyeiVvx7+WBQlGP2ZZ7N9Qg
jgvrzFH/zSTECSVPeelfzXnoFECYbLojoZw5AKUsGKid7Frd7qqHc+DFlCqvp+hYiyHsGd/5U4GQ
xSrz67AOs9GfpKy7RLqbwlzsPWOvDOFYKbdx9OZlbOaHdQ3F6PM/UGezh6QTEncTiaJFYupNSgmD
9ZQJMRsdmo4JgqNOaC+GCIZnihlhP7kPnNpGaG6ti/w/7n5bqlthaPYryYJvJ+f4Wtf4br0cFUCh
nceVgJNO86SsEmHL2K8V/g2DbtPDLIaGwn2+MzVgESrW02gYqc2wyhHPmqztciZfMOmP5yOrvTPg
/1yjc6BFzc8pnpmb36qp7XVN8y3vb9Wu+RhNC07sYJ1eaQSAyB2uSFtVRQUZD1wRfJHf44mIhnY3
bUsECELyGNuBqMeRpYZNJkySY479AWrqIZj20Ad/SuuOWWaI/ixJ/KweS9synlAMUvpVxvyNog1X
WzX3oMcd2555qBqx5u1NwLtWxnFMJdeU/y5E2pfcp0LHboq7DmmkQDO4gcLvbNT5kS5ZtzZjFZhK
iKMZfX5LEy7ZbDR7zvEAiiAW9+2CxH4QHiFIFXOluuz5eZ7tA4ff7wjnhp4DIUQuP5Y6JK1yZHh+
vZhUd1Rn35h7nTTsOdhIBfItvgW4QF1xKA+huxyl3cJ6RlU3/JSa3iUsDu4sBV5L7Asfhq1x3qGL
cvriXSjRk4kNN8jKVVhmRByjN7zd6WGwrKfT1WXOnGMv3bGgXpok6j4lb/Ul+UOigkPEca7F9SON
EsoUmjGxoB20tKpgZ2sNeWAasBpauivZ292SER7IIcn9FoxORELRovpHsNkD9MH9gG4agTLDNywO
undiOQHFbjt/23tIJstH+Ld6xbzQ/NS++mi8bHKweJ+s434sfc/7Gf/ieWlFvTzTmzArv82R+JNB
cUe1g2nv4Tb64w3I+M/89oy5+d/d6PM7FNKG7EIrSOILtq2HaEWos/eCYpk98tsgcMq2aCn8AJva
BklgJvxUpxCxaiV/tZ8OIi5USmfDXz89OHhj/YiVGsfBFtRexqu8eUMr2WouxwMnQBCSSX4nb2/m
e6QCGXAKd90UYd0iJuQY+6fWK88ds+OJQgBrnyW1L1Nsxl+1rBkqC5sloFWLs7x8F8dNie+goQ6p
kBxLG2ABhF1gLdPUmjzsYyD9yrC0+B/Z+WVko61A5Yshz+o/qPHqZJSr+YvwMXaizGzOdtUX0i+J
WtiDzw//hR2doazk+u7+PeLLrfZTvNNDTXM6/BdweKYgUT/wIh5rqGGgu+JoXpXscgIf2CHxwzx1
cyRCHUQ7A9qUfgVgjmuSkzZy2x91DdYBXyAxY3GhSbDqiIyXfvFePmj1xBL5DvogeEP16sOIE5wW
xqhM1TziCWjCbbQVM1XgI82ASYlUI453z0p98ks8mLnGbsfYLlRUMvey3/vrRqUuqnDENX7Jr89c
z5u7mRp5+izNq/LL8rtG40Z3BmeOviA7jAW2SV4JzJYbnS6tnluz4aO3C1fRqRzBbORBbFUnBzMw
dWTOu8sjY/ZGR8CZ+pOYPGl/lNs4U9fDqxBIPORe9jJHklLp7qLvQfeYgk3GMBYs1684xL/b/9I7
K813T7vA9dtp9nEerT7LZpSzBwECThxA65+OAaINOi1ElGU54EFI2i/VouwhqwnZCNuBF+8f1W6A
wwRT+pqalfZ2AD0nUlhEJ/Cwq+b5nXt8DnOCkjTsNhUhZf2oUrU7eAEfwtaiKyTQ21KDiOh+bMsK
qv3kDkOz+Z0bSxQfa0N50NbLRoFlXkDbQLagt1g+pp7Oise5PVLWtfvuVUloTgRb6EKBcT+poa7h
vnITwZ72UYcHuBpo3TBRCiIgRBIC3FsdzY0TTDQFxdv2NO3AFUjSVJQGOIqyso1Axkhgflg3Q7hW
vhr0NHZ8A6NjF/+zDIFbK+21O18r+9cOxaLOAJS68PCsQQryvsDeieoFywxPLCXbEH+PWblJY/KW
/l5pU/OZmqhycj3iYNnqNymnWwj20plgCu7L5rHffIAyXqatYBykjFzfoBgj1J1ry2Ela8TS8iKl
LHVcmN//a2TOpHMORXVhIc1BlE+mRDKZQo7fQjy4V2nQStMgM9udGa67m0q8L5vMick4Mtad7JTw
6Kl3DQt30xuu1SfwZyDSFh0+dbjtYanBMM6hldMab85mFt8IzSEeXan9gN79o/0PaHI03M9Mqtvc
dm+M+vS2e45vlIcBfMYtfmck80Z7dZBldR3wMszrZpOe8ONAYihHCDT6HQmyNZiSDVBzfRhnUNZZ
vmyWjObZxabV0xUJzzaDUhi2kO4uSTAntzBTanvejyWNPP9TVnwWmwr24rrIOe1RO6bGhRsub68H
tQEl2vkclw0wq4MocQ55+gcWXK9fQ4nWHKJ6Qcwdi9UEfvt1WKVuPnOc+2wvCMP/3bDluPlobfEH
3rKT/9ZFRpjp2itg9c3/4t2Rf/9rI8je10mLe7o3n/7OlA2+DTQXZHwKMMnpKRpb9VQABXp5T7S+
Kj6ondxAx/8rP+d1tHICjewONZtnS/FAMoPyiH0KkYzxLJp/yYgOctLNOhVYvZJCgt6VO3guukHo
aBEGDUsN7BzB4GFiL2elTqGzDg27mpROkrwM/Evb4coycgae+O1cRI7GrJMlX2Y+NJ5TG8GqCI75
zuEqfrbGd7E4rnON0WzGBNRHMd/U7vhKAmS1mBn6K3r2UMnkv/1zor4eWXYYCSfKajXJcyK6URk5
fKfzkHArM+PB/c6AtPWJ7syGHmWez06kHdcW/fOwMKa7IgdFuJPJ7DuIILkh6CVFwngXWVsBSikD
1YXrtFqlqtak5oFvvIA8iTrxsDXOCIrrqTZSGkkYHqcVzgClU1f3i073YmRIAiH/iD8CocL1lFGb
7i8RTX5vAq1WzfKJb802kYIYEf0fTnSdWqI3eovgFZeKfxsWvnrxvna+TcMZt9GCFU+lZQK02YsN
bv0JY1mw0SZ/IIqXzM3YXovqQUBgeauhUVhjh2Z00UtVADPjXJIIubNUQAClK0E0q1yPQRlNh8Ov
kL4cZiWJpNkU8a23ujW/gr3cqTMjKcGDYj1/2qa9AyMS1o7kdKOsmvrFwpXesy+lojrLEwHPbeve
hiXTlnDxYPDOxLg/Kg1Wl5fXzQeaShlr09XvW15XHES5NZhlt/LKX05dDoeI3o4yaYkvaG35xHi0
nNRmwx5eh8Obsa/hASbAF1ID7eXnoX7ShKuEf3E1El7Otmp/0NyPaiML++3h7NWB/Y3jXcUXezhb
woKDHEqRlYkKAYKTe/YbpLOcgMGWLX+n1tUH8XYTlpNPSpHI53apQkTFXqIPTSF3Dndk0Tvk4BFB
f4Wzz9suHtXuMABtVX7VpwUXqPb+h/qrxjwzxaHmrt4wjCQgqYcLKQ9EFc7MUcrM4nMa9R+5qNZv
SYuaTnGO3zie1rvvMoIOibWta726WbhVO7t6AwckPdpnc1v0ldOpM/uD7UzFaSPYizJkX5mOmnNd
T4t/OjhnNI6d5OWDXwwgkh0ufTuRrDUhiOnBFyGxjR2jOLeS0O50EmceXRUlUwpNkpOw0zPh3le5
mQeecgVHEBscfkwU/uSspIEGDOojnYfzbYnr2snSSXqlp5jOvHK+3JHwYmdx0Y7xfI1eqcdgG9wS
3AFN4PeNaSrw/0M4WMltrxHJzhYN26daHmDKvZTchCuf/4iQzufOHmckwwynUtZwZ92ahNHYMZm/
dgA7Kr/IcuywnhqWwEG0VQ6kLGtuZB4qEDvPziJPCB4pK8a0UCbGpKBx03e688UsoDL8JJ4o0Lt/
c5MLJhGNxzglKaZuc7qb/M7pHFkhMOizIxK2pL/0pvBeJlxmnoS9gFCyjZITyD6TdVUT2mglZEYY
RAuD4TYDx33nFv091Nlp6hubuwecQh9AvnUdPb8eEJh7ikP8M28mtQq9qYmPh1UvgoZPXTY5SgqC
MhTeNijVPHnhGPpLaLL0O0TbrdIbRKpvwdzesI6uKtIDIJ4mULXAkgh9ywbdQ4F7VoDj1myjJMAl
wvolLiyp+jj0e3jbznbVqKWCF3GqfI9T+gKNj36GwKnIFD6HagK9L/8TE1VnKyY0G7WezzpAm3ob
iS9RxOvhzH8TR+MTOrScsngsZGXLBxXk3TExbuaqvF9QNiosBI99sbOk0aQDGx8KC7vBkL6gjQzw
GSQGhzP/oIJ035qT6/aa77oaM4sbWuH4tF3oEqE45tO9p2niR241WA5WigYqrQA9MAgASAfXsKGH
iOfs7t5UNyCOCykTTE6RR0Dhhkd72ekmBsKFiAnrENclhuatQeXX+R2g30shwL8XKsyL34BtgS/1
6a1eGqaNoSVM5CMgZ15+9BjMZ9bLshcHZGcPesVQAnxsmWET4tyJW6pfjl78K+XP1iw3U5ONvyK2
mFoLhAUxGFzF7/TzbtWmyBlJX/u0WAzbzQBkpuhcDIoO0VYaZ8842zUiiKiAUprJSWgFJ7MDNqJn
n5brAaxqPSzFkEaRmvE1Xk2OVuhXYoaRNT0gGth98+r/XsRlNYaBOX2ks73UICnMrY9z9xsFgynE
vCDKAaNGIBccB5GOG1yYPfa6db94YG3nUE9k9RJQk9VjAJyUFFPZw0xFIGTbQnoQ+PViwARyziwu
Nt8pRX5GprAxIb5TzUqBPvRTJoss3gYhR8STJyf7M3mJtzN53XSK3z2bWSJ7FUDcHjTkQeIkUMet
7h0WAk1aoTkd7IIy5T+nkkeZ/ms9TnfO7Vc31vVVkArFAsHWtJq3S0sdGsyijA77BinOb1/8C582
iniP3UI1++wQA5FND9TG6SddjwByrGIyLSYr4AHLZFSn73pEMKKaCTtJsVTcRSr/LcpG1YNGPRU9
FmPn7ZSRFDxNvChsTF04pKoo73lPj3lK3H07naT3lICrzhY3VQJpaeFhSy8Psvj9DBXNCxnZeEq1
YBiT3Gt7pu0woUSK0Vmpi8x4lIMSipGAXFRsd/tcEbl11mVeJB5Hfide1Gng7cpU2bWZlG/fDMQH
E1eIYCdY4wMhj3d33myxmTTOvMXtRJ/NjR/l4553jL9keSQuxd4+GpJBhbCoqtg2QlTyLP/iIzJ1
7oW9sQJIfpnYAPxpZSeokVsoqHF+nz+iA/SSPU+XQ3Wy1Jjvq9vwRQ4UHZptc+K0Eo/3mZn8nsPx
uVjwhMEJYmACFH/RceF0oPd2GHQFVjG/iakrantuvh0CuORF12OfdHhYKqNpnXoQyHf6hVQn4QDe
NWnhWORkvzSm0ItJx5r/nF41nm9QXosf+L0CCyvr903gvj30eG3a8pHzOxhIAy4hurJ2lDHcG8bD
Md4DftMZ/8o0GPoXXc3Eydl5d+mTvOOG0SqgOLoNFu+/+26GIool5WxQNyY3UxYJuJXKABGaW9bx
Y/GmEvBSaMQ8YXPyTepnJGh9wKIPrxO1xt9LApfmnJhAtMKgUPimmPGZnvFKiKkKP4wq7Lld+O5T
7ZxEQKwIp1RnaVqRsADqTcUaY7cCTaE3oXP3htEtbmYW5pgfLGAUH7z49MIbEVOA6anRQec99byk
jQVcTFKV5yKWikUTQ56ypR71QbKdhkegYWAM22/iBbM4gWlJpsKpXn9PZdv/f11SfxrICSoPZyrH
NhguBQz/FPYM/6OpheKZvn3xcrUSVUpRfVsnjLmMa4iOGv9PelU/RO5qJQLDyrd7gbEHlWoSfaKc
eDee+jvnbTDIKJsUUXBTxWt4O3xevsKcMDarT9YmkrtNcWO98u4Edk6caGpq/hjT+tZexXGa5Dda
Y0nPxcIJwR3KYKijYPG/Hocbr06eAwosm/oSYPltp/42w3Jx8EhwtVUn/ouH+xvCAz2JysqcMtRM
IWHoG/99pgEnmDXi8Ts3IWC2J28D6CN55BTcOqH1Vkw7SjciJaQP3bQR9ckwYzqIxeZgz4pkO5Ur
EVWfai8d5yUqxZyDe4rxgD4ZwZsfStoSsRmjHI1PMnHY6GSZuaZKmsdZAGQDPRL9uEp+XTr/9dNL
ZYUAojtBDz9IU3DzAOuAF0Austq8KBGZo+jPZznGXU6i/myA1kOK289B63CLZFrDPKBuQldq7XRY
X3o6lnexmnPwPBBS1wxfW7Pl102jXA3/ceV+GfE4mQOEAJ8WUA5aRsWGlTTKtMxwHwOGy/p3v/Xy
yVCOkEAD1drh0Fa5MGPcZi8+n+rgB9QN83aqG0d30OV1cGPYzocVm2sRZez2zuCkvC8FAzl0FYu2
uSnyXe7WHKPKcQaP7DBqlajmFlk+yAn4U/toVroHz7OiYulSC8moQEPhymXpgvtmWKI8/p4+JEOa
kjeLrbZfiENa9lQA2Sn83tmTrQ6/gB+lgWjP2xgjbYR5GVR1S3YUdS3k/qKXYY73u0VztVoC8/c0
47VnsmBUFUzkVnJGhA2CIFqbMzzDCyZr98zSm1xv1yg4CCZgGvOF++k+jVrWBhtSjE6Wv0/wPdjo
zVJ9dBw/AlTdxP5dmqf0DXpDRihK3bKDcKCw2JzDtTh3tpgHyRFkn4UQJSty+GMQ73xjbz6Xo4iC
5KC9Yv5o7Ir8aMDKAd+YkXxLTv+74hR1WC51ZBTcDcu/dtkATXmqM+4CLmFJtpzvYVaREza99bq9
AXVfo+ppHWYzWyVeT2paI6N2UQtFd9X4uGw1TNO7pcULOC9TpMak94n+iT3aQ8KK0id6cyqEndBa
C1SWhI8J4xukdw3zEoiEnqbmrcaG0aH/FFpF1xWv9S9TYleYoZ3Q4OVcA/92wQBpBCMO0eZ+hKDh
GVAUzAG5I2sSZ4M3kMiCRkTziQGc9cfzwyCNSLmPrpJPzg5K6z5AAZahqXA/SO6Q5Z7bAzOXBVV2
fqnXIx2x0m80mRJ8jRaFGarZzvMVD3a4jva3f10U9gREmXDi1ybVg2Ljr12r7tT6GDjsju8E+dMk
2GfImkRcMIEIRabs1SDQYeE4JaIuvaZDjYHcXh2TPcbPJfag8S0nSGu98CAGDgbfQCB7icwkwDk+
CgWZGE2BcRHxbsJdNVdMCvX8NVfUgQZXvGVaicIRAD8LeKg4N+UbchS5fohCv4lTpSETh0fi9UI+
HmYHEMm3nQsDe0uyUS6iXCUXSNFUgZe6b0LdPmPBK3t54pXvypV7L5S7YbBrVa9M31FNHrIIKi3m
0/TxxZbg/cbrMHmC8cnpm8NK49aSbuS++Ule/rru+lFaKr3BraDUVJ/aBTWcVEkJEsWMnbY4FOBn
ZFsVbYFiXTIz22/uG6LqntYOIsMIj8Kwu845tPHmznv92rrI9fCS1oAqoVy6L1FGwFktX51tdH94
HG03t5Qr7r1y5ywNOl9DSSijv7O3XrkoLNILTJJWe0WCex5EDSjVqmCagIifC0FCROhTIBt8CDFJ
PEXY9PuOn6l2SDUMbSO+PTGOkBnHyvfuvhIZ0+MAyUwAypAeUGwe6+qevoshAbNRVXx9y4o4xwM+
yIIRJOAtaI5S7vPttuNY0FCNREN+zpxBd+tGeLH/BIYZriqc5EqB31yr0UCxjoaL5lg16GLes/QC
h13xVg2MNJujy0NnPuGMKHnPcTPi/MU2hKo0/2aJ6QhWsVtzbBnlQuxOsbyWyP/yLJ4NJYMj4Axs
Cp+I1egXral2G/HkdkNAbrObd5IbSF5E2qLbActUUYJAG2U8t5Tqnfm0wVokjcaRmKzrJ03va42s
pCKjSdPxIbjX1NoITK3LqjjONXUFvstaJu6f5Qd63Jzg92T8VyDXF2ydZudt5u3pVd+YBVhToR8Y
AUN5OlA3eRFSa/tpj/JTu+p+pYXize1vetEZD3XqmE2VyRmFbNZWNCKAKly1/ArAT5hX4kL0k4/U
k4yO2zOxWVRFknkoSqBg1V5wEZVkZbUcCVu7HuKmLENcNDnsPYR2aLBkPrgA47zSaDGB0ODUHhXd
OTb3L53RmX96X7wjOkSzT8AEfEDslZQizNuhiHGSQ12OwCBUidrY7+MUHcctG3prBebEXrnQRKEe
3yDFMvpKfdzyyozFg3NW9LxtHzC4fSor76tcWhPMP/imNmFTMTbAHtujM/tiumSNgJyYey8aaYaF
wCFPJpHwwm7ipiRM2hcponAEpdeQQ3MaaYjEQacXm7xh4OsyK7b4yzn6vyLJbfPXd1o6VvgFWgYT
aeVY5fVMbIduvt+ViQNZ6utmzGyy8dGalL7ml+VuJU2DBIHkbShLWPQd6j5ni0lC7GtzhI8utkkF
Fq4T0o57o6fgnXJBcnkA5xcYvX1kn+NEVaBtLm1DbVcIZ2WtU8OFlg/atzlMwJDcxkPOqPYAVaEi
REDO7LwPuPjpGomF58QIZTyGEpgJfdauyp8J7TWGNs3prntGCf8Vzo9UFdqkdhGqUqGFQITlUzQT
LrecTqvUL8iiWE6wSlBoDREGpQ+Upinhohb03uOva9kIzGhg/O7pk3snq2gOMGRmIIcvjz9vfQty
MJFTMXsDSVLKWTJYHYx1Jv9Nwm8GTOvzdMGoKYaEdnSzw0W1BboyUrGlHycM3+b4RmLZR6uFuluY
pvihO3lgIa4+BMdD93dHDq8C7TvPaHWc1y8eZPLwxZhdukt8JmszVBzewQcdqiZfDoj9gO/Ja5V0
o7hjmEqD8oBOKWLfFDJJS+mglYYXPljtg10okPc/GVH7CVp0xMHl8Ut6rkBJYYo9BSB++ZDEkpBb
Rr45b7IKa8Z2/Iu8xFYVoDl1r078FNCdPH0VO78Cjx6PhUim4+ZYz+xknwqKb/TDZsl56y+ZvVYY
YfeS6533ogVT00A+XH2T5qjrpdTGJ93lky1zQhTbNxVTTyqUL8727RmgG1589BmjARmNBiNzQwHN
LyzYzFZs3r+aqtC2iETVnV6k/1L5e7pLJQY0x32Xi4+S90WUuINcP8Khu1f6BpwM1nlod9huk/ZV
KefETUEjgLRWA0rcRHZfFKiWsdOr9leY6mpaEu6RLkFLgM8oTjO6mQ6E3kDXZyKxPpZJ0Arm3+MW
cxBlmVyAwSfmGTX7/HDfFA8NziEXejJSbXWh4ALmdqId2FpgMNHAD/GPyb0M2/wKSxCfHGHaBqx4
bFFwvKdaI9+KKEgO8x47An6gBsDxJE/dyvO0tHiuviA6bviYINHCog8m1xRXd90KIDXOBOuJUpSJ
LGhuUCrewB2jqxavwKkthN/UWiFUCrcRA7R0iHH+wbr56ftqsxB7DAslsZPlsARFBmeG71Q+aQzT
Jloq5MmQBNymYrSqdW+NiJKse0toOcm82GTVK1qauOIcatfTlrHyiNiMeCe3GzAXWiACAta5m/E9
5n2VWexmhYMOKrvemoiABQ6XlpX2aaawu6bqU3DgiIoJ5thA38f6io9bd4XApQ+4mBVE0nRoTz5x
I41usRF2/NqE0W7nli3AXODxvkO0UttBJUSMFOQCDMpHEuDJ5m2ryHwPj9lRYIb8F1u3D52S53Eg
fxuP+/kDoowoqEsPf4B+1YmcqzZgU739AtTk+Lr5l3LK1+kee7GYNl/ObtiRho8HCnFshi1XYKdQ
1GQ9afqhQ7VGzI+GiLC6xU3z12zkfThj931MHvyayHqkQyIrPFFyzumZgD+0fbn7OU8pUxYGotJO
WsVgZCCuvvpafnx5YwkqhKL2SiRD20Vqz96VVkAcvEDR00W/v9VJe6G5Ok7slX+oCCNX8WE/bN0W
OajuIs/DopNbvZDFni5RWzByb0KY4CYFFybWFVJ4ebHnXaPSTTfNXztFksvgiSTcx+Y4i3IsPixb
yihZuzvyjQO2nYmmOT9BdIfF/6MbboE+3B5+g7VvBAeSwKwMYoad8y6rm4UsZVhLmsoOQW9l+JBM
N7gfACnHRG6ExZGPdG2Gel7xQywwGsPRCWT+lxQb5PtoewcEsXhj4BMsGZQCoTY/00nU1lRFwn+0
ofp6ptiYjIEbNgUamOFHzT0sOr4bGqiFcMIKcDiySA4UQsx4LdLWL7myxqftWOwSEMJrpSjthxjQ
x7KeSgQjmZiJ2menrSyDnzZ5datqwzd04jJw/kl/rxVnw173GZkrvS90S5M3Da4SafoocYwCDe/x
Ryvej2YwJxD4DOU78DGZqA+dgzXR72M5aOyGAg8kfckDThf0JOXwmgV2r5L/fyvKSveCCAojJHrp
ZB0LFFBhjKXDzSXSuNru5BNVJcDTXVHsH7mjZ7Z9nBQk5j+CSL7kJYVD49RJ+86E7qwf50JnhdY7
CO+azH31NDOp8QvZnbd6f3hlqU63MfHC9Smzmfr/cU3697Fepo42u9HWjDgwl0tLMapO5+tbgWzz
YftKsmzDdcgXcrdmm/CvbJE9vMWBEdv8lB8ZKgxgOvuJ9VEX63XF/tQJw6+MukKcBan75v4WRFow
TXaip36r/2tvT3zz7c4myQwXBwSSDwIxwoCuvfmjPTZHePBsqNYofRdrdg6VPE3KKQJZ1x8KZRmH
8M6uA3t+ZPI8Mccre4D2SnxT3h9/BCqwNwrbiCq5GFg4CSzgFWMvJVSMB6BXv9sE/avRr/yTE7AG
zrasylE5HX0OgHCfb0qPXpUV1qGfK9fPZD9sO9X5VZGXPd9yT4rMmbHhdBCRNrwiKkumidviO6LG
u06xvLzofZ0221uSWE/sF5ZqCiQFRadU+OFoXGEz60SROL22B3E/fbLdRhVhK2G8GAy9rsfKWyMy
C6HJg52TxLUbZLs9RECcgHS9m8xVPc0wIlyuCo8yR1T4EMS1un8lUAI2scUoXy8eh7skEs2hpvHX
cpiUQUPNIUNyKnz8uIKxdiZNrHq6y1XrAwYdsL9jSjdznmdcef7b5id+fda+05TSmpWmEqYqeR8w
nPzBWNWGVhCS+f0Sd3KrV5Esy1MdKfKwcetcZukb8F4Sj9IS9NwJamL4t3o3uAjWyc8oZMRsZzMk
R8OcPazAwUSdcwvtkKxk4QSkLrYW8n4dxCmDuLXUWDGb/okiwlR05Z5A5vXmJIJ4/tEwxGGVu4yE
3i/jf/90hkGKrWlUiGwD48A+NayX7+jDaVacJuvEId0ApPJ3Gnp9V19CezCfsqFfw9qcWcqEGLGf
P31fTUldeWUBf//DLcrDzXBxR3bLO4Rbutd9ugDfmwiVt6A1AOSjCAG2yNuPSmurH55Bkb7aGkcw
WYNWRedz1Z/DCCXjSdAlkUdmQejT8ahUrN3RyXiRQP3uTtffMwAkoU8BNfW4gZsQVL8SuOERFKm6
4/uBux0mLR4T/MBouT+88ELsMhRLM46K0/B/t9n9WCJlHjxMpuoBd1WTV/VO3v7Z5f47Krnog/dO
pmUyJqEHgxtBCGPYPDGh+wsvoPehEVYVqS2Uf0YVLiv5qCgr/uLHIwaUuZQuPtrQQr1yeE5VJas3
FWtmiUUdNTbiDlU24PM3gzsLof5eBWfC7cv3txt8NpqrBfgLxP4bOl2qt1RnKkMDLW++kQ+I/+b2
TQDmy2GNPCDagHcMJs/qPslWRb1fugKIb/3mjCcy8qacr/xmYCBPSgNoxVkChABWuvjB6gf5CtKV
YCrjTkk6a1mMEnvkD7ohADRN8LPkrcJzDMGg8hnMUpxe/r15RPyuGzCYxGEABgk8VuKX7lxbfwlJ
ktnnxYm8b2RUDrZ/QvZH8sfs2k811DOZplRw7SVG9o7RkejmZSs43MklA7a7s8U+pqIbHt4VGVrs
dYpr8Xpgsri6A1pQioxZGdsV99xcN1cARjZWCn94DR8ZQweDEoltib+k4FDlr5TCaWR/aygrwgxR
ZXw0tqvkte9BnIDR9+Y6KgJ2EDtsETxTVErNF62FrwOxo0gzkPWdkXIB2N1g7NDdVlpNCZdlHEpA
KfUFXJyt4TfAR0fsImv/QSf2b27s+oP3Wgl7PjKHcYr08RZ9OIUpdHUAOrqB+rIkL5Zi4D6Urvo+
KfKMz+cxi9dZ8JGlUre/hNGb3IUemWsT0e+E9DWSNezQJU2zjs3HsTZnp2qepQhMgDGd0Hea+oUD
P5BgmjJ6YUMegjuKv5X80mJ6SZthnUxTGRa8fROHwFRvuPBsnDb1stF4boK5Gnhro0A2VwNeJrAw
b8+IDGz76ic5ZDRC+gyOzpTuu4d/SqRr6imXWLCt0p4CQYkYkoaq5D4gXpeZ2ZVSvw60Ax1DpEmq
2MNhz6jV7L6utY/1RVbrNSzl7Rp6BSfwvaoUCAI6mExNfx6IdSH1/y0/f91/kVCx/xmizMFeM0LR
miRZsjmMvBfJg/1PsZlLG+Ij6Of+orHKnvRwM4dNm2JjYE+R3Vn9SBKBA8YpA043+z/MTsy285sJ
dq8fWlSbUpv3xE9uOTTkvmdbAvmv7UQIxO8zVQNEO1mjdx09/qgKEKctF8L0jdKi+hyd+DVBjDTh
A3U5iGx+Ekf0EdxXOdG72tfFtRZijUUqG5H5ebf3cbDm94fW8PFS0m0ocvyp7tZBT3D+NwkheygF
fb25S5GenAgs+bhb+5fRDyOoAVoesq0CwjO+iVvcyU7qGPgL7zz79ylSmVW9fZujpbko7zwTeCxf
6iqvMWnTO42DFuv8gbcglBpaReihW3wrb1ssf8XLRvJideeyPMF6lUjeOuQo0PYefX6M6kcOHE/A
7jHPsQEjhCCL/SzwXYGiVgd3wGLua7m2zHAMALW+KOVii+SZjGDFlaAh38iQOR9Td7EBkz3G98nQ
j3UwB1HhzoJM8BDx0XWlzzuVtT8aJ4wUuFbXcOc62MeotEN5px5Yok5EtnvNc0IEvyd8S/ZgVqFW
RMkcbXp4ehtnOFoXkC3FP83v3fmLZnL87WQaUzr6YQLuWCMzQxm642xGcrSirG3P2L/iBmQQevWq
2h4SlHZd0K3TRcJ1ZIs4BiCz7WeRjKP3DsmGPzU/MWHgxpt5awVxrOgQPF4z83ypCgahUfiCv45I
iznb+WksNUAGNVTCWj7BJ5ugE3vIN2pujg2QBRoH/k3BzCqygWnku+cLX2F1mvyUTSq0Oa/bNUDd
U2vvaRPHbXwj+jeai/iTjxhbfx11NTLZa/zNCugvtce96qSn6JZ/zhkUB4KxqYRwIOb5FeSaQa/E
p2bdFBcYUBiM7KoH/4ih24EDRnTQDXFKUh2MMiWXCiUo4zMwTbCGCci+lzeNH7j+je76AzytE+zk
DOcsMlbYioLli5mwY8DW2wwUiCDso6biND4QWufY9GcCeL0vKtMGnsRcKgpHhOhrOYHqQQjBYkEB
tu9P2vHTsnc0fetCs/0K8OaLJZq1eTdDDTcQb42XVWhBM1ok+FT9CGaR53CmOmpuoQmWq4FSp4Zp
h33D6S0GDjK7Iw01meuLJQnykqbPwhsVkzHWWmiJcREi8I0GsuGbzhUSqkgLC2OYfGfra2K1xG94
+D9g1Ufvns7vVYJbjQIV5vrC4JE4Jg4qjn25BexeeD5BcGHEEjq4+lCme6BccK/CyonY+mwNn0eo
Ghps++FefGLAoxnvnRQtYwhdJCsdeibzFdh9VddXuydF385wWH67hXsQY9eDwdms22u23VTJpRVT
h1MRoGyWUmjvzozF4Q6qIWaHlP476pl6b+8ebFAKEJ6DtDB7T9paaR4WuMPKMpAY14l0r8TDzUZ8
mY9VLdKPfZzUrMZOs1GjTZBjV9YC+pszKaSuNtqPFnflLplysQFS5Bik4HwlxrIJZSJm8GaeSapE
bnANoH2DGp9Qqs8+8IemueNTjJ45p3WRlNOPZbZFOjCqxHUan2d8yJCZuvDXbH9jMT8fjnGRM9QZ
I+dCuzZkmp2fbO5TTYBfF44N2o1oXLmejLh/iYCU7dyzBgEextLzUCWTchlgBPp61Rjkpiq7HKhA
amcPLXABqEZMQuOqYU48sud2eIrJY3kcmYvOcfi66C/HKT4Cb1wlRo1wj7LeLoqG+RaX+YkrOZk/
A7LJP83/16TkDZlwZjqnuH3a5h8m8mc9PaLj30oG0ksJ4cKQslSgoB5YABb8qBDuj7RyFkDXtOSD
bxwGyWxGIeg8+evNIPZE6R7VIeSA07UU3ju/JEUh5SMU2XaqMvvSMCo3o0L1UXRe7Ke7IMqVqoih
VzzaU0i76VCE227g7xwFQw9gJr57H1ImS2nK7TsWoEdSa3ar1lLAOMJkfR+XThq0Uk2R2HUAdAHn
2HU5rZmxLgHx8rxwa+CdFlZowwkOuMWmczv2R7Cycy6EjL/L5JJKpA7wjtidmyyGAWKOxIcjLUxk
qBYfuW8vqHBUbef4DE9VdlzMa424uTlKeLL22TTxMT1vMokaLg3y2qoFbKAilILCr54CChxGRB/S
GJdMWfO/M+zTb9DFyK9gtWXC/6FIFIO9Xsp14AzzccpbbluiJB1irpMtSwsvlVFCtUvJNrXF2Zkn
p0fp8nfG/O9WaMnSrAGtfuZ77IJA1+5ztYJ9/L0xFM15uZMR/kUsd/CtT0IzGhmxb5c47aIf96jL
2IPBxBJc/9hLTcBTKZ2dS1igw//Us2RItZN8YvZ0xYR1Oh+C9q+HgDvRdPwtQRqHtjQOg69XzESq
BKFMoAhhVg16AWIN0Wp3ZF5i81zRkhuGVE4UzY9XMvvXgCZUH6aoBBwIZxb1wrqWCp69/5/yDCpr
l/NUMPsQcppOaYOsE8DdGmAz4EMEIlFv5870DerxvD/o8nT6ScJMAFSPs5SCYgQpoUNTrJB4t20b
lyohGIszmu0WBX3Bg2nzakaYmrq8kW0RTZbI3JRNHPjlhQ+Xk/dui9urfQpegpdtM2wKYMvmVWJu
R43zYaNy76gpXHKfKEMoaLAz1+9iUMfk8L/ZJ1EvkObKwaoj0vHtauhtt4Dmg3KqQIURQRf8vy65
w4CqXnKm+MBGvhcwA8Fbzp2HOUowIT8WCQ9ToNKsodwcU4SKVHxLi3HY2jt7bgxYzACxNbCYIRZh
zUQKtecQx9GhCjzQFVIXYHgbfPmljVWwUGjMaK3LonaOKNzjXeT72GdrSo3k6ql7Js7oRJOPvH2P
ZxwhPcDwLCk44yVTRzQwckUYGRsaTBeF3EUS5E++xXzhfL70t5fS8564ZrMkwIi22ugZY/J1k2hO
Qp97BRow9EcxkVWGu+Z75LhUXVoZLu4mVER3ZuA9ugTH5RVJqnpHrnsid2EPHToWaO6phJjTJdlE
etchrF7HL2uF6ZSswwi2uxnhDqWq/Alfj1gB/PHvYf9JQNdF98oYIJQ7KDpX7rDZeCHWfOxgHAZD
NORcgobANtf7UWsXyFSVMf7lEueNGZNQBsvo4+8tflhKEEWsPxJDp3/P1pjRSn1S9RBrxxqkWYSh
XL+A2OGOUa2TDZF7ATf4BIfxScGa/5l5ShwNGo2znGjBLapM0w+Rhy1HwiGR6xwhcV12HCyn7H9k
KC9JXAOhs02xmV2Sxwls/FLAQPzLk1pt6EjrHNzcP+Nwgfn0o7MYj35669zXyrwLW5aHyGFVeKf5
CSYgD/hYrIcvbaN9AxLzP9LljtGeNdB977cmCVWloK9LL07bcWmZ8Qt3CtOqLQniKs6Ugzng4Hu2
511fjAbIy7jiypAOR1KGmTYftvIo7cRsUiQRgt4hD5+QwK3Q5PKZa39G2B1k+wkUR+DuDmt/kOEa
znqhnzeM10PL0btJRCpHlbL0lfYrAMO2p3HVCQStCZg8y7hhp64RoUXnZ32nzOLMqdrgSuZBs/Nu
eFkFnZO3y90fTEZ29TDgLNW5OQssxVjbtkP1S9IKtltixYOvzUpkh9x775/DAxyGkxScbCvP3Xt5
pe0agUMASkbBVMBQkxut/ygs0eXmpbJMbAfz+DofFSQ+iOcUm1pbv96UJoFtcHaaSF6WfO3z/KGH
2tojtDu8Izp16Sl7GFcvhcwBlrG3jTRAny4x9x2n5lOPb2LlMOu1Fj5NX2GIReS9eb7/MXxEMfX/
CPfKRGlCSNFNMKh3oIGtK4ASYUmc8UgSvDA/Epl77men6U08SQSpE5DVgonftGD/OD1zl2w9Ci3I
2MQvSnUA2kDhuNV8f0EwzbVrwr9UzxtbXMi66wps2OhdoBcplK1xLQRncgxwNT3vjmZjtyZ9tMGm
sUENkRCqyUZqSkqUjYzOXar3vTNGWuG6Dx80v4LIebQL2O1s/NJ29k5Jy9HKbgxSIxabpmBqIL7J
GPHl4BvrHsS2mn65hMCTnxBog7xtjPEr5qxB0r0PUgh2C9iL3AWxalS7l4KUswZxUTWqrCozCFUp
pv1yeEXsWSEjV1GdtbkLASYYRXCkLOJ9ARFS1ymczSHXaiUR7ILxScuVqM5230rzFyOZ7/MPoN9R
mWg9sM/+K8tsLQfQenDjVjY2DEWqX7MWVaqpntZBgXv64Y/7uSCyZeBERfqNf5q80RPnTGaTkvPl
DTrPMI4eeYGFc6EusnOAjWMR/4Rf3gCyT+R0Z3nk0cPV+ipX1/V/MFCum3+u8+998k3z39OIj2F0
gCPcCBGaTMkyvj4XTiKONseASJZQ+SpXvKe99mktYmGxVa5gJkNFIUvUymiYfja7zTxu/lcRXqRb
izfh3aJ80UPz3hhiDi+edVpK3eSB7oKeG1QMd+IKDqrDwxb60b6GC1SaXfF6ZYPzKqLY1TCo79uj
q35jnspOGNvtQnxHXzdCBUaqoua+PIf8+b3bsfmffG2Bl3m+255Z/1qC8vOU2mFxTHKx+j1WmPER
bRNeniOqR5hewRsufO7gtuBsG6OWWeIYlWP71qM8qd+FdRg39WhD3DITNF2o+wQOz2WWMgQlcYrw
h/QFLZ9VmL/bRatmXdUZhcW6ukHy+hwVZTXSXCfTj9TZMYjSi3Cyg8NMSTFIH8MEXLvq6Hn45797
MI1+SX0QHOjizB6cofPoIg3oaqVlcFMvkvg+8zkk8bKXQ8eTydY412tcf5KHz4RfaxHR//fK7jza
dmVqS+//ISTzn5yp6TOFSYVxJJw5E2MQnW2ruHL2Kes7liaog+Mp46KjqiY2CUQFd14L2Uu3ImVH
4N32dOgilFKWsDlGDJAB3y8K2woGj4OyocK++5fKbc2zKcWrIenX28LLn9tXXhYZ9M53FWinZS3+
yREc/hUDsJaUUNt2j4jPBbb6oJm5IipF8K/alfijF2vOjhclR6dlVzWLnklhySKGStJN+gzTHJUu
jXXL34eAOopOOMRg9hF3y43rCbbJvhQ5MD7LmZ5auQVJw/cxPOJzRY8rQGBEyEinV34wFKE3/sWF
gO7wIOLQoP1wB3v67XiZyHxutHg24fRJkWGur13i62fhEtz2cid1DwzwJDOwGtZWgGa3yWZzBfCn
bRZnBD/qDwF1aYkkhrUxHG5jqF4K3cRjTbY7DxPiQaxHWosi1D1ueiP3LneaF5aBPoRD7oWDFi40
EotOjrm9yC+UYwIKyPlQOY+BO2hA37j6ozaewZilb4ahDlQpgpqDgadoqx6bjqZ1t3Y2l57LAro7
1VM30BvLMH++85P0WmQQlgVZqyb8t2q6cQlE4JoG5eELsz92DcP+HAnQV22P329UdboPkTtGQscq
y81EIAIJOB6JeghMpiZ3vRB26IFBEPmezRd/CcaClnHIGypZQckbLhCY+pfpJhyMHMa4PEHzlmvn
MDbrPqoRgQlN+QgVgs8rxApjBi4zBwhNcfITuq0fXXmqdUiHjL0cyRA5xLxkDEqH4cfPVpqODpS7
ilensOphhG8TPDCLc1TyvwJQcDwYwwKAfV0ptv5lkSnhjejkAwsLhp8tQ4x7khz1CnD3C5tRh5Zz
eBlokufIQ35aK/EmMJxO9mGIBg8nLPcJoCQhFR83cCKLrfrsUW0qmN8SE3Zo+nIcM+hvjxd7jaiB
hdniSaWqzyMehjCbZGvijH8NlB4Up5uva8jVWRSVbtqyvw5QCRg10rJySwYP5FnuUQi43Ta/hW5R
oFE7TRViZDhFAv+T1WQ+B0tYfwvyAhjf8rtw23k75vWA+q39TMCVcrRHItdO7XrbBVE1C+oJz16x
PTuCbFmM1syadr9Ewqq0Hnv45UQQKeOKmtSqTsoeidkkQOW4VZJAMVWI573UJCG0ycrIf5bMk2bZ
mEqPl9aDkhh66oiauZIVSV76Vn8KWzNMyEONrkAXHNtEjEvcg+25Sxd+yISOx/JJih9HKAvP/2LH
ZyPZQJ0o5f3iZ46sDvfkwPEMObYXSGwV37G+CqASL3pN0hfvWflizleBeqS/fFcHahqlUkRhU/cC
zE+B0zZZajxzhLsnCBALa5a/wQffuivXLtCYYWWG5SHPYHUqw7s54EQqscjXly72jHML/cNYPhi+
iDngOhSDXrFmNFXmU0NkicUafFrn8Qe/dT8l1s1jpgYyX7Dsw+t+KwzXOXCAsWVBUJISqRzGDTew
Cmsu1RejUpqmAaLDO+OdwlVQCnLoN+vNfxd1/sqGWySMiUWGdaehvzDL/0oIOM5CSc21/t58jiG+
n8jJiHnOhEE6CxiuwYmNo4Y5eD8lqdVcM3VBn/x1juluMxF5YKEtMH65+FsH6lfekSO5KQWv0rEU
JzAdMZ8tE5CxVUbL4tD64sWG8FAfAL4EVFtFTGKhkqgWndOecpgU4wfcsCxpItAwm2zS3AFHRr8W
9VXpx2RSUYUXeWp9QIrSlM+B71fkwdIkxaafomr3fPFKwKJPNgZ/WJHMCTaftgrAIKKm8xFUvq2K
jQtH77XEpiVaN7XP4OV3Iq6VY/lbZLExC5cYvW04tQSIekSWEgctJqWVOf64muY0i52xBo7zliDA
xgFZ7f6SqmvK4t1gMMx5M/d/THe2361wrk9sL0tMVDS+fQLBkH43z4hWJ4sdgpUYxum4nwDfrfQb
Oi0bP8HZMmSCx4GO+zXQfeZWbRjrqZJOVn2Lpc405EcdbcBOZZ7rpVo1nrl+45PUbcpcehbKVLFG
k1CeU6GQgCaT4ZeIH/QJSUA6g59GBYUl2llf+9kqGAM32q2aJ0zL5ABovvClsRiL/SJ+mp+Ve7y1
dExvn4sXPA2XmHjcvbVcCuYLudr/wl3xCleC1DgXhEu4MNZj6EvU702pKX4/y2bWX9I+N2EDwHzK
YLaHCIiTkHT2L0RhP0CIfCYcOcqBDX+DeuepnoAH8bc2koDEqvR4ZXWJiPZqaoa8FUFqDlHD5+m8
/IvimqS2DCwEXt58mr+Lkh9sna5v6o65017wjOFYsTFA0/ViIdN7chLp07Injg749wkCaW95ZGrT
k9WGaXf5W3ogi+q/gEM6L/Fzu/EG1+7KYS5oYBKFsOGXvq49pYfUFakvatj03u8TBPX5ij4kxF5a
lD/xXyF7WZeQKcpfC8kIcO0LiG60nMf/uYK7dOdiYNTKLMPsUQfq3muhy1j4KtMx5YXmCaqAAtf3
T+XVmlexv9SH1lh+fMyJGZXOqzmUA2cFQh0CXhU8WqsrJcHhNcuYauMEavaazA64Zx50GJXmmJIV
Aj6X7Ae8Ky/YTCHze2LzwIyFxnxxN0SiMGPEpGIFNGadj+Aax6yfOWwM5pFco6Ej8g273y7sYkle
bKboEiDQOAoihiCa8YxpXRNJvfR5x0Zalqhzz3+HWCyE2ov4WSliotvL4QRAkvtMtyaxAGKYIhdZ
d5lunImvsXZArl5YHMxNF0W/8I27+DgSX05WGgmt1ql27YjMqyWg68KANuyD677gNVg9RtnjaZ3k
GlhUQ39vWCvosQ9w149Y5aIQCgbE6wSIMJOYdG/J46JnXu3RbdZL/at1HNnY7P3UYrB3Dvdd6EkF
mYRf7vB4NJgxH4Dhdw31Ozq848J3mx0w8wbTXQxqEBKoWIbCogfnPTbDD51JvDq4DcWm1t+niSkP
NHwSiFs7RSyBccsljDanQJXJI7VTwK5KALyQgpv5J+lLthF2nPQXmo/oMIgxQE4EWRxWAmpDNZ2T
2hdOvUebtkjpHPmkZjugTYFXQsBk35Amd4J5QkQBAhfzl7ZWu8vCpQu4FL4Xuu6CNBJrhMarTMjI
0MzXRI1oChSqLXbd177RVxakc/rhG7D4VM1Q4jEio7U3rMvBfHlkIO1ins3QHmPWLoDHZqaY5DRr
TtUjs+OPkfFVgtNtVXFkIeIiaXUqf4R1yx6+fPUsVdTB11KWUWnsfL7AQRgeXcPiBsbdVXOba9Vh
hFEUGm7A+k58r77wGVIL4nHaJLXO3eEMVAv347KCv2YVzpG++VSaLVrnWYYICmXWWsJXMjVIeEaa
WxFoHmG9rEC570pRajT/MN+h+UB195kRqbxVdkFdwndTOtC1A9zimgXF1w/lnsMgtH472xltR78A
PkN7Or6SPv1+kQ6WWenhwDF0OH1ONm6D1+8/ruQjiRy9DaRLKKWfqXFuooCMq78g2MbhalrRBO8z
wNGXieKOvvPsQRimhsc7lsN/sDwqL5WWsGmARYq3DCsvFufiw9DTPd/PAqMrTt4OUmhmNXxq63Mr
bfR6BEj8+uv7Q312WA4w0lbRYW2WGoiBiBiAj8Y3xRUXUcHw4BkQJ+VbIeg9CgDfC4qwrk2wOHn1
LQbeFHT9XqveS6w58KCxryRyJvYlx2A2IID9DNtmzLhT8KRAuIFIeuBO5yKQquqRM10AS/VvZ0DS
7V1QyjjLMkURwIrXXXwnsxNTMrePlIo/n8ztJjqjoSy5/IYjAv+h0jT+FoqsE22CYxSHAhMe9BMZ
dgNynvmCbXF6kzYVLU4K2seQodrY8g/Ist9pAYU5C+u6vEy58hkYu1LzQaAPL4ypWKK+ar367Y7n
uFyLEDl1GOTWhAUWkGvfEjkA6rgbFL0XXYA7F0tqiaBIP6ZepyfVBgkzghLiIjalG74uAmjB+AcH
qOU8Ot1HrdqNkqmRuhQtyHcfY6U3gk2B3Z3tBAQPObZHAa2WH7+e7FwUQ4rqx4bI3yBwtEdtmmk8
czX0TH20pHDwYs9SLMFjHKfvMWX3lvLS5O5nT281EhRyNixQDcs3kPV6TjeBuxBUlUO62qOOMr5O
1dS9fozHbhC6DQ9aUtipZs5bsIXOv0L2QOhv6FiAZpVUgjA6e12jQGHmws78s6mIORVaVTu9+49Z
oOF2vRwzOF1+OnW5lSAK2mAk1MYyVV9cYOfOjqa13O/IkLEfgMY96GKY8/Ozr6qudoINPKsADIWI
SrlOooy05GgQjopnV9H+K8WnVKVtRSFCxXzMHzn9bN9Wv1DmYEJTwam9uEqfMTgh5JcObECXprX+
SK62YO6e9sEyLuqpsjdl/CVRVQNp31EhXPK6VoAOucPA10K0xKi9kXa2/H0mb16yBGAus3KR8Nmq
C81c0cmvRYK97GuwYMuMamuB8uClVdEjXnPQOloCaX3NJO/iu3VTVNU17LIImpT2Wny7LicUSH2M
BrZAfa+C7pHePx5fsTh02ABZ9oni+m+c3ANOCiPNX1+n6+r3A+/rjWusUPv7rXTowg3wjNl0NzgG
UrmsXG1hgi07QM43jrZTdMLSTWjBHSBfvsX5YMr+HOEPxz4gUKcOJGsUiBQXWLqz9ROSznUIsc4K
or2HqsiqEhN1UcTpBiwdShwXLspNww9Pmi0NtLHgyux5XnD5s3d4YYNWhu54JF8kInHi+TQJu8oB
xEfPFzFwNYUQZtyF08VqIijmAGFMrhhp3CbKDx6ntA2nyymj+4MStiQ+/q0zF5Sj/BrqKRePTYL7
Ry5Wi7eoqKIicX3t2i1EweI99CoHPJldIDvPdiDXoBGgkPRzyeGAo1LSSsCF6FeuMqYCYanspg2l
smqcQetegtOrLDXeKgKHdBdsiousatJ4S7+VLtx3TdIRnK/A0dr/tJMWLIEvE3nYpFWKGKWcfNx/
KvTeA1Gh4toR7Y76pqfjYJ7SkL9z0qweBsuaIZmB3geAwNAmQlg72K86kdMoyh2kRxI/6za3BcEE
TdhbEQzeV9xlTxpLXGbyRYPOsjOFtA7pew5QuV7YE1eh2s4AvxQlsJoIClkuo3KmkSuJqiwptIAJ
4vV8EW3Tv9qDBHF6Ml+aTwTBnsHvQS35eer0k3Wud/LlPjYHnnQ7LKAoVsvq2czoEgNImXUpXmfk
AtUDrDmzvVOAlaY/ckL2Z0f8KiQ1JA2/YdzNF9j4L35VMdEMLJ7IrTSylLlLfU8y/+vPm57Ou2bH
owrFbsFulGQIDMtX0WkTV62ru+U6a/FNlNiHdWSUir/BYUGihRpuAHuNIbAwT/bGzd0vw6dXFVEI
FFCgGtmPIKymwcgGy9V1NL21Wk6OjU85eMqIRmnRfjk8FvLOVpXSTrzSiAFaIYNXokUvdfqPAAvA
GRH6te8ALKC6l7lDMAVACvB0XR25GJEWxtjTPLma5c/EU+WpVueKki2iJvKtkpAx2q0c4BGx0G0t
jqbgNeBFMbQn1nfvhMGj2srX15tdBiiClKtnTyTknyOU5I4bvgREj6vzzVZRaoUgqW/4/crQ10z0
3VVTvRWOdGcvyVSdpi9Wt2Op50vZxE2LuR2/ffOqiLM+f2a8LbMK4a4uzlWObYyy8vKgQezE3WY2
UMSBdn0kIons6okT/I8ajhaHWJxMYNskjuVqj9Xyiiv2iq1yt33PQ2GM26UmaTPalfP3kqfdd+lF
jbKwHLd3M7g6FzkRcE3I5z3cgr4UDEn+7H/XsiGAQJsf+HmzGQDe/yurdMrDAMJbCpSOa5Qqev6v
0ZXd9Yt7hGlM4dFhpxlBeB1ystLvxTNngPRebhbdXoXLxiO7eOed5zT/Kn8ilmiui2YGGnrgAz72
749XZuONlVLn8h/46K8zejZcSf+lf/fCmUHPeUXyczhzC7mIErrVtQ+QwGCjVpWtjx77+Y5fI6fW
1jvBnN8kcRiy5ySDic9eo3b/VPKCaFZWAjhKm1jExw0cPLwTSbliLkKDyTZChrLXOIn3lSsAaXde
dZo8Ko0OhuMBEPaihmLNDxOngiPFXIL5QdDz7XjUW0g1ncMlGoOHlNczcctV+Augq7KiU8GrAu31
LuE+qQGnHFi+oHwV0c78sSK6xgsCRYWP5R/Y0oDjV8K+NPlLWCngJCwoyL2J5lFhFzPteH2+frFp
euiHQ9WE5RCgV0CBpwLxQjV79BgKhekKDxndvG5hWoJA21dS8rH2SpS0ECFUwMNY/ghfGm389vD3
JIx0uOQaj7hnIDYieN10eN6rwL2WYwCgC61tMwyPtHMxoiBEKvk7icyMrjEytQm5JUzvuqBhIM/F
oJspBqgjg164S94pfxHmpeazE/tOQ2fmfLVzP1hB+w6ylZRiC91v915jvPrixgq4yq480hGLBlkH
Ik3fBC3K09Nu19Hyuh3IdyyRxzJFhmsQJaCz2zUHzINHBNf78Re3WYvr4doU+EWLHo1wpjYT/rbf
YKeFXGrJUOUqaZXjs10TOqxrD7vn7LmTBFj52gj5uElUJIodNVeG93zMhSEP8hBk+5l7xtT71IXA
hqTtuPx2XU68au+k/0aoQ8zxHArMAO/SYX7p9WqLrk3yJ1JfH4M7Ax17O834vEIk7COWn8uHUY3v
FXTEiXBHgzOJ6lOhdRLCPhtWiuDG8HWNsVmNlwBe3vZVGs+H0fG0/+xeJ2FdjTKMK9JtejSAS+kq
hTeJgFPQfoHbPqeG2OQfHs0ajOK5/Yco/lMf41hEMjtRfl4uhP4F386Vk/kuKXPP09kILOdGSCFO
8EetkM1kQ1A4ZFA7GxgOZSwREQNPZzCmCjPjI0BGUgJEdZ72KXk8qT7uvlw2AArQI38rscIrI4WY
klEwgsyyLoU36n0n6vRY5JPii0CiP5j94afc+IgLcOrm6uc/AtMCJ6tkC9uZKtfsI3QbGZqGPA33
3cXl+5wv9uU8IbO2g8UhqF17VBtnj/bf77wDo+prE82mcKJsFJfM97qXlhTsmAEu91PmJvo3L+f+
tmyAtqkZM7yPgiuM5YUpwx3cRwfygUzAdgezk+uHPxM/zOyx0Eu/Zs7KGjbK2vj0gHr9vfsJDx5h
mBpOfp0Q6GQvkfhQw3vf/jR/6WYls1Q1n2DKrWZ/W9BQWUrBL491zR6htERZ3bFQIGZD8wRCmXh5
MXLifOKw6f9W+byg1GyoOKf8691MNuN0u7UmpZzX90ecFpIziwv9Y/qRZhmYeZSum8XiXRVDVW9S
maiXie2TA/T6+kyQuuDXyeQoivQbh/t6/850DWNg48VPveAVuSlHubne7Zs/OLK7c8Ry/H3ntlqN
JjxKYta8/0zBR2p4nL1SlYdBNFsxNSGUrwhke0LqkCbqRD7d8dBLpCeibGYQjNOSRCU2UjsVB6fs
I7qrOFXfAHpwj9NndmvHUASGBJMrZ7rvWuG6gI2skwFDv/Xc15vLXMr6M61nzvEZneqcZuCkeCco
5rf+Qda+mNmZwGH8coCOoLddhES1oilsywsUyUuOlHX2Htz/NnXbLeYGbF3F+8AAm9jIPBiO8kxH
wFUDmpKUdubfbB9awoMCRtRzzTc//er3N8tLveKN0nHifV78RDTJbpOe4jJjlvh4AgwebYBLEySa
Guz3jjfQGmOLX+B1nrbnODRnvD2t6Cq1+jdCOWWpKAyaM7k3C2CdtfqffClOcnOv7CxXmg35/pG0
fcn+yMfSZ2b31ye8yiIujTJ/6kGd8Sz6WQat34Bv2SsMf5xnMg4Qi9csluH5ko436jK+tHL85bf8
Cls6vEp3G12JusOAA0ZjTNdUd3oHtMdkZz2len9BvsVz+yA26PBjSf9nLo7KwYe36yqxSAChUV6+
m8mgKsC8SPCEImZ92/m4mI53fUI6ycx+fxrq4+5zk5hjqNpUxEhdikCK+2kANsiZqjyugu8fMh+c
RrBNdzTupPmf6++ryDEj2qOpg+f/ZsXmG48mJwYqO6Hc5Db4ReuJgLjyyhqTCyh9nTlYTuzxtsLr
ln3EntUu6+o4dLxVnpkd44cx4AFSicGfR3zqPS1r+AFXtKY9X6mNun3YIYJcWVU/6am9XuOlWJOW
HsafMDLOdDd/LNsG4ZoNsNzG9qRSBAocfwZgmOxKUrMYAS2K2uRKwksKwUigbsiJJWJ18AJPC80T
4hk9mhPyp0jGwlR4DaL2yl0UVQo0AhNILwwpQQrARa2j3ji0zyym9CpZfpbmY+nSY7GJER6hKyd9
CO7y2yySmKvN+ITJxJvQmxet5dKRyXv7kazpsJbCzrgaD6n2MnF746S29+TL+L43//Hnlm2Er4lK
1J/Ii1U/X2ufPWAZ0dR/dBPW2oujm7t7l7NHdp9vOXQK2Cz462alW6Fh+TPVp5Cqb1oQ6MR6wBAw
A+ZKd4kb/BBWcZSRfyRBgT//oVduNEU/BbsYI9SW3erCfaTwO5mzUZqIIauBQxAJYSp3F1pOcd7P
/TSfBPIivcnvbBq0U5wowQay40NOcLLVfLbgJSLnDQNCC0g67xx3VvjCMXwDb779Rq5jcco2oZQC
hwsWUv6rRG8QGJtgdR4AqOAY2Vt1cf/1jBtIMduUjNLq3YbFP+S766wfORScXE4y6c3IdQ4hI6IX
wkR29YsKhZz6FO5mIYedrbVoyLk/8AyO0ukuNVAVgXeDZBzMG2fA2JQ4+vPQvp4g8uEFKZIDNmBL
XkDHnMu7vk/7E9V6reX23tONHUOSrvBVSdKSV7UHpsPeVTPfLMK4+MjMnpUz2o9ANrJ8Y/2pyZGz
l+O16RWFVPirbq4KoFGs8wnoUEdfwtqJ1FcTT5XHWGoalK5D2C30uBSf4Q1d8V6qBVgv2wMuOigk
f6QTl9qVvTeQun5fX2sh0lm8OuLrE2I3ePwMDZxddnybHLo60RozDvysGnzqvEW/Q7q/uWxJx91w
sUsufCNUe18dS5ZbVP67gv2d3UVOITNEbPxVhL3180M7+QZVOms5PpwYjPB70LrFn7y1cHMZQ7Dw
939WbbLsx33MfkW8R4mN+b7x8H/tygLQCPK5TuWxq8ZhPxMoizVWx6M5OLK1Aot/mckLslKCGd9a
K9nvTj232v4IVszgG+Jw1l0mWUr4O1Cefe8hEeQ/Bn5yV7kI8ABlvcCnj/CMc7+719JHu+JCAIZo
hgat5tOgz8EU4CYfgM4TCniayyp3pNO/0ocmdPB0wviWNEnkzgPtVAWvxA550Xs7dhf+THsBzPdz
rddI7XCLwbwFhtlkNij8hxQRy+hwnDFg++A+SR+anfsAHeEhDeLKFbEdKFushHljmYUzosDYRgEL
AX5FrRYALp2+SGeIWuFWu7d6klTtWQKo+HF6ofnRNfYxEiLfF4GbIxWitnx9mgJXcf7sCF2dUZOH
IrbYHCqdnW9ttPXYXG5YZQM6GRRzd5XHnmvblqAIfSP/C2xQHjEfxYCO/peQTshvA6dhPjocYCAn
2I8iakTPMpM8f46EPvWWrw8/6ytuiCyddNaygeuhlP1eUgjrbgOHf1cOOgB3LQ4u3xd4A08HFcsl
bM6rR1jo13biTyRcx5UWG/FHfQ9LUV9N9sD6V+KNiYiNG7+xLP+qaA8Lk6+UnwRbbkRsYXoJHfWj
3TbhYn8r8cMouSDHXJewcaL+oLzVadLNbzRPHOsegX/OaTjiwLk2CF6BURLK+i0rj3E6jrEmaZNQ
8Dh9pBVK8mh61Vy14PUnw3O4Afll67hy/vcdbnheNkmGdtzaEZGgP/18hwhvkvNqxB50q4b660gr
PVa8mSu8BDpmDbAVDeQ0pXdEiAOWcKHzE8ICi+G2sVq2W17mqo8UKSQfDiTHCNb54LNIucoC6CPt
VVwJ/H470H8ghoeiZg4XqQczxRaM8vTyo/kb+V341jC681TYAy14/XdRXMx3b115x3tbZn6ubLYI
ekYUeqNQ+gDFIUefZzLiSczlj5gfA34dPrnloRQRbDnOUNTGs0BX7LKFlznbZZ7CFAsw/EgJJIik
EnZre1zcbHNIr/3NZGoSuIOS5GMrjSdBJwoaV1I1BQ53Hw82bWUFVAxll5v31QCn1lb91tO3zfw6
tfV5cjWHXNzBmwDHlcgGoXtaXAIg+qCBp55He4RHhbVl+rUWrA6ykxzdAOiT6EQolPGpxeUXYz9L
ZS3lCvqV/q3W2nsB81TsaBxJ7Fijdxtw8Z97vKNOq0FFbpUOAA+yDdJuwAlXNUPYGQjtFhsc0AlI
+lDpaO5XzWpQlSCNlSNmtmEfMT1C0uvFUmW+wXXC1t1vEdPWW/dqHJA56pJRQNSlmGX5nLhwK2rh
vDXse4RXEjYq+fjBJCO5eVNO3fFeh+vPsoemEirzlbQWD5PMby1ZUi7dsmXi4SuOx85X3wZALua/
+A8T/IZO05ptK9ehmKvxw5/NfrJ9YItfMCl63aCRh3ULepndHk+jFf31ibtg7wW7bOzyfZsufhfZ
oVPuqYa19DYos0RnISji6YpA9JkXDJLL7Xe6XT4U7TqZqPLc1VkvGEjDVkCbd3m6XKIzFIpGroqC
JSjiffF1nWhj5cMtlTjY8D8tS+2ZOXCJXAygti0P6jPQb7dlTTnWYjMR2C4eXkBXQO+cjFGPkoeK
DhyFo6cjuVNMAxY2vk6F3gxyTwdRWc6KnrO5Pdd3TTw7WZF+uQboHjwSLg74x04/W8vWAlfDYkCz
LCMFE+GlIT8Dh4C3Xo80s7/yRFjjGZNBdD0eYw3vJoy4q45fKRXCZ1w9vFhjo/yFeGrtpqUB3G0i
K+EwknZnfA3QxoVBdQlegrd6vUYdb1OgRlgXDVzdFgzbYfRLPkS0J8/jHlSbNAqzPCzTygA1R71i
zWDffiTy3poCywR1/YWK5YRXJMkQs53oqf+D2lTKFAWjKD52SpOVs15p6RORrxZPBs4LI9NuJ+35
5QmBHWVa+cTUdr+f4cSTfXWLdImDyZbo+phhhHd/kEdSijD8e6Ny1RUpwVcQ81TfQlIW6UVltbuO
+V937HHrvW7vzIiEPS+GnzABjgLRdD6a1+vmoM5LY5uduf1id2WyZIj+pHt0N0txvHrDP47/2Mm6
heyR4O+iu10F/DPpTDRdfYMKq7EoizqoMQPlOFVtoBwPtKlCvbwaRK6R9N5KreJvRkmkp10Wp7RF
gxui3sUJNlBTF0SxTthsV8e/1t47WhC1awnaXFFKWPC/OkV+HyRjOp71FDFRbr+N1cmYNeG2Bqj0
9hWbC9nA8KJZX5VP8awjLdncVL2qbTINByJwJ2l/PT8yRL/zO1h5Q27aAye6Xq18QEhojPANnctI
3sZ18vQTtpilPom6GzUxG1alIUWWVvQJ23ICdgjYQ3NRAeJGed/BhrLDo0lsW358HAu0hlg0hOqj
2+5+Vvs6hXRk8NLcXpDllE2OruaSQn6ouY4dF2HOmoM9JyPLHC/QoJG8xZkbU7vJACpX15da66pS
MiEqdKRqz/LchevXwjJ+L12D8pBlWzFrmw0exW1ECUaS9GsquF+MKfqbbeHzjVHc+pYphcU36YPM
GTT5OhsdsFLHdOTFPA2XT61aEqsC7qSKdV0/HhYTakdPK2F5Ke9fKfE2R37jh5C9/0two0CeqY5e
RKr1RldqsdX+g9b/c0EjJT3z0m5lm/f2Zv2zc4FAjNQHq1jzXsZa9rf8VCrU96PqHabu847d2UoZ
MjqasVZwIAaYGVsykFPhCejbdbtmU3Ovwn20HSNnbQk404b+MPss0lzu2o5RP+6F+tt2Iy7Reb6Y
vz0Gh2COnt6AufcQYYiSJFa0oNza5flK98igRs+PBe/1alyZaeSL1ddjVmGwPCbj9SL5fXB4CARy
SlRwimieMJ8ik2sip68IXnwSPZU9qOPZYh0R84RK00zuGHJh5hFQRDzOJQ4ZJ034bWuqcjVyd5/K
cNrE9/zRF+l9sz43Pux6epQq0aaYhu2Ep7WmdklwKzo0YkKi4lPXiavZuWzircC5Ij7my+oXWnpJ
/sj0m3oz0j/iAFDraC+0XWY6qPgqRZz7TT2esuQ58Dz/KnnpzS9AIxeKXOTzwoOsUDV6ZkUhJaxz
gCgf2FXXvCNa0zEi6y8RUuEpqJse5uPyntOI9lVLLdFKDEqJjTjYSGJ/scfVU1rcgBoX39vi5APW
zZ4N4eEWqUhYlF1yqK8rLE5hFld0wQ33aEk1ffgrI4ZUjAAp2PlRop0txp9FPYZgPYswRESBEb1B
KJR6n4IWqADZAze2oiQ2elEu5d59nLxIasrarSCUta0/1xOKupoPnD1EsNLNuizoAspZL4aYX0po
GI1pSTWSU68fPVPnesi8e91Npg1dO0J0VzfRUU5y7YF8panSclEWzz8Qcd9cLHPb8/fKlYzRAHzW
MQvCJFcCtgMRHhkj1XBYSZci7hJTHzvTEIHZpaEJB4vtqpDWrpqwek1CxVkJtnD6g2ueGYcUPQ1x
wJDPOG9HgTy4lUnnodonucY7JktNbdtpVgNzQhHk13S6Wej2OzQ/mdvJLcasaM5NXrcqKabOu1lH
bH0qWdR5dJ78a5D4eeGndSvTyDVUvK9b3v+lti/MUfvgGPOZD/xE26rVSeZHyTusd2y4rmO0AO7E
JJnkfT0cA4szykPYFEDL0vJvOv/jHxnnW/7e+HHhbOK49QD4qcG/eafFw6sSdXP7uhXk+SoNIpyJ
9SgG2H2ANTjmpUkB2JOasSaHXgScd27wpkdnQ0Nt9IifcQ5LD5g8Rfnn3+9tOaMIPB++ZD+PgYD5
Hxx0GFpW7SBxk7tV/PRvMqypMF4vs79GDOq4QVmb8lqoqfW7A6QYhWB5c3n/ZFkThZ0JRihKlr2x
GsaNcoi7y08+Xk/2fGIdjom8Dmk1d50B9KJF7vreJaa9o0F1PtclMe7cJeKx6d8YM3ynPneYzjyW
hyY7YlwSJVdG53lCh8zkdT9k6cMwdicxG7HqSQAZHIvkomx0+0Msxt3hyd0+AVYJwHLSt9RjAAaY
jim842nUhTc50TJev5qfVMy7uapVjloy6zYnLjV2lOb3QN1PEA+TvVV8cJUC3llSVMdFrbig/xP3
eGyqyshrbZNyugtH1hmJKk98HnzLvHIavfgUg3pJqxNc2JS85ny0NRBHzY5+IvfybswuTaYs++TU
hiRW2QY85hMKacURPH3JSsBDELA9Qum1cu9mjDXWfaSJtVk013YdAQhhq/0IhspMIc+yCnWZ33y9
2zys8AAYVsPKTdlAUuLsnLo8Aa3hwWCp8lTFXujK2EMkZV0hjEDOJe9hF/ZIWeV8nEiU3VF/MBlV
7jN4IaUe0ZerJ/gWTIWG+cIhCTUmNjeyPBYWjQwO56ipg6Vp+1egT8q3JQltacf4I7O9E8LcY9eX
0LIOBGTH60omOGy9XGliMtYHbFhJC1NOOw6hWYSrs6vQ2cq/sKOmJpHZgVHCPO5uZ3mdCN0GIJwJ
VeyCxziJzWiJwDwG3Pd2bwqKmdbWJKPBQMdSHnrQAMvKzmzJoplluNBelzRrvwmlcJ+SEzb2l+ix
2JGMIEDIhRL//Tl1jNthsvJfFFZHJy0UNrTpwETgvzOMJTvWdtvXasxLHiS3TjR191JjfKp27Zc6
CDZJKaNhnx5gNLmG9mstCpam5OsBgakpx33tuCmroxV2VO57lL+k0al+yb76+Do4T04J2FBS531N
FpPbs4/tItETar1+TeqgS6iutjpcTnAPhZtvnXuPE+58t9MxT5rB0+sCTxn0PBrSPWjY12Jh6Hng
ShGD8blQnCQZkEx/Wxln4Wqrnax8KKn7hdWB4uoYluRsMp+R/zaCTaf2tbyGO36cWUBpq1IDdyop
cCjzPm7ipONGcAwsTa9KvFPwQ2j++uuG6xaRtnNKLX0ihkmF++zclLXkBC+ruNB1Xx0zwnxAWmKq
sNHUNZqg3tmMGjTt99t3AF9aVCFWq3G188DlyIoXOu7NucF0mdfZuUgc6Wol2U+CIroQmJitu9aQ
+mOLGb7JmGhbY2TKfkmJWylSMdioO/Y5Rfav1Dpf5YGwybFXE2Yt8K9RdGBT3DaSkqcIpHsxAeV0
TnhrgLuLdGQTQ1xBN74hK8YSMJP3nWyyJRXXFaaLz9pvO0arp6fN2avAZHl2Efws+FSuaWGPKEKQ
KjKtBjIyjW1IB+KYNzwUKHM4FBM4GA/vjP87KjnWlZzM2HGnai/gUHeQu2x/cNV24Ebvor7MwO4W
b8ABLOSRdXaTaG+WwwfMe0ftvG0MCDhh3K0IzmZBioLY0dM1opIhzCBbrTNJPCUH5JiMxQajQ/0Q
5DvFVBAiM/feBrkBahygmg7REcqrZPNgHCIc5sUqZTBmfVEbI0dTvPmyrGFYT+NUT+LXeynLBWvK
/OZ6CKc3On+oaxVrZlmHPOcrSRNMnq7s0vfAC5yovynTOqv2jCBE85bMNkxDDlo97QMWF6u+kuzC
pa6Z2TJ78RKEHX5jUpr3h2ZLFedNElD48mHPdIPkd0Asl7u/zDq/FgUAPaE9AQR2qgMlFYDJFMXs
WKUWRkKJTYuxWCF1KtLiAY7iI6WcmieAiNJGNUY9zVwvOWskN2Qq+tNZ8eLJby5kztH3dJHcHtll
4fpFylZJj5RdYIdhTxONAIIq19zsJ1+CFXZkzTyf2hWh3rhmRF6nhIpKruYDT4eE2NzpnC1sQR4I
HZQUme0ZCvQDCH8LgYQA8bBfJp2RMdWw9m/oQTeKl027/NRDPErkef9VYmeaOWYYfPo8WILVgDOd
kw8NJyqAu9bftKjfzFqa7hFLrWGvo+psZkDLhnFL/ssndD5d103w8VQFDi4J5smpgBkCp3HZEdFS
9vA8FbYBYek9H2AVpZPHVEMj3n6MBtCcrSGapXAF7dtssYX5mDZplb44IQqjTZFneHDl2g7gxGpk
BV0Kx4o2xjAGElKbg5l1ZqqbGiPljKTHrHDN1ohMzpdFWrbfqrXqWun/vxWr/1H6BYJbBEMCkg98
9iEX8kioQ8rDJacYnjuc11YyzDFQSWKyxYk6WSWg5gJp7geITTw6eSer3jDmWfmPit2rE8+MO+WA
xiyPNWPf7T/fvAK0w/XOi5SQElQNXFDBgrxSZTz5H2ZQiMNcQ3nWR0B76rgW7R42ZPP/M7lA2iKL
FS6Wh+xBBLJb0JrKYcc6OGwd6tkbwNDZ9uOiBt4c+S9fkTTO6oVDu9SIQjwOycfN7OFQbiL11iyz
YpCQRoyB6felDorkMGyE/vUenNZEQnCVHZGDVaIcw/D5vgmVgfgjvBNFgIDYPOjTjiT5VvRodgVo
4ngZjvRi3Qha+F7HDQuscnMoA6pNNpjJYF/X7H9PWCx2aCLo5ZxhsEHzF7hjs8d0Lx0G52w9zkPG
Y04IyUUtfp1YeinNMIUxM02Cs1W89h2KCP9VpUKoDehzBb2JjHiw+NzqJzdWpJPNRfi/Ccpfxu+3
4JXXXq1Sr75bgSiIMGyHuYVvehNimjgq7iulFi9luvHFpXK89hamx8xLPyMhWGR52T6bxOkfS85Z
iXHBQ++xVNZ0W3e832PFLzWzAzNoEdXvt+ijCUYNKeh21RgQ481qMsMPzA8cC0az3p1fs4hD9aM0
yly8r+dYqv/t99HTRdV0nc6w3epqqgr+0SufEaTDsN/iVm4hibzBPGGbUOzAzhOYG5T/aG5X97dY
Owoav25XyMHvR7ago+HxkLECYFWPUiTPX7MJSc59acdK7URhiDb18B6cdBjWcsMlb/cSH2zYKJEB
dQxrkAPvPoFv1EPcHkAlNL6m9Hdv2dMVt3AFkXth5qPHiGip8b9J+zyQb0vlbN+ecUtKjHhar+NX
7dEWg0yowcuownhPlIEdL6ZdnoONuuguEvTMKIbBxDqrGQlgTSPYuZ7r+lguoWAhLUX4RKXLA/bo
l/rLMGwcc1QPKc+QgSCxHegsbqJKXECRZR+QkxxST/26vhNV3QOQlidmsb5ptRSMtYDaJoOiEkcw
Q+pzFBhvz+2p8CP/oAIUC/9+P0GqovY9wRa3I7CEcu2NjjC5ccJiVe2dsw1JRK+MyvCFFdS5baTH
+C4fu3N/i2Ace3F5hBtVEzKnq34ALHeCXIzuWyZl2OFDokmYFwnAOk8ha9JD/Aifnj9IhoMSp90U
MjxydMiJjU4RmUg1rJjFILkdgZMPbM0M96qAs+VDqTgouFBIH0tJIrTgiSZRIqR5OXQOZQrzJWtl
/ytUiP6FVJM9ACnR8l3EKU2Edu8UPpiCUJefyPP/M/qo5QcsGLHa9SE8xEgRo9N9KlPPnXRcuYcG
uoIvOgdYnu5cejlrWUpb3zfMT8hBVTxIPyLXhGrkanqHIBO1nFc4ZAYOXf5w7UaWhSTyHIWUM3l/
MGdbjz935wvwQgGX2PSILZN5xnHcP9XuM1JnkxYC1ggjJLOBkux4AZhjXcTHhG1Qmm2UitHkXeVb
DrAvBWtud5Lw0I24n4OktaWlTEX7AoXjD5oguG9WgTiV3esu4/IzP+nL1uErrMP1e3BEdDDa4lL6
0Vxgjlo3aKUG6fsD8qeF0SlOGSldU3jEdi5d1RgjbIrbOJqOtaCxNIOTUOx0berK+rXL7m7JmLjb
SgM0qj8hJUaYpZXMUQoKPRi8dYBitLQ2x9LsMemptgwA2HZuoEH52hPlinDmgXdc11ZuSwHbeWCJ
/XpFC0YfQe155oP88vmaB5VgKPmfKIEr6+eFhX+l0Z221EA9DlGCuLmib7PEMYvif23d4mtbwgdB
c/g573u4VlaaP8YwDufbqRlzvAr77Rplxp8CUYGqtVdJhxOh9dg08UU888vIPJ9FqF7PCIWnkAug
I3ARMya0+q6AC2O3VkgHS3bxEgRkmZv9/zvRSO+cGpMzRoZBUfgCwJW6RCwLWAVIue7/Q0NI/SFp
J2u3sTGHtBakVGsoFrR7Jyzs84fp1MqdSCNim7vuUiQQEB14Hw9hXorFVfaeAFRJS1MTtFRLKLfK
4OY9PzoA0LHj+uvN02wOBqv3oq3O3Ky2ML8xn4ujdt3jaD8kSNRv8LPjle1jbrKxvKab3wEk7qGR
fgzZ/Hs0g28a3bB4NMhEXhjgw4VDsmV+LBD9uJ2YqgdG+aTGYH9ydR6ccjamQtk3anFOdS+8IMk8
gMeqxePhwj03nHB9Unf1zBtqY8ONRKk44J6fn4XBThPxrR+dOO7/RDcS78USgFeEwQR2iFtiAEHL
12aDcNuDAsk811tan/NPhpdGJsoCUPEsHPO1VT9mzAqjUNweOA7V9RDWy+e/mVPKNaDuOgGxRLLQ
6RnTrKTQRzoz6rgE6aimLtVqzAjqUz8ohA2e5pS/10zk3XKir7vHME5VdYMVwYhakpj2lK4uoMSd
b4jhKDBFLxodXmjKoFEM8eNbtbheVlN700CAsJ5SXJknwRfssu2iSY2bnhuBC7/ZhzCMzld3WfSl
fGLhluoTx7Bs0VWktusg8TVT+Sc5m7iiBc+L+AtSEZCWMWWPL2SKGLiE3WHUyBslIUTRmn5Ae02b
uYTj8JFuf0GW/lX6x5vK2Z6+8jlxGP3osHNdz5WvcXWGzSR27cWftxrctxEai0Xfsod9Y1+L9F/Q
NwjfzSC0nrk7eJynpzxwLbeGMm9nQNbTbEH0nW52hgHHQIXxcV6BiaUGiw87mM2OG09dPifka8UO
VBjo+2lfynlkhnOqNqcnUyhds4m5dgWsiRV64NhDJvHjcSbe44ICLdSPkX1kWK1574KPtgr5ICCS
vR3npOLUIF3nAp+F8HOOSLYk0sU1EOCZ9JVPvISBZKNwLmvJMTtGTsV9k0mqhSTsJmzJxUZuP0Dh
W+aaDtktmOZestAtsMqgKpzS1NQ+qvW/AuJG64030f8cFK5ym6C51hFXkV0785vd5QsjfYR1iYT4
EXK5E4NFlRlGGYPDIH12s4If7/7Jw90DuTAIhqx8AWtTr+E2mUb5gDW2zFCH8/GB5hfmWqIRFcUu
Q7hwydVyQws+XAljFmJgNXgSGTts+8kiHAI5XIIw/f68g1w1GGWsnmazhi1OfOYQsC00WWhpoYFl
Ns/1eg8EPNyG3oLiaTBfBOIAppZgKI5lcDgNGl1Ytrdc92ZLNz9olYI4iK9HOFLNd6oxX7rW1o33
ghMc94BNuJHFC1P4eprEVfOKzpY5qkVC5ycz+JVIWwpgMqYpzQ53fu08Xrx/7hTkrwQnWGkjeAC8
Uq65FlbZrHbmwV1j5HyQTCtnQRQan2VTaN6nGdCuG+mSDTS/SXOG5Byb9c/FmlcyPutMXDowI3i9
MtqFrYQRgVvKn/ZW9zjSwFog+OS4J+kz4negCF1v3RDZIje5VGprJh22CEeXQ0gMG+y9INBU+Orb
KGCoOiJU06dz/Kq1uzDvAfq88SxrgJeOMKK23A4ubKaJw/x0jRDMYxPX5+pXRyZdHJWEhiKQC7y/
AXHUUV9ZMU8wGbC20ykGTOKysIsT/3xvtCwP6r6vfhCyxoAL8VS5MyfaNJ8/ll2vOu0BkxsleSUR
jzhG7WpYrYCxkC3kuoENSpRTUNnrxAn0ETlskxo/GsThkEuAbVgstxd8su4E2AdQrM1mgSdHTbnX
83saB0UrsQB/YAFUvlqWD/2AIjbHy5P8bc99lYSPormR4VjzTrU42Kp5HsFoAE+L4jlsJEt/76ia
CG0Ivmmyvx/31AJgzIiG+Yc/G9fM6hqRSPXyafvk0FfGWITLjtxIZOaw2xNviIYmDRkkpKrl2huR
NJ4pOZtRg6pyCxeMBohM5pIE24B4CPuVXEz8rppzPM8zzXMM1HETOJNOM5DspRJwvUeAEMkBztIB
ix3bNL7qLtE8TWpe4LQfbBvNZMVNDiI5JsQkrrcJhTbSB4vMOrCcEdVHvM2ioVLgJ/QL+BcYw33v
k2ASvtjWOGc59R14M0T3pVDnTMz9ZNwYTz6ueaU/qHo65DBHwg1kxtkbYI0r3iWZuGLh6mfRlCwL
RNQbmKxDK5wwOKpfH+Xm0BV7/DYdCty4/HyTwZ58gtzQNOB8ajKKVA6N/IbNFOnidaikVh+UPlqH
98Jnd5Xe6EyezC4+1pp6/PZcLAK4jCS1LgvN1LrkU3GTFKa3rnpD97MrWmBRVg3fYP1uihayzLJO
0xVbrTypbUdgzDn7HIp/jFcd463GZOVMqOBwUCd55RVYqvDz4IQpjzb3qDA4GnooCrcY6Nyy0yb0
pz4SC0hnxy+5wniMdqfimXiCbN4qYJQrn3t7m2zVxWbBodADY+CS+r6HpBaXPXahtBTzL9QEPDMG
vXyTl3/zTR9xYpHxO7XpNeBEXXJUO0y6VBF14xuAXmzLK9R9mMP6hS8PpsV4b9gW8hafwGCcV+wI
Wizoq9tic1xVVxCsbCl9qnWMZhzaSV+zWX1sNeUOZVYGlSsGDSPxwAyLgVeI47MIGpde0u1IabJS
fpmvbYVLgrzctgX0qMXfMh2V7jdq9WfoHFWey6DvZjLl4KLC/INl+DZKm0WUqmEWEyhfecMledjt
IcbEz7tGWI7Ds1kfsJ3S1HmwJu77JJMoSlVeWF7Picp7FbFXAQXX5YPqo0tzYcisA0zveiJcxayb
CXrNst9wyVPvt7AWw2xoo3b+6CUjmzcVJ7u8hJu2zl6ojtSq63H1nx/XNL2JTSbwgBJnwCZkvBPH
UXLzXid1SPmEYXJhLaPPa2LVW8jU3D+ddkrLjdNmZDeGf42uCRRlUnNdfzvTNI9QtsF3evB7CV18
HhgOFyOYw4RVHhY+6F3SbbBH9OsX9HllxKMuf0YaP3919XEzGmXD4QuzjnWjI5dH5JCCWECyA/Fb
OVtTaYbXbb5E2ocPAL7MMnoMz6AXOzE9AAOZfqXEgcT0+CUdjwD7hNc4/auO/+QVHWDhyYnHlYE7
Whvw0fpQ3vgDOQ+wQQDikTrawpToyWVB1Ie254i0fkHs63e0Srwty+GmnxhOTiZ4s06tiLvMFApc
7JSVwzyGbtMqAWfCQe9FZbh2204cHTfRh2Qvum9WA9XoxH2ZnT9IfpCOYgyp7aY2A2eKztL7bNwE
cBjF7duTzlXFdKIViI+azRTF4k16tpxMPnDA+clx4N82OzUkitN8WjzU4i9tmjiomQ2VSJ59JcAw
/FyYznciDyucvS/+3RHpPj6Cc/M7K3CD1+ZSwW6fzzy6zm3/Y3FIXKfCpE2tSwC93oDXKCk2ZNG5
LzzocraD25KG5RpWrIk7HaVwsIPlSlRnqb+Y1CYr7hIcrE45LpkOrUNA82O9Hc011umwYphG7kaS
wlFUviFqsF1mqATeo4BTBEMGr1hrP7yWm1dPskxys1r3HRvY0EtmF0YkmPasCwVXbilPzbBuDR/E
kOy1iJiy2t9Py/2sR4+/9rbkJekeP0FyqxJmN0QaH3yJWhmW4yZb9FDFyNvxRKOE3wZjFMBgTMYn
/lv6UgCWjSSagd8H7JLEWk9ZsrQr6bsRAu9BdoTFihsYusUooviiSWfGaewzN+u0kXp/+jGX7VOa
Ub5JnMEOQrSNn59uLWm3kIxqczkPCF4KiHf+jUAjLQ5XAuSu58gFArT+CEBAFF3dD+XHAVtOt3pk
+0sFgAgvZGbRGj+jtVQdR2bt2ceb7r+tCs7t7Va46TakGP5U8jeaztmQB1zmaHMM0qOognSqw8WL
wqtc/xOVhkBigM+7N98XyyCByjJgaJ3a4jksUDsWGOMrrbzVPp2ka3gJi1FomAirxgylbdgpW8q+
nsbHdLCl7s7kIkkkqYxTKQfSvtVI5jbo11CigzGLfIbAHIzEOctzHH+TdfFaOYsA1ecLCJ1be76F
ul7T3bV5HnUur+HJ9fTr2FcnobthjtCiXf5p5BYP3SqVBxdhR65IfskmhNvR3Neb4d7Fla3XJreE
a1NMlt0YzXjxgOueaktfisDZGR4vLBBCpFWaCDEQWxlX1QyCwXlAJaYBjEyG50TTbxaobHUj2AjF
PmDOI9Rpg021UQ6Y7DAmLuQP9xFoGM9EcPXTffn6Q2PSi7o0V7g+5M7Lu6eo08buVxL7HYhKOtg4
wCOO8ubKF1LUI2KHe4ylTX5IcArdOdSgK6XNfeh0Ngm62p+tEX/IfDCyfyqmnsWz8vftefBd1UH4
QYDca6VfctWGNmN97xbHdkPpMckSlPcpbj/W4795APdqz04kyDQeeSa1vQY/5jXx3ywm/arACWnZ
TqErNxmYztALsRzfbsn7Llp+dPV85urjhmb5wHfgSdumF6PMtFiZgJgDl0zlLLv6j5RjkGnFqqGI
yzEljEJMJJEVtOirxcxOOquIOD7jH7cFrRRq+T/VO+ErFZ9mrRTejSA4gD5FEAynyttY06TYaatg
my/PD6TS+kJ8ViREEKfZiPL5sbZMwzDJIxQxs7tqayNhZ8N4tBrp73Cl3O28cVEsu1spvSF9/b65
HMd9EnDshKnBpkPwMhzOqj9a2lVq+77j4vTfI0977dGspvufBc9iyQFLEjfisQ4niyLHlXHr+UeK
EUHkBKmlT3rl5Ef5Jk3s/RXAe4UNmGDzP8y67VFeHwrjT/xD1TLr0qxqIA0/YxTAbMn/J+/9pAxl
/hBIhhQJqMsVmgXz78h8SHh7Q8zv3LdY5kYxlSC5ZrUsNOMdwsJeoncil/O0QVYXtnFkIsAZoaXd
7FSoSUwqSq+npgJG7Q7+SxIau1hjvNyJAc1zOVcMWcGcnhFNWs4qgu3GTeov5w3l/rmDS5fwPwJl
GdJT22dXL2oAlsZ3UmL5cBRaMIu/Ia1XhhcEHpAs5WdPnCfVZzQ/dKbKM+kPSAxE4N+atIaZia95
3c7YBCMTXD9bL41y+YnmRM1nVB1KE4kCWaN5QZljYAfkUuq6+C2FssJ5VkGJSim6FO4y0RXVZRTM
q9PXkoOK8wHYkclmY5wMBYO9WSL+Ziq0WeZ8ejCUPFC3D4IBNkPuc/IFPGguHQH4M+miGuX+gKnL
Yk8icSI25li1Iqb63uyP0XUTFj4CWXgIu/WkmV/x6+KyBjz6WKICRTQOSAEHo7j/gELT0WS7QlFb
D+k+mtY9+z6K35a3gBZVyXRIs6u0T2zG0xsvIx3HPf+uH2zmBxEzQ7mk9zwOgIUfiXBhZXn5Q9g0
3fA8zFzw27pieYHqDv9s/JzFCA5hD0zc1MAeFzhjf9a2cOJKQj0ayiv9IetjIxi2ZLQldpcVK29D
UTpMrr4G4ns3P46Lx4B5JAZqgjZp/8fsQOOnT9BfgMI7DgtX3mZYsHUFyI7//gLBqp05/zpd83Gw
qsuv5ZYRNSprOxn1knI3/gEvUcFrtDpzwnxzEVqsERZy3QvhEMppkogY7bNM+5bm+6LZuvRpIi+9
Sza3KohSmumtcbbG6uDEMrkBTa8Z4ZmV14juTkWVJX/JPshuVnaieGDz9A4//JDpIuyjd3pHXvmE
NlI1j1nSeE+ZMZsZSpL1Qg97XqBQanwczqpQOvb7h9n8ru0hr+tiIcL5RkI7DmRBUpRr4opB23Pb
Wt/Wer6gngK1RNDNwUjVY3uZF/0JgipxKethWNmTyS2k5XaMTUZZzWQMZA2C5oksYpZK8xk0khrq
r7i7SeHZO7mbPNN16MH+zBsJFjbmvbK6nWugho6qwEeWHmC8OOTf5MI+BRBEhVs0yhEaMrcnw5m/
J+/jaljOubki/UUnfLMhXL5LVoVLYb3oAn+uthG0pwkHLM3TNoGdp6CKdgWAsntT0jRiQa9kGbsI
KaPadlNalYfqoVfQ/Ra1BkdnRnaTzrrgmed33AEICHRFSJ6WWJVebEFaOwc9QMEmDZW/xEPybFKe
VmuKJqFExjseNkilnrIKF7SZHl33vmZpwa0LO4aTFviiR6dfayWhBwXlDF866wDxmpPum2dOoYJ7
pLfKluMRLJs4xCpP9mLDD+54onSp+ePmpx6TQcciYPcYmKSdC0utonEMpKw/kGI/EK+FZRWA0aF5
Oa3osnvg5iCRgzWJrHgeR3lQQIFETtvRox1tiK2TMXviY/ZLPNJ4p7YazC0uU9svTRGc6HxNLXfj
Pg3POMTNeNC4hh0zFmpur5NlTjvWI6qXJ0cIB7dH/yh29ldantVXMwwEFUaJ88mXzZ42Dk5O8rHa
uZPlo8fEN5B14sUZ8IRrE4yPN0s5/y9rA1Lhpq8iXH8Ohk5MhuF6mfMnDR+LR52eaJ+DRyLw18o+
28Gv8tBbZhpASMha/3LvHI3X+FOBnpmdVUTXCJlQ0kdFWBBe87SLpXqo2UBUllPdfp+WGXxKUCxi
i3K+YX2hv6JoJOjjrBwlgu8lDgxu0YeNRdRk40PEVKdK61I1QBaNip0LLzj5laY+rH9Wriw+nTed
cbVRk/a8zz1BXp47ihK099dSJwpbHEt2R3TTlYMAVKkLq9IUo45gLhJi7sey1LTgpwIW83z0G0eS
cqQLAkHSYoY+IWj9bxDMYwBzZR8JYCYxs7rtDe6Ixdbw9ifj4LD/LUSd4+jiX4rBdIwkMOBLKmH3
m5Ebzg5ihK2dYc8CD3gG88HxsA/QDrBrjQt5UtVsZLFdjGNremUU9+VMH68zqkoESrvc2utxF6iy
hMtnKs0MhrfLF/kri7QDuUhHyyHLQ7jf4J6+ipkYXU52aSjaGXf/JOntBmxYtc7aa99NZmqKnqGT
bLFtyjgsG8b/MfX8Eq9+2VxohdNSRlcxdEGZgcGoknZ0SRP793sg64dDBMJ4LbnLauRBn4ygKSJl
tdP0ym0cVyh2B9g5XLKUtLDLzJdnuQBVLHNElvzzJyMTjpZYxruTG5O2jEWjUDyEbTnC+sJ+ZSiO
aqR4PO1SnCBDcAlQ3r+5et/pPK3gfqZKnIt8Lg1JhNQ5Bk3RBRxX4LgFokW4msZEn+c8IYQ9tbeB
+VDSzhg73niPOP1NUpecvajEsA57DY49wQmmdpPz/A/X83+MsbUDNUubbNvztg66Zov8Pty+s/VQ
OjFBOsFKORbheHAkuUJtx7w9xfHlLh1rqDDnihZJeXoWgttlGkcxb6kjLgelr956McFL9i3vLPrQ
8VTmp+kxUd4Rp1jR9JV5SZbwcPF3gHG3oZ2RmxR9b7SRdfH0NM7FaT9OFnoNYasa2+UaOJcMRdqD
swD99y2U5/sZWDS4+E/bv41sEF7z/VZiueppg22l5Kxy969AioXAgio8EO2KkBez2iNLBuGYnJSc
+ka0+XLT9yfUAGcfjnETYSc98IkM5+DHv/QHyLtM+6LwPkUwxt7igBSbvyWiRxX59BQXDXZDvyif
lEASJZAEEs39+ccjDQdqD7XVrDRvUdHHW/iIs/rWmKaoZNXc6bUTU4EiiLemrlXrC4WuwTEXaAlQ
XAc2NPtNq4vFU1Uao9xHR6otQdxLqmbSZ64NujV8d66nT+hBFcapV2nvgfLdsATAGXosfum2pj8v
+u+VES/3Qm+ezr0ZeqWVHjZV3QKGcuVSIm5GL0B4IDh0vCvwc1trjb+jGyV2LShq+WetuQRvfUDB
mrlxTqC4aKcS8gF9ELjIrDphYJeTfvxiUWSebAJMDreuzYByPrvmzfYt+q15MsqxDmq/Cw/6xg8P
PCtkOeaTSyqVk4sGzS7QmFp8bYg81VTIQoFa6vfkP/vO/06CRyAl/DGTzvTeSWtMDvfyMXzLaFpM
kT86ksmBuikEgEt8NUPYnCOvZnQ88CkkrbtbUcQP5PbS9rjV6hmxQ+xa/a/akcATMt8OZqpNbp5r
FTVL/cfaGaRIFGx2RMvFfo4Itl1yye9src7SRQU0RaH8d7PBPLyA6/KUUB514h4JI3a3GhUG0Wxj
1oLenBaJ2uEv89rmPzcDliEiE5Zv7Nn/lBe6n7VOMZPDDGvntagxgQkSKSz3bRtZ1bWBqPrmj+FO
LDAnJboiC/d32FNHXaUIwiaKJFC2qp0fH49Gz4SiJ8wrsR5Yg7DCU5XYPOkwtwYEK36UNQunzIaF
2/aDCuTBesMOCYXYSp1VmNLYcwNTyvvXs4/qHltIJ0U19B/ykHD1tJlJ19STQmnpWKZyLrenYKlJ
vxwXEdwOFjM9Epsp5zmIDdq3ldUlFmhxWU4xoGnCd6rcIYM8yvhXNN74Mib9RF7qtAbj5R84mAMc
LevbRcavopDPmx+YYj7gS4bHeDM1L6w1XbfBsGV5HoAjYGE038/QB+dVyNdBkXkOI2e67hwBYem6
P1ARCLkj44vlE2H8nN81MLpXbr4Js0U3w+lG/KGQoAQgLObC0NWpm/8ubv6ytIPLQFTMTc1zlIU+
1gIsDdP19PUTRU/nnxQqRaP91UBEe3rem1HLLq8EkQVBdsj1L2Kz/qaDX3P2aaQ609RYQ++lyGnt
qGTeU5gY/zsr0lGnunVzslU4bZ3SHpc32KvzGJtrls7LJfSeiWuFduX4JYDcJK+kAYbqyUlFeY08
429f+4t3fgJpCETHrvSNK+y9HO6+fkHR2GgijJL1oXfdA0tWHerpHISmxN9umHMQfbfR1maYd9Rk
SY1CHysmLZBGz0VQT9vcOQwQq3OKgBr3M1M5NhtC1McFpT3dSFzaaGiWE+0DyBKoFLFjcftKc3pc
LhQOAUEbVf9wqteCB7p5rN2C8PkTGaDo/tYvmPivTSGtwsMGeue6moRCKKOcux3yW+SK5O0ZXNSN
wYleyQrbBZAZstdimhH0Bk+NMK265uoBymMDqUw07paUtjfWH9poXXZgQGJSeK7KQo3+VpgtLZQ8
xdnbRvqyx8IFOCaz6gen09h+MbuWw+CBsmR8VEZrsMBCawjxXOiHVXbSVBQBAqBDNfOEbIo7+vy/
gD8m1pxfBxOFvIPIC98kLKIrYxtYXZskxglyf2YL4cIigMLXVieRLaBhQHQiD59OQL+v+MBIOTi4
U0povfHVqEXPVWlhkI7VhLv7qOn2JgHVxlHmVsL5Gn4fjQnV0flxYiluTqOYE+M6ZDuJWJ2iUl4V
YW3caCfhhIlzSa2/HkSnF4aw/qZ9vANmC7hXa7EKhSdhbgKD25aNyboK6qhm5L4m6pxtNKWPjMPC
JPK5QegEI+MMI5sSNH7PSr6LstPVK5p8j5aArq80pkYWcQOSq4Hd2ftCS6lF9+8YveoA2GnAjdtI
2GMJd4BodQgqAqaf8hckTDoHIH57hw5/rwnjSVI3L397dWw5dvi1fT0BKjkMzoqQJe6QX4hMQFcW
QCBd6pcNMRAcYAoImq9obg+3GLz0GmO4xuRqeOFZYWbvQte6hy/Xji7aGRrd0yQufJMZrhnzNicW
fZGD34p0iWxhlp30fl4Rk9nWg4AxSCeCPzpahgKpRVSMqWpIA3sDZn/Z4JRIc43r3LKE0WykY0zq
/oVdz8qmSLpbPvPhlWp2R3p6kmjWB7aqHdamS17jMvqeMk9we9aFJngFjX6qGWM3BYtgUWy0FBkp
wlYkpsEkCUeogPCqVsdJujPr3xKpLt1rnc3nxmkupGkuRVNLoRAqeUsVZmANrKqUt3kRksUNOms5
8x8uu+Gd7HbpfMiQWyI82kvjxdNp3rief6+DpIhlHj1DyGUXn3Vjdt6/dykIE4AcUU+9H/OZLPAb
NcSMHm8i6oVoP9A3fs05yseJ2Ac/uigiLexwuvkPI3rGyfG0/ECFaksgeC9Q0u4nBASGaYYiaIKN
ajT3CBbFaiDBVZ2je9QW6ShGB4X1HaEB1IhM9c3WLYRxR/8zC/uZmzFLTJbgr+g3D3Se9cmERRHg
MTDqHMsjAmDlPl+i17sgDnlQYRu/twVRFdXolA3g3GxMb9G7d/H/4Is2gMREouceRP8fA1gTaXyh
udyPrajVAAdGURNzXvvqS9bAqSMhj25DuIUsvM7CFKz8k1a+3nZ+G9MoPmqLNRuxCMqb33moo1fA
JboL7InIjSTlUlgiEXhiwLcqQjMwmjQmagxbEJJFNDZO2E/LVzInX7d+yuqA+w5qsCVrp/3+HJay
maxb1yDFCh3oapfMBrJbifDDKOTiTv3bNYd7RsO5TU+bMaMQr0Wfpc7WlUaGGLiKEWpBup/XG44l
MmyDGBmWS+M3wJnD7vSHvWSESjby9tg7t4AusCjic/c2DcqwSa7CAwT6f187vMO09e7mIUGEczSe
/K4641v5fzbfs7sLyXhNzFMsUbl8nc+gOl3UEo636PfpBUzZoI8Qss/qUlcIKu/ibhou2appo/qJ
gP1RuaBp8agV0VNWvEbkIDWMLxtd2YNu9iAlZb0cvDyp/divYd2/tw18eWsfc1Hi270tplmDFfyg
PSWDSXAWHNl4oZ4Klu1Pgj0P7KkQBDVneqGo2jPQp4NRKVoLVdvmB1euCKhGMf0CQ0vOOlOgrU03
ZwTuOeGVLGJhja7pl1p75kcLusIDpAXKltS+zEbU9S0QGYO2hXSDyReJzdFmEihaZ7nzWjfo59wk
6PNd8mWzz7Ts4ThPMOX4TlTNXtuyJilC1HMhTcHxJ6t+OvY9zswBMGOABrQRmPnt62iqHKBywccP
yBxPydp5VB++Lgx1wSaJyqB20TYzxpO+RVtMKIwaMt66w0hx/0xHtJ+m6cAjYgz+pvkgHB/h5IdY
CZazsVeB6vrf6wmyT7dc4goLgmB+db41hX9HlDImN7d1aXbwqryqisupDYSUNDmAoVKhkCBW9rry
aU3cbna1d+mdMMyTRHsEP23BRfJklQ69lM5wRohKv0kPvWxoAqCWLKgL59VS5Jxftcki7QkOKCnV
zo4RlkeWpAIxq9oVImORfbpIwRO/pEw7OE8iVGDkv4AQr4OFuoMZFpoynNipvKoV7HOoyTzTFYMg
X16zMUf6ojQ4rDAEWNvvaW7P7uoj9QPlyIZOyRYAmFjXkv6KZqMRdbc9Eu158399OhUAtm1AZVGq
7+gfmPQPxTBv8VcgwH53DF/BDCAmKQikl04SYV0Nf86a6VCLSYXIIVESWey7EloWqJNx/W5ybFBR
QF9K/D8JuyhuWAjXQXB0JYxy38unZR+adExNFbxzW9Qmv9mZR+xpr+UkCeU6MPcpehkVp91On6uG
8ZCJcx5uZpsn1Wd+cEE7H/Ofk7lhxN8WmwjwEZnLALaJT1hH1PeptPpcQnX7biK+2vO36EuGSGi8
3LuqRex15OwAapfGDja8uu706OzmHEE34wyOGTACxkIwwCoC0kanQYkoUuJmvaQo6NGBk9LMzRYk
53SWV5kl/nF1wh3OvuQsdpISvSnAETm4bVTD3cxW8bEoqO8wQqLBj+zNSkdGRzOjX0/GXVUUcRE3
O83kdLzRSOsRJB+0DyE2CA6g4RUSlDBbdQYDvR4nWbVRn8WUS9d1/8Z+6RAV9C02n9B42bDvA7Av
oAiC8jRkoTcp23INPMCmf80x0QMsueEUVG/6Q2Ww+uchq8ZiE6rh+hPx/EJ2YVMrxAINzU7ci4fA
q7wjdkP1G4H7vFRsBH7/OhoqwR0yNGfNiBktiXttQIgC8d2jCXKkjIRG0geHZyUG43+pYmGyMSv+
p55ve7Fxb0+2xxl28vMF9RVwgM5oYHx+u63S55yI+OD2QZquOuUJJRjue5z8NWdcf/UmWjzaynD0
4D6PiNKpfGMxp+S95S6bP6ic8rd1QmpqW5rj+yhsyXWdMU3qS+7iTOgIgJZmz6Aa6FjShsgrf2P1
pWWkbxoOKF9v6Cqh7P1rCaLfsQvasSMfnp36cS2W7PMcMIPyhexx/X9rfBBOzbsLwtAmNDOi04FO
JWiMpYCEyc0XPCjLwLEeiaxTPFBoL+wEdCfNKXGOupsJKOuSbEMeX2Du9JJmMLkqEIyFAPGSufKR
l8ngzHAniShAvc2fmk+Jd9/+ptMOzygv0r3l3eMwV3nYG0lnlAnvOnR4mnS/SOUbVl5a/aXbbnxv
3cs6pZ6PE8RhbG/MLM3qQRmU3dvnIPwoOfcNwI3HiH8lkQs0x8TdIlMNQn66RiLynq1rVfc6s2MA
fBhw79t8pJmlFXdttkDu22mLiIqzjtb7u1Zt6uWJYQ3jzcpir2DsRWKL6mudglkalmJTEXqDBYdU
QHU1mW9c6kKIEGzHhV3/eRsMpjHywy51hCX763BboS95Dy76g1d0FR4Z2zzdo/6de2q486pKEmMJ
Nh1X+RFAEBQoa8EKiZ/eBdixEgR75/4PV7Bd44pLkpEkxu5V2FfUhJV9FmU85sN6PHVHV4ESk+BW
FlNMAuwGGRzFJq/nrSks3KJOh7iH7WurZ7asGU6EUo0uEzLBCZM+gQiSqQF32vBG0JAbTuHVq9wA
vWELDP3jT+FIy3dkBQ9SGF8EArFpHGWdwpSWzrSF1RgMszgD9F5iVGa1X1fNrxNEsCQ3b52TuOkp
kvTvcsU4Bk6GvjFDJoU3Cpe8mZewCt6YgIYdALwExF0zQrI4eKkegdJ670ACuqIQ/FqSB01m+dSZ
10c1wrNjxICk4V1E1NiW+KEFShGqHOVuVx2tn0J90hgkN2zPuifuuWceHAJGbyxD1AZYqg7KUqI2
sc3WbqcAPGEfsPPtxYL8R9hMH1vWSmCs3m7Wg5aINyttceAlAceJndUJubh3hbQKnSIB08+130Fs
OiBwyshj5M1Gz0sFXGSg9krzTqepxyKuyKxKUZr4qAOg72i0ODJM10nJ28ZgXrT5xnTxCcQp226R
r7zr3cSgfCqg3ZaZ3eimZQfZ/1ssNGcqX1aCSzDWxc20H8DbqidxLY1Jm9rhB7X2XhOaJn11f0Ck
qCGqGgdLXHg9jvvkfR8OmWNcUdyFHyxD4tSQXO6EQ49t2cv8ynL4yyFh3yQLDDoiGETr7iZcyiRa
lPsjHRGV9FR75ThzPIekGoUkND3K4Byb5Yowqmdp5xEfsyC0cmAdUlrR6YvqIRzmOnxQ4QtOVbh3
1vX/ZL1gdiC70qLyKVtl6iPsrTVvzYJ/26l7fMMWPzb6baH5yxysoMSAel3t00EYKYwVUNkDyfJ1
fPUKvU+tEmOjDNX07iom7Vm55tFKlvOiCcq9GYDIjHqDFKQ1yN6yJJ+2WX1N6dhUlwUz1TxwiLfx
9xaYy0Gd988coyp9r+ZOU9ZhtWp/HCi/hQM8NSsT9n/OvQeV5KZsdp42pk/GjhJre2gUkxhYV3uh
aF8SJaG0+oHWshyub87QBkxpOAdiOP1rjvPv85UA9HZnuIo653Lt+p+DmWoKF9NcOQo/lwwHos4q
mTEjjYnYz8iocVj4tM8yr7Z39cid4/rL9W5Z3J64pSOzBUBXLfFSIHlytMH/5v4cihpUqyYxUb0W
17ZRu4A1cdKZpyd6e7E4FxR51RH9ydPjZ8fwH6BWXB87mAG0D7a16nN/HA527RuAYNIpnZwoUiec
vl08+/zalYHD9Vyj1swWly9fQTE3Z8Bo36QXVqNvqLBMmg4eL9sBkFg0xEYRtES93WowVifagSJ2
1ZBmy5987qEzh43PSzitYvxiub69+RKe589stotfhGWF+8QgjcXSbhJ+rh2ntMW3WINkcrVUL7uw
KHDiSmu6Fw9891iNRAaifI6MuiDepwrPUKA2/F6Xhc83B3pEoNqIk8n8i+JcFggWCgT464CNPpri
WTKp4xzAGOTD2S5+NLKGAAMkrZy7Z760EPeTrxV+0KdVuuoUT69gOZnuzdrEfvhxrGCFWJg0so5N
Rrfyf2ynNtPPStfdOn9lv7RtH9kOZ3x1i8ueTc1mrCE2VaOS8Bj1oejUXdWUggt31MvZpFm4DtQ3
T4e1mxtp1vMxzpfRGU2HzRNTLOkdDFQ4XMVAz8IkBBzFcqM2MaP+keg1WSxxx4kSo1jcrtqkCa4v
s4K0I63RbfIEh8QE2Pnj3Wr2Pv567TExiDjIogDLAc8PvMdkB0PZ70MA8nm6ViH6hZRfFeB/spQB
hL8+icGtt+ty/GliCRTVNjAvT3CP8Xvn0yfndyyT9jW8z+iSdZ5FMafx5S4vf1rno49bt1WZxvzA
GlnvUCFDEOhzacsFJDNJADx/cZzDKzk8vU648S2u9f322Ae+Q8lx8mQVlFcG3UAM8cJreGCkfrTu
2AQwkh4ZPJ3kXr7MX/+dm0BZrd1POruLqN3bPwW80mGXV/hsALI03YRwL4FByy3IO4XqIpyRjiMw
YLqcvDLBJd3D1yvOIBNHV1o60BtQTb2CJO2b01HozkgM//La9/yoDiyTy2ld7+lGt0RDQ9tzoEOz
OjLRbBteU01Sy1AiKMYmI2YQWyVgJvPMcG/MhVH9IhFQFVG5sKlvNuDECIIHF1kksHVE/QbcSRfT
GBxaF+rTfwBCIkURN2StEg+ZIFPmsXKa9oyAZOXc25VcQjDGkLUy8O5+UVso/bvdHmY84AWjBGz0
OXxSg9vJX+tw4LtpWzJu+JALUES1iw4muka9VH1gr1YjI0f9MD5Xivfs4QAL+ZbMDaSgmdgxjpOr
ipKWaToRowpk5Yw7tEChLb0mKA5UOvS4vx6CAYGbSodB2mrSV3+VPUyxbuYGZNVuJfS+cYJhcOxe
OQuU/QXHdxqyUvhFno5qvzzraJjukhFSj7OZ9Tf61KMtn+MKxgotpqLxLn44cHWp1n5mBVq8fzua
JQPgewngnTucclzNeUeaBnZZ1iSsauXjKPO2+05e2qKwAQ6nl/li/Qx2+GoIMgz85pbva6xwBY7G
Tb/Dq3H1JvE7LPrNgxM5/QWrWTpQs6y4nC3RhxaUxx5UUry7A4QYGKTquj+QdnpPiGcI3C7ZUylO
2FiLMZlr22Xuo7nwQNR8Gfvymhb9Gm4+U9jflQwRlrrzL9MPJW5FS6N84OIneqyMHZMqyHpSXJQu
T/iKyiXoIpuUwYvNnYjUY9CbzvQFh8MMwffH+HXhC1PzPCWMEv24m3mxb90XIpOF/KralWHa3DfH
2pQK69s0fP6fzhWYIgFqoiLWda/pNkFBvN+6CfKSer9uEhHUnHt7U0KbsLeLy2wCTGFPckBYBrzb
0M0EeAgfawpV/xSq65SnA0LZCthuIhif9PuvlryC0bip0ehoR2oPzXDpdndt0arEulMy0THr8BVY
9yQ70ileIezaFq8unf5e460snvJkEXqovK7WjXbkt8LOihd0vMpN+LeMamqC0kCi2hC4p5NUqLde
DiWhc72EcxyFUukxsL52NzRpPA8CJB9XYbZDbt0wKVEIElkHIi8Fydqk+BFx64pNWMxBH019B1A7
6HNHuEKfQaqtPD8SsF8Um3v8eaCNVcWlyUgw6aNMC36W3RdW5U9cq1VQOYOnyL30XhoT+o9fsyZY
Hq+Qbe/xtjfzpJfuqwSpGFXetr3OqThBX7/cfhj4S+NpPzS8yWxuIKcRkszaso6345SyiSS+5ZwN
itgE24CTdgW5l90kH+i0AfW6MAQPGMxKldnp8NQFPxy94mMmFoZKPXX23BfOaI1F+9KehhieAMKw
cuZeOaSwne2QKc/rDdC5Mg3yh+sRXL2GcOmQ67Aljll3VxxrevwSWK3a48MREWFQqa3aA12F7f6i
A1Xfpjg20w/p4q8Qp9C8LFFP5zYyEULojOT3b6upSXjqFFO42IdI29EPIfrCFzuMC9KawzfMarqY
VFZQD05Es5uxkzqVdQKZbfci7XTQSpU5yMHazpwYJHuShxjaQlcui7kmrclJdYyj07ru3KsC9YkC
XIxWra4ixKSG8Ys6k5h3hvKmzuAKmZFHRxxYVcpnSq+wHdXX0QbBwGw/Vt/P+hFSqmKqXf6M1JyX
G+HXdtGzVlrJk922W5Y3AMoIzXBA0/koKXEml0i3/lx6DSVWq70PnPagzWDjkwMm5g1gYjS4hcfu
KvB1NYSS6vfgRJIZkwQGSE55bf1lT5dACZ+ezxN0iT9iXdTjUb/7rYF7DTumXJN9kt3bVxDIjoOS
Z5JlTdIC2aEZtF3PHovca2iE/NkiQUSnOaUWZ0LLqba2WbVsyiokUC42PDwu4Zhp1IOEzYP47eq2
lVYph5rKph07BBoF1XaccTaf3PORzeL8W1CoV0L7kOezYTZJJR0lfRQnDvn1/JPb1LQ2dCR3Ddyw
/ENWFWoAueaE2HCkD8IrMcbktjL0Z9kUEtHoBWd6cFyi/6RWKfk+iD8mvs3fspWLHjab1XlaSKv+
KceltYLpJiIjb7qDIt9oAmKudIeLO3VQ5DI0Bi0oKDb/Uz/ar0ykcWdaiGvTaFp/DHLjMCefVRVR
lkXQEyGU2KiJVBjzdviUOgzdvMdlDN67KcKwYm1zZ3Mdaf+PF0USxR81mnv1QV5MXgkvNomYEepL
40SyzP22M/oYnQ2hzopOc4Xp2f7pKje8u7JBrb4hhTwagKT631U1GyHrHCtFLP0CJg75vPwKwOO+
xekjxePgLTknT9Gf0AY6sBqmbBb9BlMOCwflgwOmlUhEgvumcVL46XEZ2IqcY6zLI1MnMwkZeBoz
dMKcSrs8wpszni5K8K6L9OnIC99gFqB6OTjnv4A2gUmAw7zgYVJ2Hz1D0RegiaToHOk27jUMPuQz
e8gI7hbpWY0bONJ3qgibzECwIXmJ8m3DTbFEeqlMRTmaQR52V1kPik86IZNBfoyWODjA+QscZd9c
wnWohHpYZN0YdHdkETv7E27k03yDJJEqPyYrfkuV40e3ZNbVISu0BEesvpE1FKzxgFth0Fdr0Nqb
+WblU449EvRM+4fuFuUuauI3CdJVCgFyY0jYV+kxtV+YQLI1aWzF7D6XKaEfjDE8J6YtSWaKO7v0
MQA3SEjsolEeREUYkf4OE2a5CJoZIJTBNiZ/+dUqL9FOVo0JxYEYrKlWOpV4pJrfvp87X93i2WgU
6sO0jMrRbV2XGSYVI4lj9IXJafdEl+J0ToQN8KENry0bw5fZtZih0gj2VxyqvgaUCzugBvDA+IzI
aYKeqiZjk9U9dGAf1qwuWLhkT0NlHqcX5pUXt23DD0UMkevoiI+otGeluZpTcnIYPKljgNR8VStb
9nNe7TrvXYE9gnjlfS/6VXk/FPyP+ywR2QAZKkqqEbcx2ENqtFJfKeBd+chAWL+S0P2WatK7oAt9
XEo76VriP+4AQoOKORkKJrENaVPkEseKKrbNeQ4bTr0jbIU9J/V1JtEu54PzMYGc08FzY9eKLY9Y
wTlHGyH3U9g3woJdDdJEYTXUvVjyayfOdQOwetnum3B7+rK1vBoIvpoH04j/pfPtwcYnWjiUeatI
iQc/QMWIWhovWsGHR8lXoGNkyiVQmR+VI3SNtdIx7d4SpBYO24dqi8ymfUgoQkTEXYAtI7cOCIT7
3kfTpSqGzAKnjvXn1GgiSBQoSHhS8/LfZUZ//PinlpAqZ7XpVmp3vRfWOEpj8cvmMhU+Yej3QY5b
VBt1psmxQEnXP6/+GUyIJbPD6QBgBKL6cF+GEw7JcBgtFwIFsRhMQLawUgPoJWJO6D3AzybfaNMj
Lp+hsO6WctENZjc+v16T50vGhc9u3oGkG7MrD9SV3hE4HXfAnI1OtZP0PFMzbTnaYhpPYRG9EL5J
tKqg691BaOdNw7MJnwSfRKWZsQ3MYdtLOjrCrlJ233vxaScdEs35fcam+0Z/RMHb3sch9T4sBXzF
+ZD5tYti3ShaOUgipnZ9exJycIL2tG0002AL1lNn5wAYX28IVvOT9xZixFR7hT0ZFryk08wcsnXv
1Cn2ELNP86LrIV2mi8Du8T+85iZTUGXWtiYjUvlQgH4qLnchc4X9mY4fSRkrLywUryU+QlYtlS/r
tragqfEZZnV/puc9PlsqDOtBm3Itf8Bsb+0lJ+flYm1vQXO/7DPRZnbNagOcv2zd9iXo2ZdmEP5m
EIxSkzEuGtYz59fuB0FSYJr0wWPgr8oD3dI5jJGwYvEojfOWSUut3fbZAe+F/ZGNyXu7vDoDePA7
fIypsLnJUzzwQ7Cvn+l2VB8OF7G0vxEnIs7Dl5+osGM2A83J730vFwJqY1/gKT/2Foqekw+i4klG
Ucx24V+i3WRu5Trtv+8qqkrJxsmHU/fdYxzL0MziRGVG2EOY2JKpf/ANPYcEITGA2euS53+/bK24
MGVonBKsYXkPpAjD98QiM97ahLyQrW+5/CID8kbT6ptSZB1k6zcQIyCpRP2mjKdDniAwTYzLUOnQ
o19NJY6R2h5n2Nm0Q34h2bBbB2OCQnk0zD+Wedfm0WNjAykkZur5ZDJi+WzxgbaczI0r9ah6w9Vs
wuYira0ma+C0ol248lt3fSeQHa91QukhW67hYE901OpafuZYFk9oX8r/EyXYw7Z6y+klwdUoiaxX
HeXgCuYHQhgCNn9FolepaDB9QoQCr3XaRZ+gvK0FmaHGARD3y+cwWMMTQNMwXAaHGYzzB+Oo6W1z
IrJ9NdKJLtdFCuFACW9/Iy5wIWLuZX0OucKcv2ma2G4vVLovEQKJiYCd7ijEKbpSWkrSfcl1SFtt
v67h7GjStWHdB9HahgVyWeTKPed51jsNIO1TwbO4EbIeNwEt+DEmL39mR8vSr36e1TNonfn+cZtv
lfeDmXWFHHYPBysbWvATwf/GdjjadGJEdj3QPqw7HRUjYmYwVwST7ty122LhFA7pcP1RN3uDByHI
+M7P9Wt34wxF4+T/UlhtIE6BsS72BO3OgIp3olkTa+qUsAJHo+7mPUEq50czG3MmS6VKJLwKmTaD
TLHfCcE9rGPUhhSfx4qzVmVM4yJzQdOUV+KxLXpg4XKOMRjomhy1scGkG+a1mfXy2D6nyOFx9OdT
P3xcHK6D0EiDDW9N1jnO5Nokx/CqfyG0WlTzVwY61G+SKKY/cXBkq3fqLn5Wt/WTUoaQlNu5nlw1
cT/v+3ek36VfAvIni8vJSeuBNXzmItXnRT7ztmvhE0Z5jL6npmhpp9JDWtzabsIO59SkPMQVfEuv
WwuUPRdZciwnY/Skp07pa6n6CgXcSvMKVabqGSu0tk+chV7NA8sxnAARv9ff+9kMaAhTusJ1fLtj
4Htaf7pOe1zhEnI0nQmdGrYCyWQlBCx6QJH0khzDLIowLibjJau4BDm1lU8lMdCtytBr4vpGlikt
I0kM67dqtBjtzA6mmctGtVga17kqlXCcwvk8E/o8iOjuUcJ6gTFA1t7Euydesw4OFmOHfKWp0XTL
Da4L7umK3wIVTwhQuaFm7BNMzCrqpuuCzBXwKTQQdUcajKQdXyyTC0KxgZJ8Sh0AeBT3BGxigLR6
p8CrdcKurqpKHPKwAEMXh75AD2bVeRhETnQL1F5+Ep3BsY5427Mi+pnvy11Tf03gVwOU3NBLFjUn
wbwXbY+5YaJbYboLPNOXwv1+PC7IGM7cc3rLxJsB3UH8v21x/QaMtz+F9Cd9HkLAE2FU9JIvuvyJ
ZZ68MLsOKdcMTXExyQVCmj0xxylh2iD67LhFrFsAq4LPGnHzioTXy88t2WFQdoTcjyvTOAYTA/Xe
hZjDPNt49V1hdV4linZgI336XK89J3vHbasOE4kKW/d05cSjxU+jJ3v/anYSrRA3Z0uabSZ0w4Ag
qCQRGpWTcO2hQtH5KoYeALWRdbF5xf7cn9HwH08vMJfL/+yj9niIs/igplHlX1B8Xyuxra/1/kbM
dbcAr6Hu33nKLCBNcc6NFjIceG+HCKv+yRo8Fb7LrZQj8EAwUp8m485ORmEEdDcGeNwwSb7SBl45
NbBVCtoIzyRSfjj64rbEhzGV7dDB/6NgvAQYwiZtVhUT053u17kzIqJ9jEj9Uzq/Rkcc7hRcdwlc
R9SsI7KsT+M0xO8Jm85+i7S6Kq9KnppwS5TOJsjrgD43DXDeFHcXO107w0RkkXKVDEJSSuPAoxMj
aC39tPFQpGjPK+9NnIsCFN7AIjhA8U9AiA8R/X4tS4dY9iLXf4AFlRQOLoL8raBM18Liv/58E1H7
vwJ1xHHij5aJmhiWT/2qaX+Qx6ArlyENNS06AxetpVm5iPOeNPgoueqcnuX+lrrUmF+n8zTL9laF
zI7ei1EbsYjkvu0kkfsZMRoxXprvZD5xf/Gu8mhmjl/NqXYTkn5lewuAXThMxCpTTsFqvyHCKlc8
yNvSvQ8/Z2UMleHe78x5pgfMYP1nkmaWlLQREuNG3MysaUm4Q7iZbaM/YzAvnyWStFybWMbF8v9U
LLXMbg3uKxovNZFObMYyLdNI6RWtGr8mnxCxnKx3+4SYOF2ka80rch9pt8YHioRlSqKCOQSFxOSn
OoCKAWE7/SBhJZ/L9888zkL/wc3WPLFcBGHrzbDhmO1JpfvjuJt17JW5cQgqYgI/RONkdik5eHto
IjmaPkya2jWl7638x4drqCCXKdBNNf0AKuhIbuBG/h+KzykM/slSYTPk4JePpr8HDe5IK9NL5/fd
WXALBbpgiPFmvgozDR7LSe7tr0yTuyfp+w1tizKPvI/TRh2y6ghJ90ibw+qBrvCvLDqYigUR6+8q
e9kjZkLafdgpugN4xN+ZioA0XO+bLkA3PqcHfnbfDavHJEN4SZ/rfROL2dIIsoTrApWeo/DRhgda
LQHe+4pQ2+rd2t0fSstkVuH05aOHENyInkf8IKIiX5e2BdA++7CtouV5zLniwEiRyUk8tyCtZgqT
UQ7dxEWuP4C6FKPXM0Z17ai1WJ3rfU3RRwF++WFce+NOUQYfuRkh2M+OsozXakDYJfWOLAEFOnXW
8Vmf7X2wS4//ZgoXsPgjt/QY17xHr0d9JrB+YBSxZXLXPrhw4V5MqD97nLnWUAHQL5zhvenSAanM
WuASZrfH8JhBoEDUkmiZZoYPDbo274CHIVfIGPa3O8DXSCyZjPxrJ4p2epH4L26y5IZaBbVbb3T0
GWmm4LH3iDkqnC+YtHLKIYh6KyJ9dzDq513PVMFYYRpsB1ttiBi7xDn3Hf1BhmgQegUh1l3M26fU
hNn7C+Y/O5jYzKk0LG2/QA6ADlDbZbxK2VCL2/WkAHZaWSqCHuuFsNfYb4im+C+cEvqapHx0+TgN
OXr4k0A4FtsEGYB4mGBDGt1rScBpJULvB7JEBPIu+RkKbeZaquSR3OgWJe/wuNB7ums/CSSjV4Ws
W1u9m2wM+mPs1yOEnUYrFQr/KZLT9INMjL3lNAqDBAAY/tFJztiTzidPz9v7DQKAylKS4Zwxbitk
iZ2/MU35DmqosZjSH1E7Ax1uTOd8m0KkrEqJI6hTUXumygJBO4tpCJg4Tzdl3grlG6XLUrMLOR1A
ulNx9f3cxPVJl9CmVQhZ2nodNBlC6uX3I7jwTigksO4EDx/SLfbcQssvO2FXK1PwMu3AwlD8JTo1
GdGlLUpVh8luPsSwyWi4v0ELtjwS+1OGDdawKQGek0SwxfVlUbhnj/wQd0ByUdpJ2GKDGuWu09PX
8rRKuKODY6zXsmU0yufIGwSIAnQhsqxlMht7+/H51DRN9ulIW3v/eyKhyzwHWFpOnmaxfV0tkpUT
m3UhPKEf1iJPNz2Wc9r+XBVZ1eOsfQW4iQaNQkpqDxF7E0/pfccVFS7KTEeY0BSCpOeKZpKqyY9o
WPs5ppQH3CaNTNQg+f3SVSdc40Sm4QfmGnjzHl/7aVxah/RtPqgdGY8jl3iqOgybpdlH82nsYqR+
0nGdl2GkGoxZysGt39PksBprEBj3X0BzY0trEdAFj2Wk9Q/+3jWO45N6VfO0c2E4bcUc11fCoa9G
3awr3DKiepvKg498gtiZs33eJiYhX3A8zpXAa1iytJKJH1FagjsyTuQhGNOsyBuWGYa/D4nASbG4
Us+4kNwf45wIZ7L44e+EX7MIGlViJdQkZ8cpKm1vG4xdf+t65EwK4z0M0UjDsn52T5DpbxjdbGV0
aa675hfpUoEwgqPVirb9/t3CeNdV4GUP8ecXzJ3bCJ4fyMJ65CDZgEj+fJYnwkvkRFCo+xTNF6fy
AMkel3p6rvkUGiWzLsAHmBKn0hqjMV15B6MStBHMzLwSZtekm9WZcjr8EXUVbL51jcZOq0kbKkvy
FkNngXJdEKGfZpoZkYOVt7yC3JPZ/r8DWhEuKOJB0pp7IBazCaYqx9rI9Hg+gb+aNCu8JdWtxgPn
dEeL27FLDYtLZ4ArnZWOvxpHZEAx6JWkLFaIvE0Y0XbvS4+KQp+nD3J0KmkglkHIC7YWGjwdxnXU
lYeeWax/XkntXeey2rYj1UKRaUd+1gW9+qeeqLZrZka3mbcstUoBwtkKKXe9WjAa8bFE37f4ZJYF
Ekz4PauRM5ky8Dje3iT745/VDJvAz8lFWZm93zXePZqPc6bh96GgbtTWFS/H0hYp2KYGxkeXU4x6
PyGr+5D/C+Ry4grEj9eqs9a9skIj/no4Brpp73c9HF2TGR0D0izGV/9HiELiT2p2p3YCK4PkuK+k
uq8FuQHBeQ0prh6UVjWrAPjnw9rDQBuGFcL0PPkvHQUvwOnmevFhuNcIZTTRnk1MqLu+rLbWLh3Y
4UYVZAIFRl/griWnT4G4w0uHlBUmeHYc/RC1XcOVFKfevq90wgCfNaESrMytg+qC/wgeabRiMK14
yvZOGhUCwvoiC46A/PmTTnSxXnmcpovAXWVh0A0UYlfv7C1QPhtMuR/9mKkfDmrhcItghZT5i/l3
c3f0BvdoEiauGfx35y7Aty6DjgAPp5jnth9ZJeWWcvGGvAAsUaYwtsxhCXFd158O1LsjEsqtz8eO
qA6VZI9IV+1vi3UrpOvkQ5V8wBoaZZS//K+iOaRvGj4cvPMFVm5WdQxS3PxFHGl1tPVwsCpI+yh+
R5YXN452JkBt0k2NnvyqbgeHa9H/1qN8DEInS3SOOWnVeFcBACVLeo7FSx8iN0j74GPPqegDB4jR
kJK3rqZWksP/9jzHgN9uKxUIsMsBMwRkZIvny0BwWJAN7zD+T8kbfK4GSwoK5bsBVin8OuGzc43r
3bLUci3+krl9Us8U9+G7qLIHE/yY+Ui4BMBOI/FxNLKu+L3ZOS7IDAgHVaW65VdJ2e/HGYDN3HHw
7WR3evk1P4kO6N170hR+4xMgARREiSA6zv0aoB9mZ8Vj+H4r/MV9KGRliT3icC+QU0Ts6MrRoUOl
BiNhkfzMOH6O85duNkt83jTMWFha38EX2X/YhckfSOV13sV7g5XivsWg9UrssdpFZ6Y3jlqzyIXr
WQgHE0CbCvXUKfjmxyd8iEZmhasw3nyeOk3V4dRxpQPfhHbtRn/8IqEB4hhdcpSdRrosv2dyGIQa
7S4OwYi3LFXlU8Ikp/4ltL8GJ2hxbLqeZa+IYPQg+fUyjaE/Kut0ZX9pibp9iRTMsp0WDzMI48Hg
li6ObAtJx4efPnHqJ0fdSdeKbjEiMDrD6IIwtlBQ/VTWoXVGQI0ruhskMgXR6e18Mklb8Qz73U53
oa1+hJkXx3nBz+HKVwLNzfEPJZ98/FoX+ks5qv5D9rXc4uEvZDaZSZ829vKFXXK5/tRItO8BN3Uf
pfqLhhy7YrTWJZTSsg/4GUKiJySCenGzq7+gYB3z3MhA2Y89jMQhPXVj21/igDZDKXOBOtc24scy
IOr5rDXAe23FvZjH5Cq/XUOiB8HxrbyTgVS37ULYh4ys7ZIuw0hZxWWAbrIZfDhWxkZ4H1gAAmK4
kLgw3ijyKN4ugoMi4ui01CMPOkqaJPcxY9kaH9bPjeucAIQ+p1B3wnMAqQ9PUTiLV/B0SarxIrMg
4rFZunE+bXGEm8HVrknEW0ABC2Mpd2/x8l7yww9Ku/Kkl/mNNbFVg4Up3d6uGzBWuc/n9XW9DwU4
VqacqndeGdiVBIWjjf7sgo/vBNbz7tMqIq1x/4UJrwlr3WHGi+W3dNbob/cB0iWbjvLRodqd3wL9
Pgik+cAUXlIiMhYn/xVb7m6YNhiEvZsOSCxwwknMLJDzplxIn+VtszJjewu2g08h1YJLH2W/w3FF
rnvSV1T3oGeriaL8q44wXRbgEvqHLjTqctM/M1VwjY8EB1G2IfkIZTvW1f7dI/emU/3a31cDHRzg
AkMmEYRik83yv6qFrejYv2KmQmfoHyEqrmSjWJjsr5OamoCBJ0sv4F4PoALSQ/+bwfc+rgkYKmzw
r4dWBwkF1znvjrDRZ/wDphMKGTjpUt9RjYiFBUNiQnZu07hqD+IMy0aK+p9Or6k1+PK2NIgtVrUj
AwGFYMtwG2RPhHIv+pqK5WwcKATHF3D3zXK+8dmEDjfPtocmuKrl2+xAWwL/6ncsi2z8lGv/CPkk
uKeR39jUGDTEwq5y9NxaypIKfJIOsxYO206yIB9V6WKV1K2GZ4N+qD59uTmlF6sfI4atXdByODgu
EWLUMl84oKCvB7ow4iuHHoDqGc9fEjUv6mmqzeQBU/oINrikJG0in2g1lTMd/t97pNPV51LbFpSZ
LwVEVA2DB7ivpT0Wudfl5Kld+qa1fgQ8n0QkLBnbOe2zo85dmARS2u6rIMDA2QuOgCVocHyE59dn
thNFHnshMv+YG35e4bki34kA7+Y3L87RhT2Wg0FBmAegMJaliMO1UT00yfrAVZdXRs/60AbjU53g
PjJsOsHa4pYFRgg1GDwpZjQftda/EHaOihfddE/6hqKf8QrIu6YoFPemEGJEXf/qjknpJYij5OLv
Kk2Fwl80N0hwQRTK2b5VNkfM2tfrutI/xYSzpNGt9sVe53HjsRJxRbjwebQkwhgwkVYKS8yTsr+D
bNaA20hnkQXnTHYY1T5N3A8TeOI7/fKe/qLys4IC1sta+iSUfZK+WYd78B4J57/D4Vy21Of1Hn0r
2yb49beBKw86mApAsKoBoVi2XOutkEVAfThZcesSOiE4/AJtPWmqZVg6xEAmt/XXAHmLlSpRxy0u
Ka2goug1kqfrCSBS9awTZGM6FJ5fjeNTBv32q/76g2iK0tv+1Ns9lmwQMit2p0Uk2WZPRXA1gJmB
fY7gPScJqaswCOXtIkK0ejzj1IRIJW1/8DLxwg44Uq/omlLzJhekFvv3GEW2ya1YOWQrSdswBcvo
ynyGaB699cIbcFJAUnyqdX2io9iuOMV0Q/uTTeZLamigh8jh82zOEmTktA0locJAoMr81QNSp6C1
EFTnrtuGNGfd5VwBYmfugyfCtDLKmvMjVAKgZCDAsiqQOS9A1XjKrpm5HWeDHc4aY4n01oaO12OM
ThgNd61pdFbvRjEAb3tXX7/VKSZElLaUoZYkqjcjEweLhnSa3Ex4G+Y70eIuNV6GN3fXJ8Kbfm1n
Ssueco6W3r7i3h9KUD8jEYvB4fsAvkqJZekVloId65OTAAupqsKD2mZI8Gpsskal/QJTxFWmWVeW
NWaPNOiKtaA/BpMLZz6J5MVqTRmCG3lnsmAko6IR8HzboT0PwI3sMeH0TcJ3dIBkxK2C1ty1pNwR
hQ9GBeRy7412O1zhNaxE713vaPrFoWLNZjXsws7WbtxjwdSv+e0roWYHm1TMtr/KDx1tqsN6KTv+
kgU6XTD9Qsv+lbi1rMsmQ/BM0l8KfAcNdpS0ihes/PmlOoMOog0dM/d7cAi/STgdMwTeGnNpQtnc
luLfOg0gkJDd2cTJGISErLB/hVQaBLT4ODUTRvyvWDbTmzZ/jBUnGVEpbvYzzLqq+cgB6cBOTmFj
smqj+M6i/lQ+fdXpiPeXfAxyRG0kWL0f7nXsXA/MZKzaCra7J/TzBegsXqub3NxA5trDwxkfj5re
+7d2IPI4u6OOjKCGTvRsRhK+Kqao8lc3dbMoDltX94wWwFujhFUNC2wWD4qgJhjooS7DQp5YiDA7
NBYEFtYiIyDQ/aHtA9orh7P9UampVQiGVwywSY20sLyQeSblwRNFG+XtYTs6SEMQnnIM89lzxV7w
ljl1xgMQCrh4LkITXde91bPHoNdE2UwAZO3dV2K+KiuY7P+f/bVrJMsfvpodhLrOKyF5IdCxlCMb
61RB+wPs9uEh73a4ZmXqgVEHoucSYi6CfoYfhwEW5KiIdyUrLjbPbpVhXvCRlEHfUKuVrRcuWPlR
HDvtO3kYGBOQaS1A/s3pHLiqef4C+yd5fH7t+Eaocnd2NPybMsCBsDQq5PUazzawT3+6Wvex2cdk
2CILtJ99Q4Q3qgHiIToSFT8nt5b0DfpfTT5qmPYej1HdZ6/ltPHpU75nXNxPEsdeH74k/SxpavTm
kU9c4FSPiVhG/ikMtDIWXxHnGpNXn9C9w4JzqkE1gaMeZJHuSrFH1FdpQBdK6XAnhzfT9Flr3OQq
q93Np7FMjFvFuTJGL+zyHQSu6+cNEa/fDau66ZnuIL0kWUV7AI3RoCLZHj/jjAEyWqt/hQqykc2S
5cTxvzycsm2ArHU7d73Mg+mm50iTKijq/gU7ROgJ1u6K5SB49vmS7tXw37z8WTV8uGvyZ1k8PaO1
LwMJA/fNNF8hGNgJGtJ94E8eJO5BFBU6/SH3aTDcLJFwtGqlGHBB2FUhxee2SGwvYKRIWI0noJES
lKJo0uvob92pQYHjP6G6AthLwALWKwjGXI4w3DFnBkIV+6alaQBPtUqBSTfxODllh5azoN/VWSNJ
glWH9VEC+FuDYl272JvKq+TkTtvI2WCBh7GKj9n2WKJ1m0ptwN4IEQhWQKNOs8T9Bb8oaUCLP36M
ZyH20MZCs1lOgnc91tN93+TQa3Q25GyXFDRI5ah7w/H7RobEesRE0ZcH2Wtu4ICXb9vj8gBPlVHs
LYPKaSs3Xoti3pGOwuTNmXpChfWqLqT15LOUqrhkdNC/XnAhoSim7us1xcvusjVsoI6+m+R1gfyP
rD5RRJpEhRAU/mJgkaik0hoafTZG4+rfJ5FfJcEiX8z5YL3AI0V1IJ+LJYmW/5KT0VkWulqMv3g/
ihj0xfZylBUHSxo5ZEdGtJu1twIC7XUTHW/Umocl4P+QKpRIiX1ntJCdu7at3PCSMl94133s860Q
qNksnf9FEmVbM6bUr0u4TcbPHKHGWGRRSvLnDcQmY23VvGQ/U6myHGVPph4Sq6/qf/ILJCZkSRuL
pBYtbypcYpyNaYfe9XGm5PhV2jvuY3H773V2VaCXl4v7e9iEpruh2pB+4Sa4pfa50lDOZz0o/iEk
rM2wwSLj5NpX8COp6/N7N0CyPZYpwwH+531Vn1fy3L/nVE3fZuqRp2/zT/8XpkeOcJuUrbNkriAS
43t2ODv8fcIEJ3k52W/pAHIvo9uqGRMI2/Wy3exq6jxn9da6f8buFMyBEjuhmLTuMZL7fdjRdBv/
B3rrFYMbTCd2fB6cPE9smv/Uf1Gew6bo0asWyD/SzUoIDBJaT26xWA9cxz3OfqYP+bE/7fPFNGJX
ytOFIYKWTa2Yb7MeavW0457evA2UcrJWH8TotsBPcluQuWrf3aZDkdJhpAK6ks7OX4TMJ67wyMDO
rmjZ7Cx+DgUgTgYdikDVx4UQUbSJexIuPslgGTEkXcCpIRiqw8KiuEF5Fel4ickSaWycsGYR6IQu
mQhWLFk8dT4qG059NP7yni5Hro+kSUwj3WcSx4rdsQPU+u9rlNAMhl/fg+QLZEq4TtMejmJpVH/+
qyW8o2XA9kBQV2UZ4a5CQJ7Gx3buKcJPd9j2bETRNx1qSZoRKqhJcGB/0F+IQBmQI68KdWMuVBG+
0payba/TfIjv6rctDCxNYAeGLgsXABPZGCGqKlhpdxH69y8X7QyYWFbrl7sUIi25B36PqxNdLuif
afxPoGBK0wNJ4nF2GO97IZAbvluFuKTdMEjoYrGsIKNCj+eF0L6U8udUGmaFCVDhrorkgSRh5S1b
lt4svgP72Bw1oTo/nx5O3xgQ+Sk/IGsYL3U64DNstXwe2P1ZuWDDDiW85tbkp+NTRwK8L+BrcoQl
dzJNq4ZdAR2re2ag1TqHeEZlWkriRVFODOMQxdZMrX+RXIuS9hw2KoNBMNtvbuPu0M1becS3JTB/
z9KeYaKOqVZZVK+21lk4ae2gWod19KOueiyLymqzdP25ySC/5V19r9xQbuafKzkVCilzFCqilhRV
RmFbWpNe6qg6COX8I+tS9n5tKhP9Ciu0yKnREymmNXggYWsIBz2CEsNYc1ZB+7xmDc5PuOx8RCWU
dMvN6ZDy4Vk4w5eU1iWIMogdRMwRmVmR1Kgl1oBn7refviJfHrqRJR2f6NA2bN0KQXUWTeM5IT8n
AvrpGVpxearOI/dLLKptWgMICtGF0HoMb2oCJFXLw2ujBsaaC/PurOFsND6KOkuZC1Flf4lyLzH3
3SI0bXF2L+JYI05edly4AMV5XEsLlWFTgKPljCb6N3sR7/IpNBxjd36uJ8M5FRJUOcat3wzDbho+
ct7CdemYxU3PFxacyi2E40eLOFPsM/5dZYVCINAanepZqfbzkAwHsszL9TdEMGPVc99uVW6wylFn
dIB+24LFMLNKUs8kqn1tNNBDex0rszHGrf5o1RHGhEhvuO+1e1+QWJTfM/IMgiCoiA9M5HqdXRfd
VlodTD6VPBTcn3isjTjQ0rbU8EwL4bqlOisSwi13GIBZBVi4Yth5OXZLWAgJGBOeBSv6T+QW1lpC
aMDHjAR70czAEuE1ZkZ0HN3x12AvLLLo05LZt2HREoZPOje4SkzIZewHQoZORzD6AJFiIgSNRrvx
Eu4rt28KicJhKyMrmIPZRgbxutD6uUttKG/XcTiaPvo32Qi1/UMMN5UAO2kFzRJnw+UNZnZKJhbO
Rcastv74sY2TpdKmRBfhXJshn48pz9MrKSGaG9nZcsd5pENdRFZ9203talQyGtRTosIS7vwxJopq
YPsknDgENsWOA9YH3wUqBQ2bCNZjYnL2ThfX4SPqLpYl2LBhxKYD62DXmAqCjp4WuZAy3KjhgqF6
mGj930Bsizmk5RvAvZ5dvbwEvAjkvp5KgLCeNntP12BhGaKpGnFQ16mVDBkJDlY40CpWVFRh+YDX
4y79DA0XNz9a1gc71xsiSsWIFhQgmhByK6fKnMOmFWcrmbvRbE16ATELDeI3SBlkq6id81k9oQKb
Ez4W1FNJ+SSpIiglBizuEKiAtBiez05SB3+E98SGSLADVbEOYBrJB8iCXifJXPv6H6KyGcsnriZT
pAR95oHhmbWUiH6y18KL1fa1HwHkeCFVujFWkr8rvjqnq6T/O0lrlgYcLEYEsUBKo9GYgJoh2zOi
w5KEsGP6Tmpu4jtbSBpnUvjbgfpik4x7LPBxRTVdjXQ0YpYKU2bR/ZtmFhHe3M6vcxcKkzrH9B5s
x6nOqyHBlVkUimTlBe/D3/m569VaaBaMaDi6KaspXdZbvCIRASNhLQ1g0vB3//OUvWQ0/+SqG7VF
CPGweGNu0ITfmEpppzBV74cmaEWln4doUSAl6cbYjsz7aDiCjVOe3a06Abd2JmZjawXBxtkBX9nq
2ydM4+NlPX6MIU6IOeSqKPLWHH5JtCxYK8uFxw8I11Ajp6oVhNepAXt0ESXqEetQUVHOcuvvpSEP
uRoL/HAb9TzbjDnduD/o4TKeS0x8GY+fEDHiQORROVKuHUTQ+MY4XLAa+IWcuTFMJyB92we23Ow+
OZolF1/qVp4ndKI9+la/jbXUsxg9DH5ILIE7s9xGq9oPtB8O4DDehS6zX/+5BAdt+vMzKGasX/rd
+34WcLjTOtKFVEIZpmX9qmEBP/k/uMcLwMP9PrCd4VBnB6+42bKVQ5yIsMtA904CnxEIXtXyNe1/
oRAuCy+ws1iHSWC9zhs5HgVAna6/8jKuSaUwwaQapsnZf5txrdeW9fyrgk6t/wITHuYVpW6ohNun
tTWLkO/lwxypyMyvUMBO7NqRUt9wstzOchQvqCB8H+s8Ouf4BvqMpyDKZQHUouoXfqZURHXJps/i
ZamYMCYVW3/mO0bgn+I7cyxdfp3lRC/CFLf+ITikAakLNFZxTqoB6tZ1IY56GzHMxrRkEZyoRtP7
JraglE+kt/SyHgxf3W6tXIMRJtDC62Mx5t97RL+amrjrFDk3iwuwqQYtIc6WndP9SYutdCgyy2kR
Ep65tdRAU0TXJ+M6KrYJtoejZSW6xL4HzeuGowuUBX37E5XDkREDG6u6Ij4lvyGOzXcVL1rZcL58
dZ8dqLKqMoEdCy+aG7D3xJ7o2Iv4t4u1tVQVbfbJNq2/vkDF2gImu0/uP3oCb8GgH2N1pz2y0fyc
WebT/lYwRycusHJEhGXg/0LDAb1vgIQSvAUhlyLIwcfFFevVq2fBcTeg8y01vi2kGfxj7vEYexUU
BVzlneo/Vyf0tQ3GHL8ZCptpX8I6VjweR14fjIvDDeakE08dD9tqK/RPZCI6VZ7DWkInoRscsq7V
4xT6ud/GzUNP/6C6QHmtzWuklY3AteRCR26ZpUbpOvPSldzBhnr6TiHkwQp466GU2koY4hwtm17Z
BDdqaT0/HjHSva1qGYFsOqqTVcBM3O/jyLx1hJ0WMSFp+VEOV2FjERA7Yi79YkNyiSr/suI8a/v4
stv3TpzjYJ62U87d+fLDPs+Z+XUBApsBcEer6YNBfnyd1RMisnrT8ZxB517BAtK48JRJ8nNCyfOH
hEvZK8g3BJ69o6xO0HIifIV8BdfDRe1uHXgpXU9qQaGgtPng1mubgfyUkpNLbjyT8bZT7iHn9rUg
ose/bd0B4FEsqyD0zbrjBCjv1EU2kfWyIJMq7YVdqlHPSW4L1Ssm2WJjHi3tAjT2A2CVLjYb82rH
NVrIbwqfo6q+gEX3qISDH4cYNyWjbOI8I4XII1SPU0vjURpHPT7OpqGFZty/104qVrB/sEjfVSvq
MJOYxesYIKoYYBz1G2BfBUwjZX/02dYeq3tNxn7yoC10AB3kLif9f+bsi8WST7iqUp07Lf/ArHTW
DbV0jY8Hno9tGzmRFl/cm4C0+B4V4IAr3du6RkQcrKgF1EAmLVaa5OaZQO1AgjglhBlALCR+st1E
EPrDj6RGWtW/POio2oDGiILqbZS8eLGWMKlEd/mX61+dUR84OgZGTnaSbjDRMVE+6Q3J2mzRl7IS
Tz6DQCRxGzy5x7NUCWDvoa/So3LGDRZpR5F4XKFOBG+nZiG7vs6WVgXp9H8dIy1rIsaFKzUwqf4S
dNEfzrfJfBRFm6eHD9vu5B60eAcpg2sZUgXq6dVf56saP6u9fereXj4rlWYgRi2Xy+UoIK4ggYyN
j0QthGHF1LB9p1Emqmzv8Xt0DgL7eH/GIwR+BrPhBYSUF7k86ovhJeV2dTpxybMoclrpHfvOVgby
mn5WdNtpcTqJB3pb+XkJ9rdUIRGBKmhLWVPWOq/cMOmxi2dsSfltSoYrDXzHAfZ+9c4B6l6Iu55V
PYGbcn/hV4uFU9b7/A2REWS29MtvyR/DZdLs/wqMbbLCaUmmjhFSL3MestQuvoSH6H7UT3TSYr3d
XwsJlWm5s3NZ6xKzZ9+NLUzslJksKEeK5h7apfdaOvBuCIaflV8AdMnnvCw+YsY8GHL9CiESrEi6
m+gwK6Rw0TpThH/FDsu55mTAXrOjKRl/253PKwgxAsf+DP9Qw+2MjqE2wnEgmnGW7e6FwXogmeJm
qdxLeRtzoOuMuXpRTs3d0u5LINtC+neYD+KLlS/UBRqx8Q+mFtD2PGgJLp+KplVjHZw8bR/g5AQs
tmP7y2+PJ9cvNeJoSPDew1d/+GuuFLYEFIJULd8Oz6m/8zsvXYLw6//3pGRl68MmpFAhJDElsUMT
edIO4gCtO2H1p+VDFWkRBkvydWodfR1FASzw4hkH3Xmpj+UwmKmbNXUFKA80cmONyMSiw6Q33SJt
Jk3iIjHhpns2A3O/NBcPi7qsvZo5iOeJVGxQo9A2NJbp7ZIcU0MydOUtlY1FHCUHUNGvkpHqZqR4
Je85uIHod41dsGzwwjuVO94OXk2VCEUpPr7KDQ0oWEvkZ+QI0/MJQSA5S5ZfGxGEWyGyptX+6qPm
eAv6IZrE2sLvbErI6Vy3EvEuNKDLoCxeM/0nf+ia8aL48F7jrDkNosA/sVs2rGTehhA08+SxoC57
JTgWlar2NNlSBbIGl8f8Fggtr4qSVzcYeMF4k/+2C+4tL+sjQPfBfyJjAaVcdBLXEMTfWBDW9YFO
okbLg/VJC5iopaRD5yf7lTSaWW03uDtH/QFN3sM17Z5J/SVkr9T6TUBfig+vW+AgtEKxzf6Hfr90
T7YKh8P3xn5+huHFHO3Anbwy9WMzaIAtRHEV2Gjlv0fB1BfkeV5gP1dn88VKnblQtH4Y1nrXdHb9
GuiZlq7biVgqE9M3G8puRI7JGxRIjG3Q+L/5ucYvK12DTCLQ9w4LlVxtYl8oLKRMrvHLtZg8urhT
uIZkssBfdYV9jzl3vA4F4oATU7ZgUxfYMOZVa55ncXIPQbjcbVoSiBHFTKSU67n5ctEmnV5pbzKi
Bpji9prYFW3eZbgXg9vlfMLt8k0nWBLEb8sdJAxeekkLTBzyKVvtMjAAbFS2pyT12+Ktx7t/y7VG
7fnESGGLddLy00ogEgQ82gFNUWKtb0+4AVqD9BNusSM5VQA0DS4rjiIgcPKttbCLMuFVYGMb+bAP
sNhNm18t/FXXxrWblpQtktGt2iQJJE2o2LgAmNkQVmgz+p51s2PH8832WikYv2MLGbYfeDaF03bC
ApE/Xta7JU2OwCc3eUuYpjSEwqKbpyH97Ask2cYtxDueVv+LLF0a3rzzvvcNYNHdE8E3zEmlsC9r
NjaDQJqq0ksYKDF3ADNoV86VelhD4pWvJBGBo7JtJfs9+fRovimH6eh7Ldf2mja4N03cjVBbxVFh
Tqi4YdHaaQoeGToWWpIfY7iodWkqDUetV/AP3BKziosSXDNUx3Qpcq1nw8B6ue5xxbui7MmoYiF3
tk61KX05Trd+FITOVtm7acHe2aRTwHx6ofZZ9hrCEV8g8RTcn1W0XosCCebHeFivmNS6n1UL6eYH
Za3XDVYil5ZC4bqXbwtK7Noh44df3CMlpYZLE81lnGbagc/u0W1MtTN/yxDTfoMfYpnop9KIl+2L
c1fQYKLXCJi2RKA2i7piNmPr+rXtWotH62vDHB77HaZBiQRlFWnh2NcT99JBEAkHvh/WVVcHnvBZ
5iXVTAl0vtc4K5sxaMasxjujmnlOuYR5dH8Khq9vlCPDraN0lyIY+maLaRX4g1nzRQap2zx2iQyh
Lhag0Nmt6tiX9StkEiLfqDMyZOPSfAkwEKGvDaDrPcEXIU0jJUfnq/C8AIVew+8CruyRF6e2pnfQ
lNEod54ecPSMzxOAeN0F0T3/vOMktz/CfFh2k9khT1NGUMl0z+mQwxFRfJ3zbvvpkjnd2dKQRyPM
9iEavzgilXl/rHzIhqfmHwizc+vZVguaoBXhjVaSg6q+iOSs1iHdvYZ5NZUvcQxNBuh3EbT+XTzd
vmeDOW4yJZ/eXfC5UdKatJc9w7p/TOn5P8LbJnAsR6UrvqOtFwQ3upiTiCEi66dTa6TBIghsnhB4
SQ1amaNReT03Z6DQlfryq054aLQmF8HpUDSH7aDrbf6YJNBe/kJ9GVTjDSVs5Oo72L78h9T8+x/I
lejzO3WsrhdAkwO0a0Hxt6jFEgi+GXPrrsQWodo4Q08UflDnOCfe0gNEiFueLPxAfpUJ6Sd9LQlq
5bra+COGKmEcunThZ7FH/Hws289olYb6E6GXC1acIXjKf92/SCRibMQ3KGLNHMw2YQnTO4j8hTB4
HRDGHljZ2gKSwb/dG2ggE6XgpWRUgjufoMFMX+v9Bpe2OZIjxkDvmVIjf3vN7E+FggWPhw7Im4rc
DkvGoThUjjbZ+7nrqo60kTFJ3wShSfEkodteQ9Fk7iF8syEXH/48g+00VceslSWQcEwcjw0Y1BX4
6w0uNpugeHcWzoEZiw6qMb9KVR3cVj8fkWEYvJ7OrGnBZyve4pdTxKKv9nJWe27SWOsFQvccqA62
zMRmocQTGJ+7Gtkufw8kGd8g8dvzssIiJok5n64Oc0Mo1Jj5wmWiBYmUG7etMY79TV4OHWz2wIvs
Gzv/dHZv31El8OP64ajf7oPPgD4CgJSBT6GKpjWx6REPTkSU+USBTgCg6QlISNz2TZQDjB7X7nkR
iTDiyne4Sg7Ea5sbhHutzuQYcXyX2s+R3yfytn/FByMqQ73yEUelWWR+poS3Yur9pV00xvi3v4jl
visavbJxM2eH5kPaKmEjtwnVhs386n+hdmtQ6es6eBpT+lHCb1v7MMAIM/aEBTHiM8iC/nmSGDQu
pGSKwfGTRlb4ogAy3Zjioq0ezvemDuToR44qphU1etajemhYenG5B1W2aG9FjJ1N6ShgSSbE82AO
fpZ0y/FHUVYaaN7BnjKGEQFAqImNHVJSclOKgF+Jei+Y322OLBcEm7OQfkeAQLmhc834lHQ3i2ux
XBSCf5JhGa0gruucy14W9Ai60rkAk8e8DHdpIC98ojmpUnr2plDB2g+jsHTIlMaQvU7IzS1BdeNh
biN+EwCB7c62CKENZVKbIR1vwwv2RvBL6yGg4icR1/WOBY98fq1U4NyHd/r5jbINLL0NfXACh2AC
CjHf6H9BT9GFvGiTOrls7yGHLIPnX9r9PN044OjbdRdBIHuxqFfhrawGfxpU9n3+8YvLeYm/f6Zj
5iZ9RKxXoTkoWVHHNjPtuz6nxbKGHtkQJqG9r0XgFOk1rstb0Jb+Bl/C4rAu6qpd8OnY9zEdOD0+
xdZFCtAoR5GMbKVbm9oF+vNJn5IxZJXZSBBzlkwChPCbS/1Q8unDTW72L76elOj9WomLhekviHjy
vcixSg7ZsIOaYZ+bWrvP7Sjyo4a1hqwcFf3rWzuwdYP1rNX4JN+rRNpgFacfqIT8ip0hqaUY943g
HV1UACHdBcLkITrdfWK/Zj0kcRHP7dQaONAl7VM/rqM5KQBphhFk6QUiRVt7X3oNUZ6K4FCKnWwb
kQ//gptzN1zmM5hf5Mv6qamOkZ2ri4HDQyiySumUsVOB2V/QD1rA4l1/YG2witQK3JeZABTjZWzj
bUA9nW7+ALlPsft1tooYq0JbGK5wtzsoO7xAS7quEKrjqGIbSB5u+mNEgkHyjhsaoWvCGSFc0Pv0
06U5dEp7ondIKUGMN86pi0F6YvKV7accKU/JrixbeF9biPeJs5wBY41UnXvcKH3t09qY1cRKHiSs
mSUUbjoTUH7cSbdhunzbg6UpEGQwnxeX0JUPFlwfQuCNqSxmO48ZhNT1MXYxokTwOTJjeloR9fZv
vbAkIxrc8QVv7vFdx4AEUAR0Ew8UJRSWjvyvI14bOZQHerhZtG58IKCVLnqqQEUpb4PfrEYPrwHD
QQN3xYMum6f+mSRBDhmVAbBsLrnvzWBbtW/dwzuUE9rR/td7Gco+tLQnlqIuYNjF/JYaQZ4sF6Hi
/8ktJUdAdSgEk8yg/pOXcc2OHg/L9Q5GFyIM1l79p7fpQ4kANMKyHG4HCUrx/XmZQJZ9bRF9WzqT
Zrt9cbhAcaRO2c3VSXbi+ajBN9ER+HWn6fFer027rPSAWcevwIg0TNviQxsgQHC0+ONylwmQUNTa
aqA51GQfhWl3UtZn6hv1O7E/FxYvmcT+iyY/7ZI/oHE7pifgxLCdUYHV5aqqKIl7t/tBOJwX49BR
jG5u3WTg+YGsOEPUN+e++X3FL3fi1OZAEIFSCmiU/tB8TCM7R7IF+SNEGiqMp27qU180/3IcTB/9
UoHk/MUTa5CN1v1zAAvMQ1kWymbShk/Or7kQzooRLvKjHTieDa17wEYU456gAjyQxgE1C/xa6e3I
PttEdQxjMPMKagxKFt0OPBgVb917ipzcJvYpTM/x28sKxXacvFDOXx8GNORJypQdzQK4P4ibikwP
lIwTeDACuNjz2f5oBWZL1tgsC9ieWXescApnGPFgu22AaPfofuAJZyYQpfGcB9M8AuGBC2gNLtgr
kH4wwHIanFiwqDg1Mpt2SJp48IYTeM3rmWWj5AuC+Ni0H7FLFILNFxRG+xGNz4Xzwju7wy6BNxEX
Kc/aUakCWbcOHQg33HvYA/ITpHYU/+O2PZjcLEaYjXbkPsZJ9uqTdLR8ttiZTJln2ApsHuL5yXSO
dTrlTN3TPf0qdFjadLdnmzBw10Lv++OyvWc437BKO82HvA4JIsOZMtvJRAi0sXXFNcVfV6ss3YtN
ZBFtYxvqx1IP4iZCDNhyxcgoi+KAUqfRGX/pS1145/WDlPu7IELdZUnuelgDvcMtgOj+JcTOiNAL
zcx9YiFO60bjUZuwhHD3ImDur7l65RQmGRp7uac+ojqb/eLVfeQOBBBk2fhkYjleZr+FiErU37Hs
XAUJdSrbG6T/G+AwdaIQ+uoL2KkdZGAUbLHla5gxV95RFCTavXh94FFUEKQlepLnfGJFYqADmIsx
B5iq8UYbgZgHAnWBd770KvCMM9GD+JciIGgprngAUQvKJ4+oOwwiQMBFLzIavjWNrE6nUYiYgmrh
HqBhaEYOU3jQN9JVGl/JzTh+3n3mymiYXPCg4gNJaKSEr7itNKcRGYh2p1utSm/eoo0rKR5xBmqU
uVa2xJZ5V/+1Y/QHoEIedUk2MIEwQPKdX9bwCNSEF1jMlRFMobw2/UMREjZXtDorhcUfGLQ89dBM
4auqxnv53r+J9uZwKlbeDVi33LxG2oihPpxu5W31YSn0HYsiHmkfoTdlZOmQWY1CbZqrUSYjZgLn
Q/rSpezBov/ep+fibDHvSngfh2mnUnJf+/CYFGpI9y4eWzqq/dd0EbDUjEyOcDZgkPhKtsB4ozzH
lTlbNKn5hFF454Q8pw4vXNPecAsIVtfd+Eta4v3mxSPRoPVjtG6pQJfEbBGHonJQXc2s3HDNTQOo
HgH4UzGDV+Eo4S4/Y86VLoJTKZ4SckJ1U9LGKPVpfENsYZQBWcRe7oyY23B//jku0UhkxsXmkJXZ
LDD8zPN1wvzsxPP9/wLsgA1S/1iEfltMtyAH5y0jo6VXCurXjoOrJ2OQEq4Kq0FgiIz4RLhNrhnf
fTxPdsn8A2I/CWyy76hphJ/IG5H43U1WFkyjp7H+bHvYHWU963rKgWXpLi9Op18JS/SLxPu6v9oc
uS7oAMTRWy2FO7Zh87ncTmAwFdwvqXhdwGX/5MAFIk7XAlC3YDmIFZnPdbFpS1cMZhpWY//kUGiH
4M6QR+2tm9mDcutrx96Y/mmBQAeX886NSxbnPSiSTiTEDnOQGWQLyapfGckEHY/E385Z18EMb/rF
lPDeokjmHPIvyFJ6f/4Ugcp3K++FczQ+gz7EGRIOXJKVf/pFKohpiVuXDl7dLNYcxh09iJ5RU3Jh
0AXRMeCR3d1+C/36NE3oRcmCOB1EuP42sdikJHtwMBqZ/G2QRdhprkK2PTkCzPBFzpEnrjBPjRVU
TpTE/CI76idTR7PlpIfdnLAKUI7FfoMTQDnysLqzkJUxXyF7SuUg6ptlrMk6UXQ7SiwEdugfJBUZ
dn2kjudWnwTRRB+a0sRwe7/QaaxBInCjxveU6fSEJ2wmFvHLJselxEwcJKB9TNf9DV2yO4sEpYo4
bjkgcEVwbS4YSI5RdZOYSLn4xdjSChg/9lA0SjsvX7KoqUAc5tKux0EzanbZcjy1kFydBV/H4Oaj
+Kajn0JcYYqt+d3ZxVd3tXgPh7V0YmxM/zVRikyz6SNLuAP4qsgOXQBsc/l7pNdpxTct2LReGZWf
Sjy6OcYyiM+Ogk1FfI37Ijspi+h4VHN83t2km6yeJ/v8Yf9z4oDklFUsE/dmB2l7xGzZLPr6+TXG
kCVPxPmpaKbVNMv1XSAbqx97p87EdTaQw4jeo9wvLZCF3CMveNdaw/7e1SJWO9wB5PSdFq/0swvd
onjzl886A74lvSvUPaFXQvIc0TeF5pxT6090zyNP5R4RWs0vbWGFdjieXZfmUyG1zfvFWEve/rw/
UOF2ZxsvK3+c8wgD0uodJs9jwodRYe620k1NbaTzcM4J0tn515cVMT7YsnFwrvPIlvgML2CgxOwy
ZlKcNDDXvZJp+iHMnqBdDLeseqx0xZmIXfNHla+B1XhnbWNvGNrolcXOIlDTykY4n38p+Q5k5OJg
+A7PxWzkiN2O8jFO3+Hk0bx4qukF50CNypVZIvH2JQ+KZOjU7lL4QycyXCyv1TH2qXI/DJz2/k48
uwMJozyfxQZ1gMiRdgscqS3HfHcApR50qJBKp954Ms7GMo/mkOzLeMzGrQ7AW+HmkfhlqiNF36gC
5wdPs26KtM7ccUqGbJiXVJWENsnTeqpZchdX+gKBP2aKveTL951mYc5ftFAAEJTfz5Da0QBvlkku
heT+AgU/5g94DV0D6TGoLgY+xO4vQG8sHX0JIX+rAvcvSZR/1ssSKP2j9pqCk8F5WFsnZZkyds4Q
f3CiF/DVL54MqXVegXgiMkBX301uHegtK+ghOmtUzAwplHtwHMgVo8R/ngdRLvYBuiXb4Woy8YUv
KCx3NoeAgkODQqWJGdFQG6fU8S3Kkdd2a4BvvzjhsunfvnUbO6hNwdGc7hivNe8JGGrpYpIo5Cxy
I7jXOS7gox91UBTJJXN8UEskswn4t83bCapy3OwOe86/lMKVhon6lpmuyRIT8/H2XE4E2y35huAg
Esk2TmueUcxmt79AcGmK8I9shtqy+pSTB8J7H3c9NkpEjRIiJgFPn94K4d455iVHZ5TVxdhwF3Es
mY8YqmpkFRD79WgsvS6rhzuQal2p+ZvfsV7nX3uGskXXeGSrt/qxNgbxRG1eULEIWB7A+EtVOHab
fs2HZpYyJtbvTzRP1APvFE6oF1htjTRGjqc5UwcSCn+bUtbYkLl2K6AgaG77pB+V4KT/pR5NdkQG
STMtogGQKoxv1/djRgN39y6EeiJrrOUT+xNiRYWYv0GUv2Mbz8H4QRvClK+dzWJKXPgx8YhYss3G
vYEGgHLOrgsCJsXeELupo2/ISF8hqoiJfZKwV8e1Po02PBMQNBbS7jK7ZfT0JUqKzt7ycuHVLTYT
b4UZUMgvV4WXbBO7yBLfcn+xtNti9y2f9SsWOLnOBXW8BqhmXvmw/zF8BEruLWKZiuVIQwKLqV06
x2b5dd3JyKKQhMCOdNn6vHs+5CM5TlkdHDHApSR/YgA/fmmY9oYK6m51dAdSwg1JB8uxKrB1SF37
ZITcVUfKQzcWc4syxgl5CxFf3Ao7dq69fXDEb9+jj5NIk2S44uI9ZBBfM67CsdP5JSTknZRBr8Vq
ckAmLcwtDK7ZmaW8DCqaFnijT447bc5eJPwZOH3hphFJM29aGtR6UZdZG50xxC32Sm5N27asigej
dzlSjF+b4U40zHK+5AqmcUYD7XyZgQZ5Jj7iBb06lmkEuc8fsQnbXvx4Lwhbh35qA3tTedhRBADF
F6YagMf/ul14VcSvroZ2XYINXSKC/KfJ+BkH0IAGoDvUfx8ke/rDVz9wZK18PH6yze1EzOz4u5AN
x1p/uUyp/o4Vu0q3by8JgPJBpUm8zGFgeJSlGeEoX1wwIsw4i+f84HvXy9bu4g3jfK4cKmK9gLRP
CEmGb9+h+UIg6oQjYfR2CueQafnWk7xFgmUrc0Mc5xOaOg54aVfLGqyyV69bB0zNGJ0HH/Dmfeh1
POV6B03Oe8zXKOFrh0N23FmGXVqrj5peuwWJLC1iQ1yye8CuikjwlciiUwW+lbIl+VJ9rvX0i7EP
VnS/SORRXqCimT6k2iRyoZJ0vnPop5T1a0BgDaqRZFxVsoF3iXo+dRwGlY2pXHZ/+LUcXd/S58cd
htioZ795LBrnFQPeukuIZ7t5tM/0hFV6o1XPvfzx/IlJr3jhp+fuZkwbFhPyOXKLqz47tJj/E8Sy
+9wA9KG71iw+6up+6yVtAHHyLi+gShWHNvYbCeGFiPDMqssD+j5C31HyzDvKMcjmatdjIgu7aLQl
wPwZmMJE7q4QbYQH4ust2ZfJhpN2ID3assgMrhhXlMvewlxcUAwGzl0fss/RajuRZ5TiQ9Y3ekHu
oEDyXSAsmrpotxBrls/vGsSJZGxU3mMJWcDqTcQOnsmjupf5/MgzFX/TLYY5+YAyIUwuMgVDSEAw
HKUijqWMHjRxhIUIZbD0bp0r6hGw3YxgFJCwphe/n9nnb2u1Kpuu9gC3+pnVi59QW9uFJOyBhe70
aDwcb6eY9p60an8xr1ajnidoxs0sJKOgzbD7Scs3zoVy5B/n69PXuvXp6S8yZICTnDYh3uJvlRYT
Lz+gruowYwxPg7RheiunKDsFQedcJAbZ2vqaRdCpZXSrpCCm1UMKScmcd7Z+weXgzs6oxS5W1uJw
TI+U1xsjj3oohxDJlLwYWN+j45xIp8xX2lFYIqzXNvj7rWB5Vxdk1ruxpfCF4w/utp0zkHP1cqKn
kSoscn0psEGSE5Z+3pwhu+wacosrzT8trglxRcXCWTEpEe/or+npJ+eXOzxFEOrAkJJ3LsRwPPBE
KNcYdDnhOeGT/9lyk71GiOXmBnP7zPmt6UYgyq4U89MEmrlbJ9Gc+usf9ElgWINIO7w/ttfUf50a
JILBna7siHSmZRHXj0R9MV3NYQSLgsB7P6WNEX1gAv6EDd+tQqLH8pqrWhJ+uyU5TO2oS3FEgUKf
CUkbUu2Cn5IwCMVzG3SqKzIem+r2kGf+0Bzpe8Ee9+plNslgRe60ZO09+KAh0bPRl3u7LbQawRB0
kamuQQLt7sD1fTGEd/Vi69YUuQpdmbFzGuxZpSEBIP3TQK1XKm2ha6IRonMCzT9uCMfBcHp907A4
+e62rFtZe7q4IkisH2oSBxiLK55CRXh1GEE9sqsvKySPoSjGMUiDNHi4ug6T1n1x5pf1gn/kjVL+
ESdCmmRDuwVjkngKwTiFAPD36SMUVTWO8SHamLFfg4xKtI9n4GSUeYBKRFRDSKrKaC2tIuAOXEpO
N8H0yOOS/c3zZ4fBMtrzdOsIpsi3/58p9tcHiJfpsQkRDfxwaPXedbSvw9ugIbByFx6ZO7dsGTwJ
dDApz8WVsuS/pbu5ANwOE5IAna5KUGBzkMcmWOdiYDA+KzFIwR4+Odkpbd6ueWJ9l3eKLMt/Q5JI
i4WjtTOhbnKEa569vtYoc41l/7FL1UNEoU29vYoLCa4PA3Cyoj3K4H2Yb2VKGE9WtokKFQNmdEad
hD/hSGukZdSR04vVOssHo4CZyWjrWvUCxjPXenB+eP+hYHpirOcbbgVEJ6xJiHAI2EkB8lNGAGe7
Fq/obaOZblc9hyQROJ7neMUk87ODIFS/5Tp18TWCUo93hCVXqZJ8l/ICV5gl9yTeJ/zQNQ2JhmoT
B7f+xyC/2jb/cvvLr61YsIBpxeoHkj6uZ1xOLPM3tUPk12rlMOQhx0drWXxADu8w/ladpmq0ubCX
ldxX0vDLvypBZmBbu8EzfMqGG3DwKMXZtCfbIa0ceE3tNAxcPnZrePpAr27Fu284KpYCQj875r5E
mID8M/2qej4/Lt21zHxm+u23sFNL+sioKud848w4lKivTmPmSKswh58u8A8J89PC2mUrV4Nr9vJr
341CAoN05BeZsylt2b5Q8v8qplB2bAd+NNhYQ0sfGYSfCRVdasuTQ8NPVjkUaEC9d2p2f30+p/px
SCLBx1/zLUKGuVW6zOq4IpAquhAwx1XdjMVF+E2NGVW0DU+kNvW2foYH/PTUoFA9hp4Eys7TBxJx
el7KtQ4ZZwWq3i6dd0PbIQcX8s76Ych0Si/AcjVmm3Fv1WY/R1R1uynd7GkUiv8KeStT79DKdaaC
icJehNGv1Kt+G3kWfmBPm7a7+yemtLIaV7HecmeQtrYHU913vPt3g4uqGcZpxT//DtnuBSpqnUgI
7Gi8tO5UXIeoASiXERIcrVM2o9ADq22I5XIJCXlAFX+Il9MizVXxLIXavQstzghbpvXoYO9XfZGr
PqxCJu56Fq0xQsMlMrbdNwnJgsq7zG3pOZB64AEMBHHMlZJo356aFRNboWZSMMGtpfe7DQ4Xu7/G
CfQh2PO7+Bn6aNd2dAXHqHD0vIk1w+HyWkHGUF9Nw7e+vrdZx8EaDWYkqFclK5VMVDpel6IOAA+J
bTyLEBWiwIf+7OaPu/OSKuSwEISfissjfMt5KTHkcACWlQVMnHRDy6thCKnREOCMkdAN+oNhP6tT
NbfghW6R0Iq+Ep+ppaAWQHHbHm1avUgiezdkGoDWQxHPnN2WdGb0TmfZ9RMuQhBU6nW70vW6wA2+
icUPnhwCUtBFKepl75pbDG50cxlQev6HCgfk/1NIfMlug3aEom6Y5nX1H1X6PJ9WnkaJJvnYuOtP
FncqX1bca/V9T2cBXBji9GzlWaurgprS18e9wObckEnQCoUicexCKvcjQOqo7MfLAs80WtvI1Rc7
craIZwFD5RKLygpsch8PVpO2iEiTuHcZnEd1KnZREziIobp7T0jPfFYsbUcgraGYXnyHfiTRWR+f
cxT3wZqbXEFm5wC2MnAUn2EE1eB0tB6VjWNQRt7iknm5J6hVNfapagelKT8BdjuXTbxH+uG0/zn+
k1gynw8bb+ij4EcL8bYE+tOTq/nnYv5dO2p44tcsIz+WJzx0AlJVkJ7XZtEaWkYUcIkeAnm9peXk
Gdnbx86x1vvsVTlrdUYhLQkgeWE7qewq4IONO62FDLB+EjxXLPKlG+IT97GNorNsq+26HyvSCOi7
Kv8ogsA4bDabO7mHeCEfYtY5Fp1vabTmE7Y8tEvV1lQgL+j916iuPU+B3UOrC4nffVtrlnmyLhoa
0eQRaX/YH4oYeIHU11DJ7rR47cwEiX6WN7sGeUmexucA2eGVdRtkVMnOLGDmO3+BMgXJEA+gmlpx
aNYC04IK9saE2w3TrkhTecK6Ss5WKxiz6xWPBtRgnKyPMYT2EXzpwkeyhy74fQ6aykKa2tjB5BYj
y72kgUZoSu9rB/4Lzhu2+LiuSmzTzFGP+oaKSyJSwCcO4vlFo23i0lazNvJ5EgZDc6i9i4eokXU/
3HFtuJLQpba/63uuLBw+Bta3xK42bXJl6gNNKbHXlMco4SrCzIPoWquRnIZf5W4DTVUyMFOigoD3
u9cJRF9nPE7+0Dkpuk4BcBmxD83mDhqHvd+ciUN66qtYx71Y8RfiUCIGCgxNkK3TLSDieZRjy+Ju
QLUdgDZdHyhqkd++rep48vxEmacvUZ27QsoLZyS/9n/LnldolRjM90fxALkpqLDlXyEQpiXp3FKY
x+MLxCfSYzN7rVWYSL9pXG7x0UmXSz3lM/qCvh6QfbvOJpd6TEmJf0FYGD4NlvlBjfEUj5pLZlbJ
T7aEZ1zFYtjAVnAmvW7LM44m5PgH8vxGFaTP+308u4Bz7m+B2y6mJIFu/fbLQ2f3dbkcHsE12AKi
2vLymzKNDkz3xJ0MRWuKUdKAryYh7lxXXVpXrrACGmP+EqPeS9o6mpRuLqcnXmxyYhTHCCAybqEP
vGfM+PZgaXoHQEC6NULC7u0i0fE/yxJUdLhoYTl1b0GOj15crn5KtGaAZUYSuMZDn6WCDMjtR6sk
xlFJQOvi0qqaic4lx4/Wza22uTtw11+IXcub0qFFL6dPmkQABXv88iATTazhqA158CkbkC8CgNl3
l4xCTwJDZ35mH9qZhKFH28ySZLtCFQOxPQFU/iUJezyFrY2a8O8R8u83dY9iPF44PiHcZwFtUGBn
cuSnhmHx2X33o22kPxC8dK6RhwLAj8G0o62f6+ViiUrjy+/KCwuRu4c2oWgZLBc1kzVDfR4uAMa0
CqKxPTqDqP/KNtPH97fzBEjJqlsW5uZN1URS1m5B4QNSo9b42aDCx8Ax0PS/xgr4mvqE6vyzKvOF
4c3gR2sfjcVa5Un6UT12yimZjTij1MFobXYRVQzmfOBszUL36504tKoSdzAtFBhum7k+2dWo2fN1
b5f8v31yBVJ9BIyy/VEywNWva5YvY4n6NTs7Uh45bNYv+i63zczeiAbbu+ycPgG6ujvBlMuVBYDI
L9GgFXmtPU9tJkiTBEK2Pqzrq2dfxbthzeVtwU+w2J/3y3Zg44PkPvhUA2pkcOMnTU4T6a4K1Au3
DJHmC8u9PsgtkJjJgIxYwE4Y74NhmX/na5mfHO+A1lgjWofuUqSMvdkbbPMcKi2c1TKq03lm71DM
a/5mXyvUTt0GWZ9mTgHN6TFeXBti1VulkYqaSYCm6HlJw/Md3lt5Thg04S+ZwA00ZTsz1oiFGeQk
lbM/T1aFKNm6c3HiMdeNeUG6UTT+WHvLQ6Z8c0Zl89D78ag9XeijDgflheJ2J3p1ir7/2GMJfHiB
2GxcX0kh5dbszLgsz8JJOK6EPHiEGmtWDU1sksR0QjPdvSK4HuSCNI5/ppl3aIr7XY82NEPrAotF
xtp5AOmzo7GoLZrw6gvNfMa1xymoA47YJCWNZ3IvWfY0zB3jzY9VAxZDk9E7iyMgsI9zOyl0KEe5
GgRRfXQvIblrv5xl3Zv6qXBb0lgzqBlT1Jw4dmfenMbZ4r8VnFEmL/Lt/6a2s5X2lKQj7RtWRBE+
ynCFBQ7z3O35pnXIb/b6DAMjyD+y834PiE+yMgS5omGPyR5FRt4R7zgFJEsZehrjelcn8RbJV1dv
CkHD2IQ529Wb1agB66L2R8Pi6pYafbWrHkmV/sYiZQr9R1ZeVObmZTLAaV1abiRq0cglsGlKkPUO
5CDopB1m1CV4NIr/0lU7pQ+zKwwd6n9sbK9NCVkQFaJcs+r0g7hoZMHN32R2W87upCwix+scPB8k
MhcEO2i3SkWmzRgWP1FUnEGvmueODecJ8qpOOTcRf6B0QBQ1FK5rdzYjKsRKn8rBmIzDZCcFixG4
o4DAMrdjxp7AvIECOpAsblCJ7MO2e4Lvg534QEtNQjd+cunPi2/dJ54PtD+jJGL0NOiduOpUOyOM
CH+sPuHV3CF4f0UAs7JsiFIfm3abtWf0oHi4iWr7KXbC8oaMUR8V2YQleM990MNUcJjkWSTKMpH4
/fRQ6w9U63xrJqBQgEQwUXv8ISaQ5R9jtEoUClbOD6DxhOkAyo6175MQqldWphEQ4rOoTLGDBKQE
Xb7yroYys75TKMSbEILyesWAv85EuXpRhQDyf11VqoOtCuVeXoiYk8AI4FM4MWs3OnKntbBAEk65
V08a7YF8JXl3tmvzmdQBnmHSDdCtsdoNOlUUhToQh8Dv+czJgDWRuAg+6B2z/PxiLnoJyg/dkPVm
wCEyVZUC8YbsclqD8JvfuTpzCVN/NlJWZYisWfHh0CJNlzt7pZLs02R7NcrA6rv2dwJ6x+Cxzqo0
lrgFuleZb8UaZ686QsZj9YVH3epW5Zb1OAyzAJ0ILN4t50OjGnWhgzBTuJ5OigV9lViHiJC3+Il1
tq1c/4AM2OoQ4GLq1ngHksfVCZgJVFLj72y4XsqGTlikJx2IGb23xhaWCJn1mX4a+P2+gPxolM1n
3o198IzSF/xwCARIpOh9eZhbmZeotsKfzGibqZ8JwwziZjRMoNt6zVmmX45HLRX/0rUD2OQ4mYFf
ip3tN50v3DZPZtsassRR4UTTd1eIZWcJ2TLiOOQbEYEHvcxpNK6CwtTxT/X2TRssBvadnq29mU4b
uxOKyUy7tpX7gHsW9wXkqVlKjKUMzTO1o9+KJgYPeKSVn1etFe9538m8Ta6XuugkoOykmWDpnqUP
xuremQm1HrGJs8ikoiw7QTQAlsHUnxyPEhFYhsEVZrhTBKJXy/AmlsWU2AJ6bFysqQse+uj4F50O
dF9ZE1KHwyIxngb57BUW4XxIloApfISadqyS0AvhauQBgjlRBaKV6SxYekbSzVIDE36pi9AjDXxT
Pa0sGFCklafKSdMftgBD2dYsxDkEE2DGf/NH7ow9l7FBdMDn3JSVQiYXoPnEsr5+iannrhIqn2KI
pfKAFKlYoMbbcD8tZACD6CSeCjQFjmFXfV7OPA6VhrM4bowvyzsUnYVh94lh2DTRTJI6bGlGtb7U
KAEiiKSfAcP43KcH0zpIJCmzIJvd8MFYaoKCvywll+IkgVuUCtiKfZhWtpM5Eyo/FhQakLg/pfUp
fBeoGyd3DBqqhXMEIhMJts1wAfAAH85biw4vEcJED1WypYSPRWO2+1W8OaytvkAtnuusohabsGv5
aD0ge3DoGFf86g1/mIQtgb+2D9bRihW3U4IBa30EFluTIlSJKb7ftEUoXO3YhAH8MBLqeZLxn2T0
lC7GZo6vOIWVqhkGGXxPN/aPx0wZS8JrppAzGgyFC8zbbw6j3ptrL8Q/5ADCZ64YFEvF4c/HBJ00
PHMaV533TLcf3YsVTLTE+Bi/xwHZOiaeLdaB9xo41RJR7JoHch4qSg8WbSveJeqz2n4CxKQlM1rm
lHVVkgs7hNrao1TYGN0pVBguv7pyM5xmtnx8NKO0+vZi9pFbetmSzo5RhSej2piePFrAt2EauLU1
bdWXlBTKewwhCE9T0LZa6uJkjIojOdf1ueMG7mZ5uIc/CK9yNwcm6KH+Q5JcLLUkwuPhUtjohaiv
MiAyfHLWQnKZ59qU1dZdAnLIR9EWuiRJgqBiWmEi90H+wle6j3XdbLiNQ6Pc3lsvLf8FT5Cjsaxk
yitePmaBH/detSyJRkzK0mfPDH8chy2YIfdOspSD+A4mfkfb23mSx/S9fTuI05UC5gLRrQRm7+vL
80HxImlwiG8x9JCaS8z6wO9MzyXHDWwic2GLg/RJ1fwZpsIJkeofsxuu2IPiJQesacWveMV6P7n5
u4B48uy0VFbMCSbUJh7gPuL+COqRrgFpTvhNjIhbqenwbfOwRvZxh1IBa9Dd9yBfLZrFFRCsJ3je
EXjLvllmK/7kuiJIbWW229hZrrvtVWhk5xSEaXHymYAHUEQ8xpM4V0m4YIsSNec/M24/RItoUwkq
S/cOFFrmMpgxBpxfywvL3mgHJ8/j69J8d31VIfxUUh8AjIjB4DQaEJkwitNCHNbmRVHWJTH4FvMe
+k8IZEsjJ3YRx3GkFuH4x73+j7mHwVMtnT6NgxlWd3CgGEtV8MAtzUPFNaSJOTWjCfALm311K80K
smCOfXNKJ8/fS9J3no1p2jTHbqgx7cg6bRceL1wE/tMpBbvFQDf+sC2Cn8sV8yghjxkrXf2AK9zH
7dNrEhx0mbuZ03im8TrH+p3E1V+833SyFCwQqNhCPHsyaSt8JoLCNhHFCjcB+OKiY5OTp5RaW1MD
KTnYQsP82lEw9oi6eDeTqDof8d6EIw/WN2BdA3/h/2Iqb/drkwRW+taMDQ2Hfw7Tkp2yx60nfkBI
4OJeKpG5zD3bSfGfWxTC9J0HOSgsAPVTmsKThUcMm86zB1zZRXlewsFQ15quFUvAhbCGAm1lSUaD
mIaEd+JZVJ48ubb9gVnGLpDpxV3a64leISLbZ5AOjfo3HpFE6DmWf30bUE1a1mTHzhPJmC1V5TWX
Y8h8lLJVrwb+ODsPCgUebTm88C8DPEYH8WFNFTMvp34Z8pWk5GipQF6tBPqetvKusnaqgJnAA16R
lkERreZ+OijiYWPn1v4N13La66SPDwHePGwNsEncVM5zpFblIeRRkYgD+w/qZ5SXa+l+CYuyTMRN
Y6sSFIIyHqoZywdY4Fucvog8OnutWcGYAYcwP9bQS/CJNpKoINllgc8xvJcklo0tf0C1RUqtxQ+J
ufINuJSaE6kAQRaN39vfaLj9CsgHSxQTyHiDGNsAJz9y1OHwuy2kE3gkeY7SjoeoMUA4NLp4oLdB
+rr06sMAl5uVv8OM6VAY6RP7/v5xr0yLc8GPFzY/6JDaSC8NCiro043RX3hR50dyK2bRTAfewLz9
1GH9n0ygPAyJxkMYJvtHVl5RCYGvh1ui6diwSfX+2LKTXWSIJhwirIFcl3TYmsaRMvLTCtmq8izy
016sNlMue7THyB052V1wJv3sLyNMJ/06lb3KBQqecQherxj6ZT0VRtwrQAXxIrJKC3NYpMhJLUc1
D926n2KTmbaHV43nLx5iJhe0YzHCEitq71uut58tLKg0aRW60bVsu1aOlOY2xyfX+/o32W7ZfcKS
kQMmAezZvs5JuxpXOFSLdKMaUu6nB3IWXMCu0fKN9PRDZEuMmhM9NReMNXh981xsx4Zn2jIfKJAj
2DPkC+Ef1p0a3hX4HvFuZ829jPqOgGokvZmecfUSRCN3GIrlU4UV7+0iUZ6vlkK3XWCSnlu/PM4I
HCH6Mr97uLRiqERdX73e2bfWggbtzSCHNyFxHAABg4bJ/0N9iE8Af60sFkePlookZOQcvO3z6Eoy
3xQK4l+8xj/gsu0MJLxJQ1O5CVnhgytjQv43JrEs6XHDCUFTvBzmxLVUPXFtCFHHnkxWsJR79wqp
JVn+n1FNDhRCRXON3pBMJJHlyRAsRQsiYzlPpLaQraLrqFk0v6Ym+Hnuw/6Qyri17Ed2LiPfe2ea
W4IfutuIW08b3lD9CC3jV2fbHbe8dWq8YunRyCjFTPSRyHkT6kq4ISw0HA27fgLKB4kTrJx7Usf/
ym7BFR92+hw08GQQ7ulroNavScV2ZGPfbB+sV9raCAOfvaVda/R8eZhnDr3hTFSp3gHrMHwc9ZNo
Gd/GsmVrX/RoRZbnW5nFH2e91T/QjnzGIGl1f/J8SxcId6frPhD6MppjiN+FJz8+PjmwhekvylsH
6hg1XNLBMtXOXPb+FXgn3tFIg0+68crNQOgar8uWwUD8iRcgmfrkEoEKx1jSP0yvS7gzVfmCNoCM
571Kj1PX7pg82D3F0lzZMPLuxIdlISTLmwHxz85aYsgCf9CrG1gdS3Vak2/HJorxAMu9vQri/ojQ
0BtlGGIWEhCraO9d9bx2esGm6KJ6FWYW0xyp2sPP4RwepURPJD9kP4nALYzwVdUlxJR1HppAiED4
kgbCsqyZLtV0P0dMIubK8FJhypuKO6drC6SC3+JtjLEkYrnbbXwEQ0GmwxJP8atC3WuDyGsGigHS
jW9FED9t9UEfd/17i5O2AxkzffVGKEmmSyF+t2yu3v2fTKBnz7MkwI4bSO1rryqeblq2Hjw6E3jg
rk9TZRie5K9E5WZ7zpX+uS7gVSunK5inveQWMFWrb+uvZ2MSlgp2XyHSmhUA8fKuJMZZW9IIvGuE
hVn1m6cBJ9VXz+2kIxhrK0C7l9EnV016d+O42HKEqxHlPCONmiiXkZud9VxMKUtB2HrD0tvMt2bq
5HXdso/6Pcv1oKM6jHl1JAjgo+yfgjgPGyiIydXFchq+Ihi0rB5lhyxJP05Ut9hE5tiebYhERCta
HpshiMVP3qY5/6BE8yri/tFKTKU6CxMHIoMYXerB4XfJRiJ6kXzQboUktoFwY7Ix0o+ilFP26767
Y/kX9pqk0u6PkJQmbgYNiomMPfTcY0U543Kzac0MddCDGrXTqApLmmqzNs5/+yukzcatHBsd8h1k
jEfSafTWMTHOSX9hsqadLf6blcAhFccUFhif3V0iCNDTpEfzLHJruo1ljAj0yJ7eMYzjOUH1jNJB
vwbCp6zbvMRMF4ut/4PLpcB9RRi77HlxQXTORxBnTM8O2AQXct9G4B4hYFX5HQtm1xLFCtUfXfhM
yAZOKfxgUcmwUakQyFiATHVXb6qrnL6ctSMPvu4rBl1ZghkD7QXbuZL+C5zEOUW1/X6F19R0L988
q2gZazTFiJReMwmQosuCBOC9T4ThX/wpc0VW7rkSzF6w3SmPe88d6sPR0upiRSBsMlMXERNfunRy
q+JmVzHA1cyWsaFq1rej0VJdDhXbI+WVKIni8OWSVlw+JnHxyQuEFJOzOseYl227LyPIHs6GruwT
DN/t0/EUuWde4oRr4+2yJnxi1ygbuROHXOa8MmwYxp1Jw3x1YqE7JMfTKbSaB6MI4P45prL+nTSR
/Mpyf2pCtqqL1dwCMqGdFt1If8YvEOLAcmkn+tSWfsIJO8rEI7cQjMA8lyJmpihfbDig8SLzzZ2c
hw9YIJzJqJZkH6O5EjXjYdvwE9xM8s4/36RIBmGlrNiVxfr//X1wrRmuQKp13fzCsKIrhMLdW8dm
cc31aUGjvshG4C5uQqbqa4wntimsj8j13MKMMa9lwI3yV3m40hh0ehVHDh8PSVo89V7wch0HBILM
NVflQdl+Ni8MoOYqsiB8/gt9f61vR+l3vMJzJbkjr1KymSdOuaY9O+LNeM0wdVKxIIousyVZebeg
eeN1uGJboX3BIiBb0MoyjGgbGEuueB2wEg+QXFzGyPHMn8+1EdibG9gl07VoCCGrrc7FRZSeO8At
HKLIGnN3n+eOVQ53h8oSEpO08RqzHVC1rL07wcG+SnBMn+YioOLPMbaRotxp8H8qrxCvembmqbDK
8QY8hLNjV8j8KlOeoMCpBdy51kBZstYvCyQIFG2xkpZv/xSf8lC7QNE08DJp4yjBN/cGOgSfl46r
GvU71Fx4jtg8JGxaYqUSqiPm9m2SXVsYlILFxz02uV+uLECJGDe9L6WfOgg38udS7bwCYSv6hWXI
Vg0IGWPCtL7vd3xrrjvfNpsTD3Q1o0XEbU469X/urS8FX2e1VG17MMec3NR+Cy5wHdEX3XO4JQ7H
Wwtht2UPrqAN82xwcP/bdODlU1nQXZWsmqBWCLGThcTvfUUeUIxSiKdMNdNlSD0Phii8RB9extAC
cu4wIjoDCguoaA04KDhfA0HGBoCgCr7u2iB6hiDF+9J8A9e/kBk/WbgowvW8NWaIo4k5CLK0/HVJ
mCEApVct1QRuwlgww1JPr9Tt4EFY2tJ0GTtqcSZ1JOAEaa78A85NyeVN6+bZTDS/HpHqsklPW17z
4cKO6pxBShRI9WumQFW9DQdDU1sl1gt+e7GApyaxPfMk6pnPw86f2s8wb6uKWB6xVeb9+AZJNRuo
ugmMQaQM/D+gjP25Iu0hkRe5CLarrXsYLcj6iU9DUgndiUiE5hG3ObXVaqUfykNVO5Gw3Hr5XSVN
oVt0OwSYmHlZG9GxtmhjiBvhf33fZl7txUO/JtsOYEz1PuieudrlnR5TP/fgd6IrvDOq3TOwVljm
aMbVVrId8TDcIeE2egiryFKaqiFTH54//9iRqns48I31ZzfGozQAVrZmTJCZto32j549ox/teB/a
uXu1sadp7WnWM/FQaBS7RzZI3appRP17+4clgmKWXWi1xXzeVjw4cb+tTvxB28m7G67WqX9gj4ii
5MLfnOzKlyoqJSiG3+OXewnyepmKixUvLuuRiQDIqN4+hzhEj+3QOBylrUEOCOBl0GIG28CKRSnp
ktCnLWXaVHbXgrzWNjakemrBQ925/yz+2/cPJSJoOyBhzQoQ+VKuvz+BlQzzr+gzBcMapTQZILeU
xRl9p1O/noV0/rB3ctGu8yNP6pNpFcJ3+UyOAMddpIVsOLM/qu3WZ0TshSedRdZO4+IIDNTaX74j
UdvlhI6xOht2hySsBtyhmL6/VuQCEm7EgAk+VcSYD4NhxoQq5KqwBztnqnanT8ttM2eP93x3k+9G
dS6Ejp9SCpY+LgOD7YPsqdIgmmLQZF9H8rdzXWpHw0CbIQuolfERJzl/nBQK4HVSFrvEkXNA/nyZ
IHz+uSUue0h1j0PSG7lbrAMf2lrDeWn9ow8cF4pj/ibyPZ/1vqM/jN0lsyqsLsFztrPbzH1Dnomk
yZFgSbCA8WxJK4cLxwctFEL79/OhlJ6foQERcNiPmNVjMFHQGKLT1+4Y1TK+tnrLpiTM/Mp7nQc/
y6mH3ToVKfnqzTCGH5ORN5Kmf84WLNkJN21VTOCPAlViDCHIDp/f+50/S7gyb95m2xXQdGXgaU46
nvk+yKoOOTI34UNLinOTepjv1pY8C8DGRpszJ02qJynYKpU5ZTEQKnk20++CdWywdYFvtvbf7nIt
ZWVMf5D8RRNeVFOjm84wPbs5cTsKRiedMutXKRxPzn8/snT/CvjRPXD7L+1WIGlRBagayrYUnu59
sRLRWYRvZxPyxPYf2eJaLfhjXGndu3o0q+d8CXU1k8Fu3AiWZdsD4hlB5g05njJCZFKjHmV2nBtu
183sNkyD+rx8UMt8/56My/4Q90Kbx1a7YnzRnxlXrJGZbPg645OQCQIhU+CMRWT7NWllOXu5u292
ecb59sMyWmtyXbgmbKE/PXCS/OKjMNPQDqFD1a7AMl1HIYvsxEkNc2SvKsbSQFSFeWPLCyHdq8Oo
Yxc7SUTQgfRI/EA41jFeu5w0kGuDMOw1FLxqEKyGksSz1N3OfcgL+wmp21tPeQ8qFypyMJ/fTWXt
z8QbMR8pDS7+Tbv1GwiSj/37r79kVFlWIfN1dXu0UFokljM235hgmWVZT+jTFuGmYfXGlSrN4ydp
Ve2Nty77rV2G+3w0Gsz6P/O3uY4X5BEz5LDaNguZ/UlC8kUudKSq1nJjvb/X/g0h9kQWf9HCVq7e
bihrK3GaDkFQDyYctbqNUBNiDhFfM/8vM1XczhMmWubTIe7u5Wd+T5tW078/Xs0bd6CWxZInep3A
4ylSDf8sPIoNPs/4tW962MjorCXivUvt7eQdsH9F8z+CkbWauSl1hiyI4S6nwzFNvJXHsfPc/Z7d
G/jfMxJJMR/ogJPUW8VWd8oFtBp6k0tjvb1nnC+8yq3jcJrhuawge92xGv/8H8Ewf3GQn9SoUUpw
xb4cNZKf5R6W01KO2bAWFMO+Vl8/qqnH0ExvGPjDFbsiI5WwM4NTZzrmrD5qeIMvx53/tkFX4Jkd
iT6+GXBPjzf1XYE+TqAEzJ6PwSrwqWj6wLTkmgvdWb8VtA9IfeRjQX8lIOqgEQztYUjRTPqyDHXh
sFqO1RnnP5PdEtkTb+9KAMhqm/RFvw2vcNJtUERl+VrTb6YRwiZRVYbVe2z2gdOPywMyefWf4nNG
N7ULqgufp9Taboc5pUdLsqemVK97ZVZ09+JTuYNt8V2djfJxrneqe178CMk591wKqAA1tCz1tseQ
nCK5eoNYVME7DnCmAsXYdP2wnIGl/bL7iqpF6v5oqsSOuaAZxRSx4MvCvOyLcIdZt5iiM8xheg/n
OuQZ34cQoLeoIbu/eUS/kv7r7UC1/qLbsxE4DKzxcxW03gwpVuKV2cKOy9sDnw8EMW1hoc2nSu4c
hf2ztn5cZ2hTUzulldN/X4ts5bA+S/Jo5n1D2JapucvLzaiyRuaVSkIrJh76mp6zjY0yqtXLgDOA
I81UVHmjMAnK/XYqdt7/O0tHowu/uV0kblmTzvvHFBY7PM4TE0G6etk8FPfJqhyKKEWxgVgA4o75
zmv7psf0p30jBDUbUNJg+3HRlGJs9t/KwHb/os4tliSoZTWvjpSwYYVYby0es/QR0IDKieTuwuaV
3ukxO2K45kQKa76TnZ1mBWATKZedJbFX6RBkMTFa+3UeD+Zofp+xwPqdWBTswKKfU1oqyPntqucc
1LYHOHUiHVNebBEosulId2miTeC/zlKssx94Y179azuZ2BbkJ3GfqI9eIo72TgEYx7lxJd9HLNnK
s0Qe2T5O6siEaY8o/Htm/4KbYADuHpRJDfaxJj+9XyLSbENyyJra23VSWlF7jsaH5qqww9mdZKaH
DuNGn78RYsbRR8ExM0wLtJZ1ipQXR3sxjtJCTalttvwPT3MsvGNYNDJytemZpa4/z0gOSGcoCj2u
hccg0+Ku/Wv30//H/PPGcQ2GUTyVTgDBy8ePBii60jWvI2GpfTp7jn2dLZUtI6IRCE7pd3/PCuRE
Optt/PJFGSVal1luq+FnW+pDkqpDqoz5ahgupKzTcJ2faaCHkg2f7weiOKGeOQ54E45TF5Q2WlSM
cxz4IdWpCLNG5IyDFSl9YrDmnvwIu53vmU2/u5iLiGQeRDGIoqdeDZMUpPnuX/RR0KPLd3CXWtgL
RKJET6V8qXCV0oKK1YGPkDl0K1/u/3YtE8ZdjureIVUosjZCYX4wwyBV6myG8FUD+eYUY0jIb3vd
tFD1GTTiFUcG7fifHblvHF7B2B5qEloB7AM8mgCcQfoMI+J4bmhBCDE+h2gqaoHR9JjM75i1D01o
7gPKjT1f4+Q5rn4dXVCtCuxVmMKXy+gOWkXc2jblJDK0IWQYnRrqv6s5zBUeuImEcYP1NxU1bTaX
KzvZYaRENK9iaI4CS57ynXfppIMWw+t98lmACFdDrLjrux76IaMxRJc2oYg+lQlDsru4orOe6r4l
CKAZ3NUccVHTmSOX+2M4woEkXkOy/xoY7Gv4xtsoe188wjzZfrTu0lil1FEZTg1VyO8QkKHQNZ4z
PJfkuTwU1/IUql14rQxY9k16A18GcJv7/GCHOfB56RLdy2r+hUGGsKUoPp/2v73h6NrRGYJ4Tm7Y
SfheaNdi/pH9SH1OuSWXC4M7XmEkwfW+dtsFDrnnb0DrcMBrZj//te17SWto2XPeQHnKaqNZO8LQ
SXuC1hgEgoHjSmXnA+J2VLal2tOaWt+5nJ4VSv0N6TjAsQLU+vJEfkfMlwySOgOvOx74D/yDyQKn
Xuw+hWwFku4gfYop2+iKPwHqhfIAnZ1cEIWUsXczVpPDKBduHhgk+hdsHKzNOMMalx3of4plgpw8
L4Bs1au1TIsTNhdO5C+OtxU+5XZsri6MNyQILpf+RCk5yUMz7ip8MQujPDPKUU4+KJ7kz0dgyW4V
UbavNgmCqbKarQ2Ru0XLNDd/I5Mr5qrivCYnyNXZJ4owIibB+S78J4ZmGd1bsh0s4UDZtom0HiVs
edqsCvIpWONLuPc0wrhItAjvrBJZ2y+hR43Q33ra+/yNVYZ9VkVklBhu+KNIM1UuZ+McH4WDZrBd
TsjP36+dzfhAhQz4xPQtNu8lGzZFU6T60kRj/YA6G5AhbTPauthtYdyDZvz5inOUIaVagHO27drQ
q/0isiof22aVGRpA1FwBU3SGIapRmfu6Cfnq7DGVJxBNSctUrrLGJVDUFuB/H4sv4bSlHLS9mWqq
ItitsqDjfk51P/1CgJOL0Rrvp4OCxzbQFpenfgTt2THU4vysqfjycSHM0W0qnOG53qQpvNK5FNKU
BkNWuA3TwkmO4y1VTuGQqwFLP/MPTFquguuKI2xDq1WrS3Jfy+Yqf5xYYs9HgdvM/2njZEcrDEFE
rGRv0vKyc0TUmGfeKZzJ11olau8DYtjUfPggMHU0HPXQGrwsjld83muvvVPP/vWIiA7RTRN+vFlP
cXVOs2RGdBwRqtm91H5m+EH5Ty/D41T9J3J7qBeR2hGXkvM2Vx7eG3qjcbG/eh5by/UWzOZyFQJ6
JyfPWzsPl/Tcm4L/Ksli/F0zvDi9vSNSbLNCc7/D3E5oCQwexQPF2AuTQa1uCg/ysNV2mBkzbSZI
veLQtRgfTbQ7U6ADA0aeq7YbDrxSBDSqNWGT1atyeXBMdz749+EQE7VAsaJmAhAIGMVG9+xCvJmw
WSKa7DZVq76CJ85cn37Rb7OEL63MM/nKGsqJfx8efn5kKPKQctGUk2tSrEwn5dJTYataPEggzoEj
QueHcJ3gew+B9UY+VMl2nNel6JUVul89yJkrZ07VBb/cKZyIsyfIijUs1G21b4MPgpB7LoAua8ph
ibZLSlFhK7m8PVbwIcwxI+nK0hduY09VUbHjNR0l64DVOvKUMM2fD+bcOEacUK35Ojmck/8tsZou
FBOpXOlV+hYeZj2dZ4AHUdIl/vcwm8Nq5+YP/mpzEbThnWxOaOwfRgx6D27uNG/k1Ecbrz+QkLgt
T5IccVr4Owwo0Us8wcTzIR37abuwhM82mo8MALtr97BNGOMckI7NK/eQzqfLdmfCep0NIITERDC5
zrcijJXdvZPB7APTXXVOqQI1kA08nEVlw4UIj3b+hCqoIYFbSD8J8MXIjmDOzmrq27ZysXoiKFB5
euVspd2l7D225Nis5hYz0LHA3NF5n3BfBqFkEGylhHhimd7v2A66EmyJOKnWdv/k5bGnjlQFoiBD
UPWdApTJ4VeiPhvFo8m2QscCabDHn+wAW2haDAwKoQ9hlqoZe86GvGvF+h1S0jJYU1rhcczL4mtG
6DdljxdmW18qJUp31xWM4+cQlvRh+KHEip24T05sN7qjYFiFqP3NgmJPIYQqewj8kW5JrNlHjnus
wDA5kaMBpmofxcBdNkCVo9ZrQoiBL/vYD2WVmCEwdfvPtQqF2HvP81nDSr02leLaNNXGyaeCE3XW
tRNe73KFV9YSbaCuE26tde7Bb4oYaZ51kOUIt51VWT6faCgmJTOnQHFEe12mdKq0uj6M3vV29Vea
Lo2GI8k87Ch1Fmh+/qjol7yXs/njV4GUYccAMO8vTzMYzoo4Jl+YGXJ1wxKxowRvyuCpietrvGaL
ny4YTd8s//ViR6TBT2hSaxZpGL74tgrrp9UNWzUzpyjNRSTKFWgV+Ely8w8qvf+R6q6ExrtoihU+
bcBCX7R5a0zdy6DceoU9eOWDGIEI9WzjRCC2nYLMEohxdR12dDjGNdUbGUVvoQ0krxLXoKqZVmKc
sUt0FGM4ixdL0cZP7S2aNWioBiKMn5ZX741PSxzupNOqUdbo0I5wp2AM3lT9/ylajj65MaLSmaI4
+OXA/2fqrVsF+MPD1IaYD2Rvs026bxrgTU51tACSkkMXZthuip6LDwqxW432OZ8NZ0sQtti9xqWV
lYoIEp9HtG3bSSniqCZFRjdQ3okCG0JGh1QpM1SE4LKBF82omrF73L0o8jwGu0AXKMTJe/wyltR9
hhdtuAa5pqjx36I2nhiR58whf1gUcrDkHxEudzOgP+OT8MqBtWd4BoTpefBVcmeSIcULcCYvZU3R
mxrrdrc+CVoiD8Vk9XVniIocbScb4PHerTRvOglfo0GXWiN+5GHrUlIPQoYiuzdIIhv9hiM+9eGb
shs1JbNS+sCiMYn/z0kzZyk0JMW3Vnt7GXPZZcCFe4A9WoBFlNL+vwZ91A7//w1qh9ecmZWPVMOK
0/ZUTUIwWW/j2zUijDckxK1+4ekFdpbvYV/NCVHRgCUsPFw9IFsvYnAhiPEWLjx/ouB+nyn51wDG
Gxv7amOdhSjN8aV9zrNXBdcN9Q9NVcHgqm03Dz5QrRhdxhvfdvmN4R3YZmGsoq9GwKjV13Lh5gfM
v/qz8EpKc5chv712OMWOBx/hhsSvcgBSYDweungQU0QHTgpuVRklyZjAnvycIMTDBnIsdoyD/q9s
6KT3/3HJfYp5qNLwzcUnYUl1YTO0vlun6AKAZubNaxAjTZyj7wyrvs+ijdLcCPU55kFtdMwleDA9
irnXDpsohj9INI4mY8TICJwXULpDk3XCxk1TCbVhGCmlHufd7qgTW2cA5QwmVrqXK3OCfkpWgL86
GbQZHMwJ9X29NzA4SOTSpSU3ZATstC5YFbGpWE72IdGkWcLLi/K3vkAXV3ETBuf9B2/9H/o6jFr6
apwy/qsezlXgNlhnALSzh2MkaxoLTHtUfuv6P5/3vDR8QLeKu1ZOQyvYnk/ZdK9C4Opn5ZnqfGd2
GhjS2WZXJVbHjupH2auzN2pLhsStp8CHjs8HBWOO60v1hdi21ruKIIhbojMJb0X6q8Fbcv1vOi3P
V4x6GkfhxIjxZAcvtGF72+LSUdnPPLtgX3G86oi6tH6utVN25HGfJJWmy4e1xC5qTUNYhT3UXohW
fJ7tvnprA8SQ6IP7Ta4GqsoNIKSpgAtT9rvQMwJEWD95VooGJ0+ubLwYdtfFfIDYtDsNGllNi+vt
vkYtZTcWn+8XkT+EuYJBp10i4ovgCrFdS0QuzvN5hAkPnKDKBko7jd1MFrNc9qPdHS7ZPXbTmpBg
epSsDhcpyrYtV8asSNF0rdVjMy+qDbYpR7C6zhIZ7KMehblR4Rlk1kNzi4cMsPRGHEC4zFysrlUg
0VCNgsUhXcgtcunKe7rowU8yWzmso3T9dHXQhkXhFsFM22lckiISEgpQv3xvSd3lIeOR98UfMr0r
bPcuOpZCVZi1aWVEmZjRTVUD1V9Od5lubk1lmPUB6G33QiVaaKJFgWxaBwRn4+OPKlhICXa+ycgd
JcrOcrIqrQksd3sNrVt5oqUB6hHXNitf7h0+gGhJGLcL8TE9zltE2hqiHu5fs0F4DTV5HOLAbvSm
ynEbr/zVtXrtuBudnxxpfwMDuBt1R4uAgSbjVnD7Z1QamGn6KY0O7Wa9cj3Q7b/3oXvqRbfA4kB5
Z6aQBvblTn3dObpGyqEJcYpr4helEJFwPm42FbwzQkbOypT1nuML3PsbOHDMFWdBEbe91rXtNiZs
w0ZY8e8Pl6w/aWHRP/jPlstFARDKXHEJRzGQapLoWzPeQh76xb4ndsvFCke/heYJrqjkNXOvm1Rz
i6c7ukGa+Uy2DQm+7N/Kh1FeD7Z/aUsAGteNhFMX+K+B9EQ0P3fPD2rK0yG1RZirm4RTzApAtYME
KxUPqttYnDjtaQvTMo3UrBB5e7DTjIPVjQCSa6awan5vmHiFcTufwDlBKdBpzaYyEb9B3LwqK3ic
UEYpK4hMMlBeCWWOKdgRwmkd4vrMuZzru8JlAeAoHDYYI+RpG7vejs2+lvO5D3DdGcS40FB2a312
VV6feWnrphIPLVN28YSlO+fQpZriXMxjQHtLYj2bwmgaWJBE2mOzbdf65Mt1FeOqa0wKWxBkxRgh
moWJjOGCXNUVfDShH3mbuZXMBrTfLZhjbojYJLpV/FTdsp65/Te8N+9YrtXT1AqpzYiNHi9J3aJh
MlI+S2HvXMd5KdKE0irgRbX74lnnEvQoGGJ+6YszGkueiG9DMgfVZPxKT3wZCwP3JN/m5u0D7W0h
b7qiy35f53et8XjVaFpermMJyUK34xyhqsh0l0mw3HS7KVEhZO13cN6rMVkwCRiD0nPBt9XH88zQ
myfR7QtsYERNlvXlAxiH3l06isKpmVEAQeC3YMV9i3wmZLiSWu0NdG2U0WO9KHE6lj97PG4UnwSr
26Jqoxi6N3tl2nS8j1MR23KAd9PmpV70WJec+1UKDS3syL9n8xKZC9EU7mRChWkKJQBuZ9Ez9eta
LOkh7cFBp3uOB6bdwC1d0Ak/51Z047hx+x3y1WIeheVyQhfRAOQpIyENrKcXBvPfGAwv43htU5EB
7lN1NRMjqz9a8H9LJlz+TZUQTzcJGyY36DA95ND7bB9gkWlRImXc0WO8m0AVNO0m9gD1uwo5nZJF
VzS92SotgNsN6UcpOcI5Zn+Ido6m73XsshtfhdhrXtNw3dfChz3wXsnDSLyqPaBxe9FhXB46Z9pr
0CPpxjKpcGCgfJBGzAjG2yZnc2RCzhLRLa7SMhSS6TsAe6/bjK8N0WRK6Hun7BMT/j8IbMrsWvlH
vxvcXN+hs8LFAIXE71G1vyfXd2hsMtsi1DN/rWXa+y/s7029+2B3tOF9SduyMybkJjPnXAiM8Ego
zxaLx+NP7Iu6icw542M23blGKVIhjOL+qGFkfxkra6xEpbkjIdaY3w7wOXKBInPzJEdP4CEwVwTC
FI+e/DHm/A0R7bpNOIqgAilxJD7NToYH1He3+A39+ksyay/XrBL+Grx/Spx3YHaSggtWmYnzi0Tm
6moPeDpONi9Vz77gpi92jcRbtQ3J1Jme8z+k12s/4HmVdyk/4aI8jNOUv4eoKphBQ03mIyLrn+7j
C0xOSNz11EWU1Afq6Nw/ed8jNsDWz7bMoj45aI9yZnbk8nz9Hw4Bt5mmrdNR7U7u+vlLxvVCsCLV
FcRPbd43qC8x4yfOT1Q/M3Va4LLrziaye2TdwwuJ5vy2O/AEJgt41SRw8HQ96RtYJivSumOuHcQE
rKZy0UAJwtstLTKA/Dwu3+Dt9SxL9Gg4Cnjn3vBNxJlFS5YMdStzvtbdxtqH5zcfcFe6g1ZafrnI
5OYX+YMWsUX7ZxsEju5BjYAujosjJroieiODk35sEni/ytNNFf0uTdT7uxbzgHzg7VzeNyd3VtSK
aTPdqJZCLI7LvgszDhjhXwu8wnoBD3ZXBgmwjmhmsxPJ1DMQXG9+cA2i8IidVeSkEy6mkfkaCc1B
XtzCANhHnEy5vQDynjWF4umpiAd4bfRU/VVTXwSTpPx3Mz7F682s73pJrE2ODfqq8pNfZzm9lfo4
Z0R+xRh7Ygs/frdpnAUxLTj3LRYidgmG0BgH1GI1tLvQDySBpDjX0aTLUb+71SiPRE4i6Uh9zjjO
AD8ZCTPyaU2Ct4GIgOBduP8K4pG4+fUawqj4GharRhETqXTtczJBST5FAMXIlbMD4/X8BHf/AABc
acfn43IM1iKhTkeztPStQ2cP69Hlrpmm8TOluNLi7V/fZJXSi2e5VMMo/ob2MKFm+aSwSYGUpfhe
z2At58U+QM5B8Ag+C6yjkAQ5egOpkZBstzC9r1yXqkZmoCx76PWiJ7RFlYdr32DL11W3XCKMhzFj
HzNtX+cjU8zNbwFNAMca+/nqT6QC0CDap4Wwo3VWHWJHrgU8GvCnMe3JjIBeRJNrEgZ4xmsHAEP0
tJ+F1Er34eqCj8oKjMCS/NBtL6mCo7jbKAvTjzj6Ebx0Tl6G3p8D8JYDCyAPjvcY+5qG2TFZlwhN
xdv4grLhY+i7ffTCe8OH1/e5z0aBTNhWVhe9RH/orZPZB9TGz9eXrT2PpVw0Dik7M0OPp6fWbxZT
2F4Ocsiak9Mr+izdJ1wJVCWhEt0djAIfcue1qb4fDMyqJvv3oONbHOIvHy2Y3cVRm5b8y+W58V78
Mv3TUhXmgclECFnKrUb8TQq/L8l1L/+/mCMrF5bU7eQne5CaxyMQfKEhG6ckGDH6bXEWqnIlCDln
8G9p3yhJh3QqSJwgKkqXUOzUQwbgp9KWXgg4e80KaPYRPVKEGx4kMv1jsgixL6CK2NYdHYEjuw5f
AGwi4sz9Ou1pegBjLaaFXfcC+mHPbCfqPYUZ+sOVpXuN2uBFX3bdM5pVpJyRvfF/LX140Y/i4m/3
8RsthkBWhe14PAdVJJ0h4YKLJKrMU7UK8mxlUElFJpH4Y+rqV58ZYgizOE1uwTizL5neMfdClgqi
ULJyrJct10pm8gqRbV4/i5RTFt+px+pWdIWfaKOnGd8XOTmzAA+8dEf/U3hiC+bkFrGECzy6VgPn
MYIfPBAhUn0YBzFt9i6VnHagQUQ3f0OHPwWT/1kIzKWuazmM445kADZ/liGSOU6xbQrSIXZgX8Z6
MUQvFbWJ8o9SrWr9ZqVDOUOXTL3Hcgg8z9SPlPlJJ5i2YmRi7fEpuu9RcCHY7pqnsylYJg0LNF2v
zlSg8rRxYL4PaxIaMbcEQuOvjda+sihoVnY+6ThlVoKC/RWbVcMbVCZXqZ/IW0Mctd3Lihl2FhqE
kIIwEnxlP8sIzOJgtPqs+7sHB+UWqncb+WfvMyBZLQPGYm/LNzZ9Od9/61Z2pxdLHr0Nc5/sW9Bb
2/oWbnZMPF4TECWqn2CR5LE5rS/vMAZlEvmfxgTZBmRCAzfG9BcMxevUUQ8saZWGuk16nV/61bDX
CqDoOqFIb5wDQAH3Nm1hKrikyDGmBfwjXxwfz/KJg5/sVzrUBRBrwN8grZTeC7kiJ1WvSAs5MME0
npN0CE7eQX39InaIc2FSWKjrurpjwrEMrAWbCmu9mjmENMSQDt0GU3e9UX092Hd8YC626ulyMNZ+
ERIWViA73c+tSrVEtCKeU5ynVVVXnz1II4iv9rtqhKGVN/s+puUTIfo3x1VAH7Dqk26ehf0+regy
nQko3ePkMaJnPnGQVr95CVHcVPILLYgz3AtunaD8jcYbuv7ChhnL07y9o8fsuIyIp1oIpgbWYI/g
IoYzv5flg1Gm1raDM5+EJ9sT2JHRaYvPV0GLqUY/HmZJ6IjbHkXdb1fKNz7zO+ALnC4FFbsAv8T7
XseGSlxCFZDuLBNfXDmNTEQKcZRE9vqTN8faT0DJQcdjnKiSoyNkiOvsIp2jJDVMw0f5Hbu9p7It
qcsLeymL8xS16JWPVMF3X/SlL5+v1ppUpb6x5Yk0hJa3G6Qc4cMAkXz9gtjNN4N5x+MrMuwe63QO
Pol1UxXGCJ6OnhdRL5JjzsPGI8tTYJ2vxQ8u+SecS870xsPo26gqCAsqZ/inpFRAFTbQSVgQOm9Q
jYD1nQkNQO54GO481bwKaDDy4H8JepddaB48Y0yN0P/3LqrmtIPU+jEJpoKHkCUGlk8pAe7fQxPu
te7l9uZanEluNabqg1QG06D9J3b1/jnYjXMb2cHaSd1QzhA6589+xb0D2iegGqWxiAexfZBL4pFc
1dX0JO6HNpXbgbwjaW/2baRKhwV1fc5SOJYM9NtOG4E/cVTTgQFGmqBpivspn50bJL0v/KGOV9iq
aDcOUljZL/8qKH3QMxsmdBXseKlaVobvgpH7dBO62B3PnfkH1NCeaBcVJ8a6fZC29e4oVE8q8uVZ
ht2AgZ3hlGDmRfwyex50bwdIicF8w+v9lYuhOC0PPA3L09+B5MO8PEgYfpr/oGsOzt9GxxBtm4YZ
3PvW64jPrlzJA5+GHDFGcy6Cw9eghkpXyGkU6BjGihyC+DCERX1qjqyS/EPE9+YZudiSQtgw+rrJ
TXyQVuCEUiVOJMH3FgaAl0AC/ezJ9JXT8he43gf7wtXk7shdjxd557uSeH2WEQ+aAhqLBC06tlb8
FoxKx9jMHeTdHupsOpGGHwJmQppo5dDVRFI5bRTM9VK8fXcJ01EU+4rpQZHCL945pvE6ou6weZuR
mGtETDPpLZvYGhmByjfYtD6n+0Vs1h4vifpOZF3wXRAoFSUsg4TTGAapySStywX0ThWO2fCgX6A+
Uz2eS6kLoedzPs5pTOwe2n7pJBqTg3aLr8BOxPQV9och6mudEMR0jmmLYeODVJsJAYQQrjGbWOYQ
MKyrd95+gqGC2dDlbrY3JKzOWIrJzwpsvakRNtjYLxQgsbdYU/aUmGAsZ6X1R3N8Kk8thCaaUMzz
KUqJmgb6pnm1oQrwixjCJp1c23U9+WxhYwBwaDkrA1QDsH6W0TD4XzpuR0TMwE1YNl2Fj0cG+cmC
CL7LHgMhDsScKGi+dzCrjgw+XxunSTi7CWP+wisDWJ3Y8TTWw9e+Od1PJ6Y8kkbI6XXWB4+Qmu07
mFRWozJf+lrKImFeM4KBDzx43wtWzTjpdf5p7d5zGTpeojLfqFYH81+U+F21E+EZw2ETWHwU3bmj
tykYJ3Y0oqujL4iZIR/lBbksI4GvqkeD4bxEvHSp5oR4d8GbM2/w0pWWIV6cKakb1rdQMDiVI1JW
EqClWqc+jIBbV4OclToX54nqRXf2UMOL6HO+9preO7HUlIqHHt1h8sQK/i0d/pNVZmKyIyLmqXHs
uWloIs8bBddwLDiXFYbyU++jPZrLAfU1ior8uXgbYQivi7O9S2EohexDjfsfv6AGQrH8/6KiKoeX
rKKFw6qADo8TetupbKzOk/tAAU15wYhA6SdCyOIR3fkKKbucUTviitUWwY1Ljk2gNGDxheoosM36
acr1yap6yyCFNFrMko/pHJfINAhoPOYBRnIvfxD22SKEKK9xkPcw1D7M9pS4Pzq7X+06beSv/exv
3sNA6G2Us+vPnze7EEazjJJVQvLZ1UvzeO7uniR+icnpwHxEW4jB4vrBsOYlrlJp6vtCMyB0Mh5Z
63hWaNCphBf2BBdUe3wpjz8i3K7ClzlygEedRPknmjCF1tA4WKi1oePYh1/I3U66KYug2ItZG9j4
gDhthX696DqF3+RuYCknxTIgwrVNy3GCLBRtJW2D+G6dbUd1AnKHPIvQkWOWhmFXIF16oTo8Ss72
cok1TUvSRGOGX9a7SW1ZQciXyVvRRvLD/Xn6uNRaehSHbdepZ1RvNpm/oUqaI+VFSMQu4TRiDfdn
hDl8xnYR5cslZKTkmwnUIr4g0CJD69jiAOJsTsWYqmjwe7brHPWHcvcThiWNMcaFQCKSB8qGRhc5
5m5A54W7fNA7sAkb+T6dWMpdhiiCtvAzrZMjAQJDb1AYcigS8/kSYnNQ6tDDxGGao/2pZSqNBtqv
+N7KWqHAKPb/ewE84g+sd+OwCmU9Gs1qO/QmKdb50tQ1ktP52194EO6mRWbAzXEMRYzBXwFJn7RH
bGqjx5qQDlC0450N1zX/p6s12cwE7YPQcfG9ZK5jAMYz0rkEBQN2H9cUUWD1qHAK6PXWQcBNgPt0
H8CHqjKPdAzScxqD6irVgxV1sZAZ9qPJTyDaC/KwZ1zkmYpNvhiQCgT9+200/F+CjPy3M0UGMOzX
mtppnq81DWiV2Wolv4FWQdKzvz/W2K1OzsQWojyrc8DSWKwX8wYhEizJ63boWJThNbAHOq/dBYxY
BDh0xrO1Bhuu0JhU9/6PLwqotbrOpQdyZ9HMnv55Mw+Xwd2Cs65K/HRDvZCsMe9GAouJO1qKQD2/
nfz/64LhtgwHPQ3xugqWrC5jOHVXBt34NmbcRaNYBpjy6TsmJgOha7I4RGnjOO3Mkx8S1WCjBZBu
YgXa3bpUWuL0MAC/wp6ou1J0JrA/Zo2mdxwAUQC2w3TD77tAuE2ak0N00sDUwjHfDVGhXJxQJgt7
N6EXYzxppwQ9TvS0wuOg2bX2RknhMsxi3xLd8hA+ehADF0T6eyKvrwjhUdDNhqnI9le4w1AFvxrL
RGaOMx4/D31igpCa2X60KqSQDMt6YkEbikw4VeqyHUlBAAnSvzbtuOz5idy15nE2HbgCmlF0l2Ky
nxfyehlhFZpIX+Vicft8eOoMBL5IsZvcAE5BsMIzHW5ea9WDipYfrngd/a+0g/guN/qCXwbzqItX
IYUbSFurOeMJWHuBeQ/T5OCRfwmkYtJDxojbvILNLP8Hha1YzFTzootx2JSBPUTSGyKewF27HNyo
8ZucntoinqkzhMXval/b3ZplK7K4c8dlW8tcwoTjWelLha4XLzOs3zoFzHC9VeELI55lqSTXMBXj
p98ZngPRIKAXBMss9t0n8LdIAtZrlRm9sk4XeFLZtdawSBoUgcr+3Z6tok596XieQ8YMG2AHmBNS
1H3UoqDqIDElBpcTaqBdL2HQt3uZ0vdhBTiLoJX+9vZNxVCZB/fqLpLWDE1C1l84pg8Km8Q8mfcG
d3RiRhst2SrNjF8vrp9iCFvIcBMhbnU9nck97KAfXtkd7+I/MKHzOI3UHaO2G3kU6tdh0W3Zj5cW
pMRHcn2e8TdI9Ty+kcPkxZAN4xf1jXKAeNI4X4nGJ5hYFKeGtgYFy7UBM/CYc6yjMNLedRMd8Cf2
6qSf/c+sTFk7pO/g+XQYwPL994MFGLpoRnTKPRO0DC2HJEV0CbHvV8ttiZXGQQIKthsqYAGH0as2
A4YYBUYB4pDPb+xndtDWSgqEAeYUldz7Fa7yYymCowhu8lcn0jm6B2w/dh8H0UUUdPwusAbQClc4
AAVvluoEzuP7yETtxbF+y2VtNMoIzj1nZ2WxYSmm34Zidj0zWHbCORM5wzEkkXmUPp3mXlBRVnyR
nsaW9ssSDDj75MGel0otsMRfqu1ngn8rnxp24UXvUENFYQFmDK+cms6dhH0IJ7MqGN3sgGujd4YN
out/FKc5uzvCCIlaAPv6yqFnLux2mE+sTJLB3KrebuInobe7Slkql8VC4nZnhRFGDDuT/N287lN7
zVm7DtdkraAOPJ6/WYZSoqYfKXJq/fAzNO0/I0uu71FaR8zH5Btf6JUbxi+VR6rsVi9do+0KzFR9
tzc/jqh5Z0dw4YUIs4T2vCWgpS4iO4vg1YQ527EgIJ4+Saitsi2UIoEpJIRvGM1p1/gfB314aXpn
tr2Jx05WiESuXj7bK+Xp0nyBKHLF2TIT5hugkXNHcSzJU+GjrEpUbn7NgiP5pYbNWVXdbfebGdSy
sjtmFqFjrpUBElWdTZePFZhz5RANrIjYjs5HS56nPKNpHwmLhVXpbrpJxDalKZayf0w+TqHpsPO+
PODVRg3vg+75OckyT+Z8Cn3mF2R2XjhfJNKTaOuCv3eX9vFlgtsfZsO3difPo8fonB6g/hpr13XJ
xx72hulttGWCQ3UwLZCeMs+4sWA8uKoQd4TIWZydne6fgpiX9G13u0jsEpMAij/fRYcbrl2vpmVd
cNzJWYxgn95bnd3uGYVxBEL8xwF6UQmuUgM628KN0s3zlNCobknxLpj9oN2s2QrYXZoDcN4WjkG6
QodGyHR50ZOoiKIZNOhRu1IZq5QrxwTiBw15An3i6ir5qLXOMW/NdkZCQ5inyG8IIxbWBZ/08JwR
YaGq+ZrYVLOQPRnwuU/0e8g4+SXqY+aPvsTEWNZcj08OZieznuvBmOU4gkVnSsXG4vXGOnsbQgTm
QIuSmY7KxwgHIaSVks335JpTbT96EJ8QBNJuNskhSMhqus436Zsy3mcBzPqqz3m8TI8w/Q5Z/ZZb
J5tclg0Z95IbZbeRAprW8xvI5aWBe3fUlqmbwMY/ffwvUqid3xEaseGdQpl2QaN6dxfRayHae9xv
scuG8FyIJlV78OoResOcSsCRd4O8XRzZwKdw8goBmW92vt9h4rjr8TgwdZWnWFHuQt3pTpUpssyG
d9yCSsae2NG5KwE+d8AIvfxAJcY/hs0tq3alILAY7vaYl4xf0mLmQnXgSkShvEYGcddbeT3CPKrP
vWVHvo25MvC2Kjy9srf8r9N1ooJcgDZzw9iJaUNdEIgSK+6CTiyPKTAPdRkCCbOJ2LLs/P+1XbHN
T9wLjXfONtGf55KlsGOP/5l7qPRl7S/If9tRo7DAyKlWG8nUf5lEuYgt3TMk2mE53VJkqrnpwFzt
NEdLPVsxvkyUvViemqV3sDZiqYoV6pmHEQRsC5mxI8Tj+p36o1poQgW04q+Tx5JeAkytsQOB8llr
NEml+5qDJGke1Vr3L7LMX8Gx/xgMgaQ/gelnbKGu8kTB5+0tHxlBwyqu7jlbuwWxk+vnUbuCRmeq
DjDWe5DY22Vgn+5HHU2CR0MGODU88jsQvzLYYN1JkREYsQj+aHFXUHdUvE15ycQZvN75ViG34uve
DRjzju4pSZ6ZSO46Bymk9dYTlm4Odl+S5fqgywhUb6s1IhXTF32E4I9hO459WtOETU0u7NVozvXV
Gu+W7W4b/IMhwM/R4IGES/114Bizk1geCER0aMpehk4HNwwOe6hZfRcB7cAOC8MeVXMHEwBGfSY0
8m8CCAksSbwwSaP6xi9jUuy65MsnEWj5EVKYUThFFU6jOb/M9iDtJzyfhHyZKx5NOPQgx0Ow4lBF
yeH1hrVSHiMdDsZ3hoCluEgXr4vwatrVi3u731a43peq0b9AvuZOEsW+mYTjRN1b31Z5weqwd9NK
upnSRLblJyeyTxkMu6Kz9m3MH58sZFoqq0V0f96glkX4ifClOtjOx+e8Ucv7vLww/O/w2ZJj9UUr
7vI8TWZ4RAr0GiAX2gzgjkFYnr+19zCiV0YWKN3j0QR86LcRwXp5PUj+Gd4MHFhIng3fJcel8p55
6n62DPrmQjj1UjVqjfx3bf38YNblQHHmIThPiXVY165i6GLcNnE4KYWMYFwakEMAq+nSzL7oxhZf
sMLaXZcktWZkH8cwU78AcaEaLIwxbFu8+iwZqZ+qFC2SuG74m9K1VL0O9kBp7jTUnyaWZXX/Q/Cy
gRNAmrpJ/2CEU/bC4vqXiwAcGgADGsSAsKnFwpj7mR8T9NIgxgUtZhbJSYBKXwgBKLPpK/GVW/MB
3HUS8SY9o90ek6X3rCVJaiJEPnz5SaptLci8YLXokt2Ca/b69mKZFpVzHciYukJI90zV4XobAXcg
onBrWVj9dKsmN0WfjtU7/iLubVuqelcX5C+TTxsKKFYwEP/5MVarSeygaSIZE4XLpIQAnm2Bmwzy
W/1vDwjm8BLBRaPCuXD71C/p1gXPDpzrUOLOn6LybWIZiL0y5Z1p7pKweQUHqeXX8KbeuiE2jAhI
UYTI5V9Vm08VvxH1y6OHMrDQWwKbw87ZAsy4J5T1efkC/8vt+OqQMQmE2YrNWi442zk95XAplFVA
RtkdgQMM6IUDNfH52++RkP23C5D+2YyVIHMRuYb5forAr9YAxkjfkUryFBjsLEBpAUTAbVS78H4a
5AfBlNifNKj9T1smKj1CF7HC/lxf0LDEMCixTSzOSA0yUYGFcMiVogclySdQ0zFi/zTm4deOz6aU
QdPy5EkQbZBccgAfkFQ8DF5aXTjPNQoLtGX0NAct0NfrcnKfSNk8PhWH/JYzzF8YL9BRC9A+jyNh
fuHM0lC4MmSYKvIK4cnsbVra3+X4mubMJ5JtTYu0+rRRdawDiL3NEe0Ho76jM55h/xoFtoRXa7M7
pqf7AHcjST42z6GmO/IMBegaw1KVYL8lIIVvsgrt79o+aLUBtmT2SQF3x0aG2v5hPp3VZT0o8MZT
diQECge8jOtReBFaZC6nbu2Io8k+xXEQsIckc45GCJqf92J13QVxxeSsUrCOIkjUgFRtpUixv1mg
NwVc63kHPL5/qzI5N/NN4o9k4Jgqhih3Hl+9evwR+dMSFfRfH4qSjtsZ3JyLQmvZVyhVKET//Oll
KytElIaQbvdlg8ndnOu4PjEw02lSOtH/l3j0t91HZZAIub0mpyTPu4t8GXa3qBVeFu5XQ8s3KdIi
UvKeFFF0mRZAivyUzk+FRZxRrIewAcgRvxebIIL11XxOS/mmrHKZfKjh3Y7arlx9mUP7pH2i8UXY
NbGxw5JubLepBvfCXE6DZiF3De3mfI+7EdmT8559/h01Ksr4DQN5YgVGhjgbAPaXXzc9I9muIYin
mnA2Gm6C9GpWI7R7qJ3//GSnq1vF+cZ9p9mp9yj5of1kIlTgKhYCXK542ckLF6gJyE0ABN1Jr/B3
9xIArIkHPBHgSw7MW63hzoQPCDUsoBHL09jAksb2bri6MBNsrCbktBDWcTkedCWLrVGxQc6nADCY
2E9IPB7V0Kr2FBmMCwHx/A5hpew7BxwyAu2yXZiebiVBM84Vkc12Wen8yN2N1JpIkmlTok63uYSu
CRsMUqFy8G9LUt+2hQTj21izm8iNzP11A7dYdEGCsD7TTpBn3iKr+5bvep6nItx1LH8pSuG2zB/I
y2gYdBowSBzmoHXQ2HkcmkKIqj+UvYljT5doXE58ekJNsgoyGqYBb84pFktYS+rAMK8ezFHMHasA
zodg2CHFz8IZIp1c8LRgZvr3bKeB4rqGPoDmCMFa4HKrErq9cYR7iSQk1S9di2GP+AbdUJh3Fq10
TaWCjuzq1T7X0stQqBmX3zSp1x4a8rUlmPQSHqljM9s1kiHP/WJxHTZj0OZNtqw7uZ1LoAwxOxo0
sFPhzciiNxbzedUSLvQZjbOo+ljbwb7zVvrPLmWSYqIA16K0p8ygqh2vfOKA+ldJrREjN1fGCFUJ
7gQjbg9zxNH6fjrHOogBa5Dz9LI9+AosOWPevnZasVn+Grcd8/VpUhSXrpXgUx7SGicFdiSezZlb
MxUF4jhMYSZSr1SKSplH4KZ18hmO3acrUEMUAvSN8rTAMiuaeZ3gYuPkHhEY8WkonewNl2dGAKqZ
3N1CPQYtkKbdR+zN9VnezcfdrIHc4CFSSLlBMat7mljA8YE+k3V+Kd9CrybzYKvyoSqTiRMp0LKh
P87nq9Oqg0gaBG9RC6A6nUp2Wom3w+8miQN4GKBNTAkOgNiF9k2xtKgqW2M7N7HPHi0rsUrsNRs9
yU1rlCyTspjWiXac4c23jC/8aNZuXZqYzxlVIryIfxgGgRHV5rbBeF6e3DdVceBjpLachjklA0ce
ktStX68CYIVof2T4ZMO0892cfbmaTgF2d5A6pS7QLoj02E/0hdXlxcQ3YaBcKYlyCYXCTC+OrRDo
0HS8eFOQTSh5Cln7Nhl028Xm0OEfU/xy3wFUKIXM9V9U/1+HXlblm3u0KiaNaZd4CgivXttOyzXj
gLV1KUazgOAupGEunvEs9Cjm0qJQoMcQSarSA0OMU3VszydBDDQJy+1NEuKioDnL6SG6FliXYs6y
Jcf9ut9H8EDVQTslMhZXnRM3KZVFrwNWI7sykePPq6bWXzJ8AWGvc/ce1zWZu+iw2nrbF8/U5D1a
SwiBIP4/to477FuJ87MZuOsck+ZxLpN9s+FmRStZvkebhsLOK2EKtEpxilL1ozaKcy8QvB9IEKbg
RJamfvBYZBlonHzXVz6kXxWj8mI9id1urkOaZKH2kSOB5mjhgZS3inXcGvgsfJicozekP5eN8c2z
z/puhiIMPxTXEYbcT/H/yXJhiPbKJ5bboBF6XXDy/kD/Z/w7CSl1i8c48sqXXoSz1ZcANG5gf2K5
+wamPFSTFnfahMmcC82Owr6IQhVMYxja2+UVTMz0adbou4klbdCvVzo3v1f4QIWLv/DozKpHM+WT
+xr93YtWTLmI0j4MxhyWY7IQxsl0VKPyZFoxcW84bVOnJE3HxAAniZElIyn0BOqG0j0mbKvWnRT5
ZeKzeBY0SuDKHxM0xq9EH606BrfFrJZuRgy9SodEjMWqV0GlgJBzJiMZKHm9dl6hc81dQwHv9Gih
7MI/wAxsaCjbjnrC3Kb8mdPI6AxeMoVgk96NYdAb3q9E0B8vfL1Jx4MVAEvGvVh7XorRQo9fVsPf
iZU6CkxS24vTyHRGfHvW2qUZ0g4714o5s4UulYhy1OKfNNDCXVw0EZaYEvXCESTn/4dvIfndYUXu
+cxkCfiN7Psi8sc6y4VGbAjEI4A7KTu4wGDkuo6GjjhhN9L225czFBjes85exTRUKXsd7yFDrQI+
c314K8h3rncA0v+SgC9eIoruqphC8tiTngiCeJJ/Mji0OSonscmBIa23wENTPsD9WmjTFnTC+BLs
kZUivE2caeSicvlLFhnQPYd7jl3plBuA9y42/pIcQ/P8AWqRFQW+qVjo3DpX4viPkFJzRQ6eSJhK
9ANEMI401k2pNYAun3/lyeiMCkhnFZqz0hyV+RygSiBtMJPOXpD/Eosi4V0QmkHskCfz1DX5GY+n
GNWuHDRy13VWbL8vPLeatC9F1zf27pcaLlP2N5WegKHZOAypcezmOd2U73k3PleqyWjrcAca1cJu
mZrPmfHZCUrMrPYPhmjWyF53tUDGXjUSfCbHZRAM64/mwDaF6wMK4c7CHT945i4vHgw/UBcrRAfo
pHzvK3mM66B/Rp9hOmQkjGiipEkqsDt/RDJydXAd2FaZ3Zph72q7f8f0VY+OPbOVOmrWkSd8kGi1
hldaLeBqoYjqETM+Kaab9Z11IWAK2t413UZ43trJiv6ybPANqdhWIWKvSzW3leHZS55gDzCYqMtW
k3XJvezbUl7MFux4GdZjP/kNuL9Z9/Uj6sUbXyCYOpzIl1ZjQx+4OIDmkR2V6JTVBdCg/3TiezrZ
BhL9m+j//UxfZ4/Y0TjnrP1HY5C5lWlM4Q00YQdsr46q9ALl9yePke6CERe4D6GiWGh7YjcYe/Uy
IrcZnxZuhKyjA1u/Jh/Cu9LL+NVlD5N3RIq9/r3i18pPBWcSOikH90Gf5VT0u2a7lDyirszHffQo
odmYUIKiEAKmEBRDsjztNJIUJMi3emT+CG79UhstBgj3+rUQ7zmd4M4D1ojqzR4UnWnb2ZPGhCIf
76fG2DtjLUzg3siLw+FVlbylUxAV8SvtLBKdlfOKaqMvVZI7/4GTJWWUMxhuuIZEbmfL45fsfCfU
7MkYuxwVLmjXqwRcYdOLLxlCB0r5srRnPj1CEnNByn1OMTOtAMC4HRfCxgQVVZSXW365fs7Gd/Ak
pnAEB++QlbV4XWFiv9J8uVV3Dw7ci2NNII4fUwxDN3jUTdzKJxQuPD0bJ65AeI6Go/J53J/dTzqD
bNaEmgNsrgrLKu0a5tvSb4pWuLi9NUAx9PcrM3lwPLC0+VheC9IfUlZkaoWS2x7GTeBUWZANu2z3
imyRpHPBs9MVeMRkxtRn9Ks1CxJDItu1jetg0mA6oGaNccw147TdnXpCpmCphcFjsh1EAHjbLpSO
IWuHmacwfXfRSjA2Ge0D6ou+dzgGJfrjD3nSSls9mfOEJTPxMvq2Kixy7GWNJIoHKgCM8CmQNUdy
iR3GmRCnhS/CY006uNDZRzqjXLanFibMnM/HytCFADhElz/J7xClT1kw1+mV29vHmYxQOw1PNysy
hZhnkc0HhTZOkUO9NMCxtvfVy1la1YRF4EVAlAgF9SvFsoVD4PaUx6YAe/6FnDm/JN3OpBqdoJJV
g80xHoCPAMQWXShvlNwhXU6Un+RV9MG2Als9UGw14CuRz7UG/FMq6lSZgEvsMIl2r8Kj+sjusOzy
EPnJWJZJJ7xu0noWg1HTAC9p8RGiU7vSCK7HJZIJPtnxEh3K7H/MZSGrEo0osM+2OaxwDpV2Y52y
BByjzGX+DAQ1IAqQnZqcO540mtyxSiCI2sTAJLvV39KA9/DYxSkl7hYmNP3YgvmyWjkEw1hssQqO
QNCV7d6QiWJbz9UcFkcigyaY4x4RxGLdXHWe54T+l08h2KLCwl540G1DHVtDUqCp1+hd9uQa70/8
696Tb9Zr1VY2X93CSluOp9l3ePcsMvB9Et7DIX+xrvms5WdR4Xbl7RiKwtPbQtnFib7/wHgQecjf
3BPsGj2+E8N5M8RfseT7+3do+J++xmCj0zkTLAuaDDQwCMutU59SuAmmdFXXN1OxFPeV1kuoIihY
Lq0CpRRojIqH1MzBa92aAqN/O71OeoC+Zgifnd5vsm67W6cb7Vqr50/Lvab9CoS+qhgMmdqI+KUh
j17WO8wKUzBtSYDtByKw7lKUB7qo+ui1uqCivjeRJgsNN1oJD2nejjPzOTCGF9F0to1Kp6YQ/nfb
467Yo0s8Popf+VILjahIkE2U9jNR5rjkj5QHA5bpfDR76VfrQDZMo3/QuARR3IUacvcYk9l+OIIQ
SRVbQdJfJ70j6lxaqtXy7Keqgtn1NQQHGHTY77eBREAoyeTOHe988GN7ur4P2xFFJJrt/zZ789ZO
nJscUzOqLYwxX13MenO7wTl+xOmkvQSNZU5w9MMmw9Pk3Z8oOqoHzfjW1Hc6exaEgYxo/xmCKkvA
/OQBN6Bo+UP7lPjFiRLg5Nxi3vNWOO4e6uScK/NK3n04kK2zgdYJ7jj1t3ebJM7SSYiNslPX8nNn
BmlnFbaxYt0j+MviFTpdQ/aTCSS3zCyHh2HIYgIyXBEfe90+wKGdfrNP0YHYFAACvVpkGlnGbYCy
geV+uaBU5O05O5arKW365jzm/Pmn5u52dgn2zIwK51duQ94V1oTj6CR3n7kD6Z+0G8DMqJ+UcHog
PyginkBvrJBppKOstlicPBiwMRFp2XsPUdE2OKvte9HE2A+3AYytbnFibVzfXT8shwAYJ6/JV7fG
abDpmjIkk8jY6YohsFF+GDbYwBE8JfA/qNmghdbGTHrEwLGBIGrBKh7/rSJRLb2K4fN9KaQFvhIz
waivPFX6xNpehlrlkhGtTz487P0XpW31QS4WKudMFL62bdRsyFCektgGUEQKw8rzmQIrrGPOVYD6
qmmKhd21EpHeYTnl7AG99QA2sX1onh8hX59wqFqUosMoWGP1Vne6WYoJnl/73fUFlUNldsgkuKSQ
1/bYCDQSK5/eNjBYCAZK/W1RS1+loxD8tj3P8SKgPhwkJsAICnBRyLOqbGBkBEIMWXSJoasUE7C5
KKQXqUyGClZphFLZVLwY+u15977bM1B6j6eDTRIfB8vStb2vhSX7TzSaYiwYitmFxH0Fo7KKfk2H
u1mCF1fZM301QvMbQPXrP7LTwUU7W249lwpjQCwcLW/fqJZbdstKXUmo5Sa+FuJXOMynMX6DJAwH
QheI+cscGzXxcF8/ogDexmWA31adK3mtuThGwwsbk2fVjpQRI4d3663SN/Tn3QykUwTal/8C5esa
Wn0QlZoCJOTBe0GFEFyR1vpfooCo39to+tU/MN3n7N9HuLnuHRBWVGfowSNi6TcFfaX7MhuhouGA
kW/FdQRHUib8KjpuGek7o7AXsODGwPl5OSi+NsQYorupkAyDKTl+H5+j4NieXmD7qZAfYKmOkRD9
NVuI97DXbNy/LR1wANXRJXrWUVET6IrH9OveM0GthSQx97WFsBaXaGFhqgaTsXwGPKOu5hL7q1Kv
a+ZDoB3rR/ArYRKuk55r2KsdJgLnKyJX+a+lna0gZm8Y/8Ot1M6V8Fh23k/vBOVcSvgcHf096SQe
vnOAWz8bAIcTZJGUUJ7EzKKqWtFLpFxFtCjWJt7evohFg2bLP7eyMkT1dlD+pQCacAp5BRtmGiZv
Z0ePlksaQ7XwnJRXpqTkIAx3rHlt9rFmMoh9WCmwxJfQQqycuMBBUQp0VeB6yjelU6l9zRaCWeq9
V+Ospbh+WuRTOCWE6SJ/rcNkQQe78sDWwIeJxlPeVUSfPScs2ZnXiXZZZ6lKB//LCJWzUhw2h65O
k2yyW3EQeK3kUf3f4NR4m7W8/6lq3Eu34xlaFIHnp7sEA0Ga+QIWqW8F9B+AdGwsx2up5cbZBY5E
rQlnW85teIxsdErph0kbBEV6b0+jssr+/uvI51DTgKuL3yfngUCnscfcSG9RuB5B6RiFYDvpcQNZ
vnwmylrVo/DriMJiWEZkX5HibOcLwZoA44vnOXw6RjYaX3xwJF8VewvmY+vezZRpgqMHM21mW6PO
su8NLaek0EbnZt7H4v1j+OQlPQCyAdBun/6t5n9E05/RwwoHVqUYJ7XnCnVUa9k3Q9pClAYdrJ2x
G9qyita81Fn5h79G5Tkece23rcfhWkSSy1zORzHolMT+Em3b+AUTH/WWB8r3c3HfxigqliGT7eeY
l9DPvIW5o7Z7fXo8fiFncdnpJf9ughDTG6sIHLhs1PfyJ09XB6zZZHzeZb+XyXkAvFL5pKi8SvEw
DjSuzUJRudznfvpO/w72LB34k5DFGfD1rF0WV44bjJQucl6jPVZkWYrB6rZVY49zto2nHEjfnlpC
Q6vQRJCicGISuckgPz97242zt2EM8PYuvTVqzZldtuu29H1288I5N3db6V135gHaApkI1ZxjqYdJ
AlPGRJnFkb/ZEgts1w+zkasJ7IrV4iW+B7RjQosuSgOG9ohKSXJl4irel2SOTkuAsQTfRyXoviqO
8UqFHzYF8OA3i8w+3EX+QRPzbWjJUAYQ51OMbKtDdQvRKR9xbuYmEYpVndKzFTSgcFNQCweioAPN
EJ0ZjV1XMpVrD9Jc8LMcFQJoP2mqaj6qzlzWiPisHbGHOnPkBKl6gNctN/C0p3Cys7XRo1O+mry6
h0C8KmKiemRRxmvQK/ixCSDQGtBuIcGIIFOfNQqY7WBdukHySK/HRupBkmjxqKFPipMu8RdhoDv2
0WQtjIX5+eKVq6MQnaO0RCNPK15tWRNths5hgBpnOz3I9tBtaS8jfmtUmm6zzxHVc6Xkaj0gDOGI
t85yF7DrFMNN5MYADx1YkqQhhGd4TTSkpoPz4FTOCpUiWGO0wQlOEhac1gRZePR54keq8d4CvyiY
S4hd8nAij/TUxn9uq8fiD6Lv+8E3XveGFBLWo9PkhBfFqDoT84ErOpQU9Bncs14SIweokkiEUJcp
knWb5sO22JFyX4sYeg8iurIpROJTuABq81LIPrQF/NKFrKdWxErct7fZdCnZ91X9tqyVF3MMh+8v
g7FyBNRMQ5wyXURA5YthN62f3oYA75XB14fjAMt1HeR9fN/kUziA6sQE/RG7QnkSOeCGusRZp3Kq
TQ+yd7libLCxvQI1qFpsTqjb6NuNrk33l46TaIAgo/c9wbq6VZR50UmWOQfxNab34y30gUvgNszQ
+ewU0KwelYjtaeVaXIvGUCipY8/ok0fHJdTZQ+0o9ItMOTPIZ6hik4bUjZ9i/I0jhCknqSAROpAV
OuGQmn5g+hu3cAYHwXtaK0Rr0+O3y90THeqy/V+8OxbboLPg7WYbS/AyuWFrAOv7cv9xOGqbew7J
2DgN9aYGtPXIdsShJvLfEdoP1t9Qbseslh0H3fvRIvLnVcohLiUo1v6ZloL0p5M3eEy+woL2iLrd
63LFqlQqOXBCDLn6PQU3eUHiZi/9LvzoHeposf8AqZEvR29CTR5IM8KQ1vFK62fUpmE6fVlLCtCR
eLAtv/KiFXRJy5eXqyGlBG+ad07fFTcBatyOUqaOs1SimaEV8B3ooNqm95i4+W3WwxPtB5EEi5Tq
YIwJ98i85e4df4uYRqGMsw3i5A/+lxe7QohWjs3zqBaOFksv39H/FMR9iUcGydsH19mIbpRUTAT0
6pN951e9HLLd/vLpza4kll+YEkEyRw1ntzwLdo61L1ScY+AfOo35RLXw3M19QX0fJzZLrwkHbF3P
emc52aTZ4gWgsEPf5nyal6RD3TLA3t/TVjeONI7ekiqsSTER2BOgcMiT91LRVrP7Jvh5KAR1KACF
obvbNg+PYe988b6Vpt2OXtm6wUVdWTMAA2CQmWNCOUKkY9bGCG3uiDDpW4kGnf+Ey9+3m+hppoCo
Rp9nb6gyd/5Zl+QraJgMO3V3NPm8hfOTYZ4RrLRgJdGNG1Ci469FSbQBLcY18JeccYsTiMPs9VQj
vDvQh1R8PhurMVC/JHdQ9vxmf687dUdchRrl4HHjOZH2qzCq828EKqc/Xt4l4Nm0aedPDe0kmkve
FWwQr5nv+rlec0UAEjo/68wbjt2qgGkRb9KpI39e992f77fW6w72Irt+jiYcGQta0V87YMZCOF8Q
bv/uNHlrUi1f0Znjsdmy0siqKMfATx4gVQJr0YwU4Nl11HqgdTSy1AhN1BRJ8729z3z3RGhc/P1t
z1pLttXRpuJQQ+kQ8Xv8J1Qwio0xTx9QYUimMnElSE/xo/bEcatAYuxs/V7lOQfOqFkd+az3wUyo
J5RzPrO1fRQJTNRZ75TPSHzYfzna21HAZdMd8JclO5rOcDm6fgsCpmlasy1nxO2+1li5zBmXeth4
YdPNe+LzFeltEliWhC7OH3n5Cirz5aVpOWcc9jHsf7STBgh/4Os5Chaf1JeFXe8X3pTgJhvU/78Z
2o7cstpkvCV3uJTPqpyPC8QJNfWfUft2DmtulW+qlt9SnMOtoupwP3Wqka22qFWTxxgc+5Rh9all
bj2OmSe7n2leUkR9C+9YR7CFGTpbqBRp643lRsNdR09YfMmK7iKi91teTXlJiwBh77RmqXPLJ0sR
5SfoEi++Ht8oc2rRDhshkuHeYEU1sibJXqs24rmLmW2dW3Mayb6hf4jMexmYDGvArbD3Zk9rtgub
fduiIkWDWnQIREvDirEVxybmLlbpDgGW97qIgXlDXVGruMhK1nI3ck4i1pRRSAiLBN9sCWL6Yhaf
fBHsDF8AKEBzXKvbGb8cwxnxa715UXEJigyu7mVeVdvEc4d171HxdZElVPfGxyuO20bx3RzXPXzz
NUS8pDA9ZYTu6eUYfBibINGvacClRXY1kb1lnBvpIdrqLCHruZvoiLHUHvbfgVyEIh6YlW/W3NbF
Ekbm5BsraAY1T5mS/5OXB+P1X+NorOhTQV8uEDBZ6Yt/fsRcKnpOloucZITLxexOiEyWeGYLL/QS
J+HXkkBQdpxRo5PwyBtoo0dD0gg4yQHACZ3+7uP92mAgYNLL1E6BhqKIRPKL4ANVoPAgFLiTbeYu
X98/ZcBGypigbixA4vTNT6hhxuPS8ne0FVemhVBmugL605AaEznPuhOcKT5ORPQRhKBBJDN3/aXg
A1IoF2W7+e2OaEkPzzPYDsdarSpPxNG+OSu1k1AeE/GUxVicmpW3/eni5gtHrTrNW1uDt73oUJ5O
hi0+NwiiePvoPemtfUtcDVaFqiPIqJOXK/bCjaJfzNZLFcvViltuS3cXczFlC8LV0l5FDED7bWuj
TUb5Svv4k9sHVjeH3/dlBqjgy1Yj+tLDCBGHh523W/JGawPFAixCSttTXsu4rfVX86qaR9M7hfs9
SN857VinTG3DZYX704vK8wtujM782/tTqKtpAy+FmadOGdSe56RzT7ykN+JF+ygXt1G2qMxehRkJ
EWt5hIl1qF0+cEMZ3u4tc4i2A6ToePz4J0SpbJh93d4QBxaB+V+9iKjOUvRww1+oyTmI5PPzrxzX
XH3WNQl8CRtf33NNeGswp5yv00ohtGNi7+2/CkZ0NYhCMEm9gur2LzDEyVzgyMCXklRIXHAp+Wzn
QeELKa07WOPDeb5SWJ6shx9hC7EszbHz9iOq8J3B5izSoGcJtgmUnpQPFacUvQ1/u8pYwtZp7gOo
XcjJVFBmkZAHajyQihBFQy4fcIB+GnyJM26WV2wrraxR3dY3b7qxlzvPX9pLM1JJ8pA3eowGyNzF
1TFEonUekfqvEGSfd6t3r8aNfj513aNNKb+wCTXTdM3kFJjkSZOoSreyPypX69dGlKtMP96q5Vwz
A0MpEHwhQ2bfZ4FudrK4NHmlrCgc4ijZ0ouPOZ7rFWm3kRfHpp+oTuJ6P881kciJXEyGeDMwinw+
6eEZhpak+8xYH+dcyKWKpCL89z0hCTVAVUXNvsB/X8xUT+OdjMWJko3SS0BNqNidLs4UeEVA5vrx
UAmrdq/D4sX6gxpq808gLpldUGSojvmDkCN/tE88t0/iLpkWuN9ocuJPjbg9r3zUeq+a0EoxTZkn
zGMx0JKcLfNMnf4vLG6lcf2k9iejM045KIik4y2VmT1ZbSU31ucsLlujGs5H3g4OJIehLroQrnJ/
178L1wc6DJTTSc9lW3Ng53y7HtB/dqSVgx8ag1N1XiChCU1SnMWrLXlye1dt/dslU09JEWPefkby
W26jROEczU0IKS/gCmFWeKk0FSC4Mykulh69Ixor4t1TLIxWkbIsDqWYol7Vw+pEYY1KD4Egj0KQ
tE18iwFKSNy30dyZa9ZGGcLHP+5g1VUDM1J0/mHTBF942inBBA0wtz+0ZlvcINtDD0iBDhVk3ep7
MZ58NWdC8Wp7ChOmWX+vMfUycFi7qF1fssU5eK7AHpjWofVwVt7B/Wh6iy8oESRkZK+PQ3sOFqJ9
FYSUxnjLo9RrzKBK5PnT1nXfh40/VTtCSVF1e2UsSEuUUb47V+c7pXo3ZL73lVPlZoC4nxahTznF
7T2wZVzxdn/1hyzXQ0OIT97P9xIOYgA3qnTnJkVivZjGqSk+EfGZ/clISbQ+yCdkpeD1a6K/0EL6
q6Qxw4r5N+FuydbtM8n1/DFO9hLPzNdxx2QEZ3atqFMQaoq9dNxzOmbFd0OcCjfNqq0B0wKVHeIS
u2IqppnHm5pYwUkYjbOJmprIlzy3ET5dgLUmqa90fa20gA+lbSnjH4c3Sx7EPSQuK1iDzuFWxzvJ
m5j6oQUYqi2hnjB/VScJ70nNcAzybLXhPQZzV2qS3U9qMJsCjLj77LdG1JXvo71oqQua43/mSWqF
4nUEN9+QofZa+vNpa2MkElFlOkJCmeoBU+VadQII/RAulPasndKpGvxBuFSupSDP4UzVOXZmy9+l
j7cT+ANLnWMtbl4JQaH2sb1Rb7+ITSZ5y23Ob7NAhquJqIvUgeeFSZkRvFq9OURN23WeHCymnQPn
j/aFmqNG7ih8ugXTt360DLwJHeijpZtT4TxTdLEwETbriXUEFn40h83NW07Kje7zqz2EKJs6YTzi
TCbkEK0PsFMs4hH6jQ5deouKQm8OFHT8ugg2ce8eRZKuPqyh9moHNK3W+rwIVkdjHFT+JsmzFlOl
fOfGKVMxOGbP9YHXd1WHU02pqTc+wUXGmSoSzkNypu0gWHWW+gZuLhOdFBy5zOch2303SLM79jqv
6CNL9hpNmo4tyf5sFPfSd6VOIqSzLKqMqP0iftIwASpxYKYmhitx5VjT2mlmLTjx+AvAQWnNavzY
UuZfsXVyFP4v6KaL0uSqn700FBgIcbpb+fnss1RrV8bEOu6A3H6+ac/3eWzo44vUP2J84RKglIHG
rMzinYMbd2MaaMAYAxQ8slDNUHGBtsYkyGRscAbsJN1E0mc48vt/x5YyCvzd6NB2QMHlMMNxaWQZ
uzcXv0KXeXcVnQThizc2DkBDfr39tSnQ8gMnHE3HU/VDfGFE5xgJzlv2CyKQ8ByqGrlFdz01sv7F
Qlcb4Dos3x14xj2cGBnziPEtJT6Il2Cy2RL0iKj1g3HG/oNhqGycAjlFbrqftaa7jRAFG3ejQGtP
j6PwHGxBIxhzFFCH7k3gLE1ueXlbXCtY5y2phqmWHDt2ii/uL2ypFaVW4yZ4fCGWNdariBn0gtzM
DTjqLU8x0u0bM/M2NRbb1iyLGtNNd4l0E32Z41UlgD09KLBybeYf/QNVgCqhZkpWJMa0JQ74sQby
84owk6HcfYRATZyMEUgKZ1MY8dOyiZFQBlh04aDs77WIogVxgnLs2UkAWdlalRKwSGxxYHkZJqmn
YiD9i/RUKGHy4i9rJuBjAb04pO9/DW2n+/nQaiqMq2BYFx/DoUq1gbdEMMihsKemZAwhD8HBOgk3
Y+LXGqJEnyztH2sYVoRFkT029cDoYKpn/rm0ph0bvl1ptZlSYSK2BU8+faSi5NUYvQ7ylQS+w3jH
iSMqUXuk0NCfiIkvm5HI1MKOKmKGESZgp2uq2z1bjl7NlA48WxwIJ5MYKwggi7FspVZQbO6soeG1
ZfnXmk/cIKt5BbkkM5hxbM7GOlV4Ohyh2wNttpeXncQQ/1YPPdLhWsjJr2dYViqnwIXZRPA9YiIm
u7DJBhaeua30MU4k90cNpxzbuvNwJTAsd+QvoPMrhRTWYHhDRpyeFn+7GdtRZUOVRf3bCiaJnY5v
RhCLTn3xj58IoMujCEJD/C8tcSPhd2TpPVYHAsbqAW0XR7HB4M4QU31y97RNYEHv34NwKBiHmD3M
xrmH0QuhoNJ/3mE/FDCGqksVqB5w9NfRbsIlBItqEMhLHqzK5xDd9UiteXGijcRTb4TS5cn2acz2
OQZ5rHLSMw42PJ5+Uz/NL2D57KgLmj2I++8o2ut92QEIvj1D6FtaiDMale4NVGxj3xOVudpbJUYf
okXM+W3bCySy+M5CE6qeWIFMMklUoPEuju871k7CMZwv1YedSQvm3aazUsJSR8ZvTsyIZwNec6XY
Pk18yo5vssMza0DGXQ6Hlwt6gi8aiQbdCQI831dmj3TLBDCw7BY3VGPoq1ubN8as9jcFDJC2TRrJ
dvN/0PY4dKLVzW36Os7el3+1YziefrHqb7GyjtsoARL7zj4rQpEpaPIbkwdkAtTYG3yAqz11uuzi
Awnp1037pkLWIWRMw1hmAPUd4iWAeluaA+2KkEhMWpTVMYeuAWpOnQfrVxr2xhvfEqfm2TNpkF4q
juejAxV2qkPC5VY7TfIJs/I48hc0m4eicsMM4VS0pHRxGKnlrgVwVdt/7C1I/MoTUSJ1stE/5Ati
c38HDhmysr6LRL4Ko1FFUsChqr2iNp5W4B9PnEcVQRtyLTj9XomPwMlphtIHZosXfd6W+8wrjtzQ
MClw6FjDUyuakyYj9OwHf0NXe8Q3RmOS8L211w23SPDGojp2U54qLdcbSYZRIfXbNgLDySYCTvqy
0oQFFh/r4K3wADS1rN/6cES21H0WljRmaUOieqevdko8bvyyoH4dA4MTAHK84h6V53VnGR5MfZKw
SbMo5YbuGzjrFoQG14gsEZFk9OoP7RoAbPl2g2YH1gGX5eYrrWmU1Zv1Gbu3I+l3uqUSWUsza4th
xkC5JFd1ngZT2yLBzj5xcANkmPEtoQbNbqL4noJ/T9H/PmGHELcSKeqx17TM75nRMF9X+uyKk3tz
Q7xQGB0cA1Gpek6IUWAINZ45x17ApeEfAiNDfvaS77fvzvIDVcq5hMGfBucVk0wt2jNJM6lDVE3M
D6XtD9qpaA1WB8IhQ944D/7H445USBoTijyD12GmIIVi/nUdGdv46BweXmI14FnWPglXqQQ/bvzp
d+qsdjPzeYRH4Ax9WqXS78NAwP1rSE42G1Z4+lhHrqPO+ImaqSC4Hl8rNW6JopewAhrToTYDVTiK
iHLVgnzpSOmyZuh4rkBTVEbqzlojeIjac6z+xRdY1uAsVuolWgnEnCM/IXX0JZ3vRS2A3B57lE9E
ncICXyMCFLCduxdeo8abo4BYxQLkpwH11N1lF3+W/2ZG+Q7eUQTV8P8cdHgRwGFhzvrrhKjtxb/9
j6wYWJGtKGPBaUFdzy5xZxRvqg2Swzgj/hR2U3dChiYIbxFA2QpPErJ9jzH/DBvmzM5RTpeq9M6Z
ma2zVvPypYklkCGUWuDVelh0kGCjIp7iRsuyNt3eWSEHmP3PZodyb5jtYXZDP85LAWaJqPaqtFBb
38c4Xdf7y1pYSWe71+uij8lPhMklk9keSiIuiu+rTmi78rrV7LyxV5hC0vQxscGncBjHX1OdRwxf
aX1YgmE9VCmFmtdww/CFNtqvXtB4O9P4GYZ7gjyXPzaTS9gOKf6jxmnXtcpt5HB6Lfvx092yf9YR
KFJs6ce8m8u8AuN35IgL+g80yObtYkvIVMpCa51Z/Ikv0HrUq0PY5XleBT+rRhW120JSFnOR8Glx
ePXPa8knq+5OxGzLy14pAo0zXS9g1NNL22W59Chh8J/WYnDLzkJ9dMYL/dSDgU65px2dJhTGExaF
j+vRVpmDMrD+A/60JAlu56gQ+hJKsDKxIXW/dBZ8grpDXHlQbTmo/jWTlm4aZ4CAKoVvDv4LgjBj
i7T3P8s5wfL1Zs9YbyI1EXApM0aBIDDutcFjQ/19gwVLix8xWZPqZTTU74B02YhT6BH5lnUrrpX6
YFX8yiitjroC5dUw3AWR6xLbcfz3cMOq57kSfzvVA6NCIOvLo87QbXtphmd3EmA6P3pN39YiLHqi
mLkSRwf+ufqVQEFPDj8AUs69FLwvysMZ3Ljp4jeX+AJoFgYBoX1cxQIjlyN+UeFxvCDVYp5Gt0JC
GFeSsflz4WH9aObmjQySN9Lyy/eTl9BBBQ3q9vSM8BCgIvO0wpORJrgblxfBMVPXqp00EkD0YDdy
m0oqCK8Jjcqmk63IOUTAbjU2qYO8mwjcEKSmN/2s1pay+O6xdTQEBIXoO0pZxLH3EuIXzt3fRCID
Itr8O0iokZJLco5x/goAHxjeSLoIfvmE/+vUo0vEKgwKNe0UeijGd4NNebgHKp4ThE/81UL8GHSt
UVOQjo8W1xWDbUc0eLZC1PmQxPgBR3Z1+aXmsCsNjLIsBcUZrgH2P4n+sFkxUcJq1W2XtJ1rROTz
bNHlb1MU9BfXZRWSmelLexg9c1ulvv2p5a7kDgOSIEBf/Bpxi2Mq6EiUFEkioplQ0S4avqrWm6aK
9x6m9aXRnvWV3AIIwpcD5YSSncUFTWL7m63pY3QvwS4BVK+RP02664ePmCuxKxfJ59x4i9QuXgPy
rqIxZsYNmdDFyOcmUh6WfTmKQ1AqR7Pr+9eBRgPqfMEB2d4X6bHNOL1gAoGaNSIhfdXO9yUkJBJK
ZO3h52iEtuyQGgA8zLKucsBsRW1BMZvc02/8W1reBIG0CHZp83ZQ45CwUbVj0XweLmySK2ID71N+
WIxMoEEp3d2nJhWy9VS5gZGTBE7YDcRNbBDUfN+0h4X9ZhG65c0yiSRFUzVYv1mVyCSDzLOeKgKP
PJ7ShAg8eoAUx1X6HoEcJOXuueMO8dJlQJjEpfVilVYQKEIVZ/l1iba0rwA/jGLcLUnuY3+kXKAm
1r4p5Q+9sKKxC6Xi/NzWdPdfWY8AF5ovJ9/I6TxtHOC5soegO7DLOQqiypMnTaPikqSgxt3lJg2K
svB57c0+rE03EIFEoR2HFev1mpoJg2SGkw6yXdWcEO+PjJgAEkSm5W3u8OUKICfuztlroCZKpz54
CZq5LVCwHt7A59HxypQIgudU2KLoS0kozoZIf+DCnU1WAINJ39Fk/eGkizkEQ5+3+5vC67QJdpbd
NEF1TgOLzwxM5EmopqGe+UbFOxVR30E2ZaF2MYEckhxTw9noE4Xq+hlE7mY1yOPjBI8Z/OhcDkSw
x8wcUyVnE1UW2k7DB0/F6W2pIqNDAMZcE4FLOEzCoDafO6uMwIp7IkWC5et/5XN1BzSzUsrH5S4K
aD2p5NPRA7V9swSVrwHekt2sQ/7PpTZp4mT1OayE7WKWmvfdoYoLwf6O2x8A35E1FEMnOLDz2hlv
CtgY2HUpstzBEUQtQKgrZLOma6WHfpLl5+hSd00maDJehpr5zWd3r2y6vSAQn1OZJFXU6oK5gUaZ
rUIvnhzBtyy3BqvOOS+SbIKaFL6IffhTf+lc4kJert0UfGwHvAAMEtaEinv431C+0nQ9qVfLQwO7
G5svuN8L1xkHSm6ngydRWuBAZxJDeKOC6e5/KqCbxZXz+SJ51gx39Z78B6mADL5VkSGtuIQWimPq
5l7k/eigJZPQNmFXouJPnTEF5KOsI4OWZ5zB1txn3EmAyN4K1Ywuucm2TT6VB3m3LJbP4xK5mgaX
C5d6XyfWwmk7jmHuez22m7PO00VO6dfdlnv0tp5dyi21FtiEyCzW0lgxhARBbWFwpvUy7nWXjbXH
UpOJYnpNHIujCv5E+Zy20l73Yh5eQSgHpo6p3P9Ha88QQZmNT52lRHBRBm58T8qIhN/MypScxTHx
as/tAiWv4/Py2ab6yigrIFLuXyjCdxInQ+E9dtFSzyNSO33aDyL4KDMCuoRmborxQpXQV8VfchXL
HIl1UsjIeaQzlEw3GORyArwbsM4Ki6aFIqlnlai1uNjUl0GK4V6lNA8px02j6eEzZ6SzFfMT65oO
Os4OF590d0Tj3UOCBGAxc34hac2H2f3pLbA+l/Oaa1b0PRAeGPAWNPY8XadKpoBjPJ1P8IwsA38U
+iImaG3pvXUCLkOpM7CBKGwrjQdDZvAV3hWndj0SbQSSO0gwtA6DccSMNkZgymVPkY4TTY/yRKnS
TJDHmm+l5+jCgEugVTtasMAZIJIC44uiMO2aToDZ1g2sHcZPo34Nkl9ZEIAIwB+aJnKVWOwQB3sA
qe1pkG2RVXy7W9F3ER+PNsS6zsGfrgL5bp+dNp7FPXRT2lVij9bliW7kOeWgQjWm0WG5ZQTJrzx9
uXd19vyS7T50AK6jATZYxnEPR8G64MCEOjM0tqN4fOC//cApJSCrPcVzEocUBzQaMzwT42WRlnAH
agaITitsvKoVKV2qVRKKbgMVSlWa5lW7vlsEhk9fnVzUX3k8ynljscAGilvQB6CGI3/QbzFIAJRR
lhQnutGeYHHHPS5I/jQOoBfGTZojXSBJ5zgIQsm1O1uAF97k4WEg/BM4BzKwkA3SQbfFzDmmBE6d
VSVz2clixEFiMu6QD6itwxWW7gOuXEQjwQar3lC9PplQW7ykEuxWibxaZ97imodZW6OT1Pn13Zho
IK0Fef4svxPx0d6o5iKEWMpL/f/JGHbIRcwVHFgs4UD73Dn5wXXzCMsyXX875rWUh9J6UdlAswLv
4rdTSg+GohSpzLESwsajBJ1hXRVPffZ/CeiP4CEpA6K3v4D7lUkpZxTHmNFM2WkkBg2hdVavTw8e
rhWaZjnki0+CreJSblvl5ekF46RGplk67Vg3+0+guDD/AMDsngHVdyiGBGFpd8TO/ASEyqttQI/z
Kz9KhT4XvUzA6QaOLWUkps3jhcEQpzfVXp5e4VpqqXghtUWgN0u/BLB+bACTeRsuSE3BE6Vo6/2W
ubXCxGoLrCnYdmVnYwcifjNPGpqIPf7tmODap5B1wM65Jg6IyqTiziyXF0uqs9WELUwM706noQZx
jOujAR87iLCMoAkIW3hZyoCGae0vvrvnsPetu0S0E4J08zQaYMEVzdcwsQxOoX/aotOVdQ81/hww
9pemgB3Pt+vQBbf3/558eUFzUA6Zt0HuwW8ncEHGZPo9QvSFwZVl2G9KsEt6VMyldkzZ5TlfheOX
wDghj0vqK8/qzCl2MW+1jvhRg5NZ4OBW8roKC9N6qqkvHN0mSIIgVjXoaW8bM0j0UPX/zu3Ggqt0
0jOkHprrC4nHOJ9gKtBbaCgtsVJuPuceqvnalJrh3L6pJfk2p1DmDR4A4YuB1AslqmJ7h/ucnxAf
CI/EJV8bvBNH8Uii/pmyFnMIKr3tKziVD7qp2y+ogVlhXGOn0hQWrSEAULJ4T+iXijGm8XSILKpf
YCPVw1smjHoaadx8tOm6zPfQr/hXIM/PydtOCNeqxD5ImFLefXhwhdKxwT5b3irgfPz0ARaT0Ncv
q4U2w0TV+cGo1LPlCEYykkEywL5+PTAk1g8SSuXE4xXfxUYMPGxfQSdpxk1SMqinjfUf/dUAfbfE
4wqYKoMQiVOtd7FIssogkGgvbr8qxXCHb3EINeGa6qypdMjfFm9osno5259rgjxKeQS8ZQKI7tkK
W9Zi9IGOPhDo8eV+o2D73p3+236xSZeyoIMlAYEL8/0pNOJXSz5n0ERK8UntiV5r3YAGrDaSbCUq
KK6VXL99GcLn7+01R3qV54nlG/7XG3lImcVa94kFecCPIJSgAeWYS+E/Zd+WKCARUDaJ7PycU1a/
XNfrECsiLVPJqwn3X6ivYyNcKgzcZByog3RcFN6gJPKOgUHRfiIxIDTHxqIrAEwHLlnDmqHEGNbi
ZXmiAQtRwIAxamJRzmiCPziI2EfCnyiVKYeRnwW1iZkFbk9sFR5URlKRxRqCEqBFKzSGFtWsslJO
zoxQC2Ga66ck5wGfPyn336eqcuHfpnwT7y5zkPNN/GuatN+3Sy0/cH3uWYfCroAHnBmu3VlhBzXv
ZvBugP4JqypemeVJULBr8MpEbPFc7QLiss1dh+12+FAgTxCtq7YX39vW4qY+pE/c3KgYjms9p0Ex
jv9wZQ0r/XCoSZNbJBEk2qMIV40LMAFZdwfE70lG/XCM0uJveZa944phapJ5+sJtQGL6e9kNMTSu
j29cBFG7nNbfexoYIb101G3s0Z3CkTF9s0R3WcritIUWhNbDAggCFyRaPH4BdHU1r70oNCVBAYdx
TMx5CemnwJXO31uF7e0mPJv++iUOXGJLCC3KRvO96hBiLGjFVzjgg+10nFf8uwmwsThDPYWxURn4
XAttZFz5/V9nawBDZrrPHNZnsuolLEnuJ9gf/J40O7+VZQKucIkAqP3wES9s63K/Iiiq4bEwSxbj
Np0kM8WSWzn5vEsHVaFwR/mgyr2CW1f9ytmR/T0u36ozyrWZs5oy199mkYjHEmpnjuP2RwxwYvd8
dlm1sibAqM5a0ExaWl9byZ+7kzqkWi0CWryMHx+5CHfBDHKyVSed/pF5sXpLgFmA50At4vDswCzW
hIWv10xXbfrzN5Zb5My5nQVVRqATv9bdQ+ho/AROzo+CQEztjf6/TR7z8XQJP9PR40p+ODKVJTKV
Yel+iXVqdmd/lGoOjRJ15e5T+0Oekf1XS1hlqj0MlpsA0/7GJR4Sw4D8ykNVJrHuoeCZzjMfSlx5
yZ+t65+xujMg17+48BM96oAgy8OXm1k2kuywrBeFkVsGLF3jgMWmeTHjlPbr/GsXcrk9ZeBq0dzl
ua9RBwwZB0iETBUS9aAt9h8ztW9LuDfQedBcMQpX9RcRBIyNGNHPRY4x3oLxdeEzYbcPXRmPnIrB
BZ4le1w7IQAt8LaUu6kPLxugg2yo6x4Z4mg/plrVHivxaboOGuChle7NfO+RUc6GoljKTIXjVCwr
s2/e8AH8d9Hy5pbYpmzNBLJ5l5j8WkT913u/q2P36m24t0MhefR8der88A1aB+h0Ayt1xKMGvt6Y
EGFKtW+7a6sFQ4jPHlXfkszKhOkrjAmYDWJIP5Bvq24M9RD5NJCb26N2TC6EVVu34wJxgAQdZxh8
36XLj0Prq81itysjS+Lpggq+MFrDFrWT5SY6bfyYIFDfNhwN6DX4NMxym897o2KC5p19L1vFlM5O
noozK8vaLoxI0vTMdUtbhfs7tNChmupRvXURMzMo6RminG4N5FSBImBtdjwIZoF0l2AFlqu5AZKP
QpMcXcyWuXS1cRGVFC5SRPDo0FMcKbntaAnHzMHPlt3gXcuQOoolGqILIyoAjm/ipYU6vb/nk84N
F7byBOgbDWHUg4GH629P/1taBhZNXctyDNy9UJMhiMFCz+MHhSHuFWnC4DhNLyNEyRAS/hvWk14c
dqiFTuXhiKSpmzxRMxJOOUseTWF6KH2nSnBmw6zWDPddVgLDaCx/MH+/y2YQjKnnexcxDuJ2OY5m
FUpPAtWomvZhX5KhlALwlaFD+z3/Mwnr3q9xKqsZjDPdLs5J0njFNcYwpEd8syuw9dxnx31elWWX
eU1kX4CvVWJkcLIbzVBO5oufQ9BC30wx7KHMvPUMA1yxwxrjT51wSVVYm3kXoF2G9fUHCYD6kA4V
kIimOlwWbGNejJ4to196O22PdyuEV3EsOrcnbcI/TEWVl3nwMI9dg45GHwZEqQhoA7bVQ3A8h3DV
UUHOvyv57YrdUV0LtbdXeHfJreVWwHZjnBk8WNCDQbU0+BVDBGgfDwlrhCRK2xScKBFkkV/eMNSm
+qy2agfzT2b2c7BrQm0YVVTGUrw/8Q8QXiDlFAZOwPW9YPmki/WrPh99Fsa3mSYU3x2Ejx/3JnXO
4JX+mD+CQzNws4DYDTi6ndbaNwiSbhdg8F11Se0oHJTyonsnvzKT7cxTe9XH5ZgjmAgw70f1u9rk
SE4YHfo4//GAvZH+QW3ApFcfPpxupadLlXSsNSg2qcIX85cvyIKkCpMV6Q36+cZn2F0uZVLnjZPn
RTKb9OOq48tKD9w0vaAcLCPha23xu11mxKWaqNbmJ79PdzMmgPilddE7FognO1gPDITshznoZOv/
2peReeyPp1A9bCNnTxnzMW8hKmCg/XFr6UXZCEPH45S+6RVT5fRtmT3mnki4p+hjIQZEKHOayj+5
0AYk1aQQsLyhaOL2sNWZOJFA2VoCRJzTT+AFph7rfdS3XAJUEBI5HheWzuIoqbGJsjXmrYJsKzDI
NSBJPiixHdOpCLrQGRO6wDwiFSG09wb9Ffqg5M17sWIJ3HqcARU5caMlnAYnvfxMQ4/lD3VC+ePx
LJb8+E2+7UxLp1mMXWwSXZAtV8VfHn+9LNjMmMyVpk0WlLxmPhzUONYbSmizzd5c54BXYSkKX79U
/jH6cTzcRdgkdI0o840U9WHv3vpv7NRB6+mMKCz3W1hSemtWkIrVp46uDI3c3XihEGYGJ84cIQag
ADLAjH73QvAYenAZxGOUHqsf88mIr1n/1Kl5sbh7Hzj7uJeQp3vFbPKIKy5X+V17wueea6/XDO9Z
2uU2rPvR6V5IQK6UVLgwk7ew84CgR+lEK3xi4dgb6vglWmUxbrLZkcKIA61RXxPDXqBYq4GkXvK5
rEYx3s1zs1glh9DqPIk/YUtyWdKJoaTy/8NKjX42nA/4OVRPA8f0Tcb5NJG27ovB+XuvzgEkYzkB
bvYJI2MuwN/BMjJ77xACllFO99lu6vtS72uUtPBmhat5XDbr+nNDqLNFKAB2b+BPvsAjCkYU4LCb
i63Np/klI3rgVSZ3VS/hKaajob6M2sBk4vbnmY0eRNQenzDZOHI3KRCWMGHheOrcuxuyqTTt4JGL
sr1zc+OFZ5Cqn1V0MQUR8deE5XkpqQnXAKy7Q2Kd7SGxdG85hZc02EODSMDhFZip9w4q3+9vxW6j
1VGY/UensonWNXKG1DqtqFqowO5kKsVl0c8KGn0sRdb90tsPayPr6NSKaYsHeuMAGT3AhLUZuLHl
vGDV5Oj0tYlI8CtrClRedwkbQKvJ/fUTVv09THsm18Umq+5Kia3tkTmwuUHTP6C3b1nlfk/dNWjL
zm+fcEDRuOSVun3o2Z+VCf3+bQ8IxiudCgQ0bOeFj8p48H2K7zO6y3mL+/Biwq4cMXHIvd43yIej
RmYHLOrL6juyeGz8z4L/+ipSvXvg1EQArxs/zfIiq7/KV7Uzix0HOlO9VpCBl3iVuHszTJgoKTLh
Ct1G588UT6EWVNILWbNr37TlECEcR2wPGk1b0XWYuSBXHpgf8cg4oYPrB3f4ySOcJBquGJ/LJrSn
gjEDqDhKuwrBh/AzFd6g4trtl+PLgtkienOdYXAwo3NQgup3n0wgV/dxl223cwcornsojDOg2h8x
jhMdKcesaD8DB++sA05Ovu80fpT/vsQftktN2QwgzMPKeL5aQVCqrHEqD4htvid+WmW+YdxhMWHD
ufNbEb3yXhSOfUaBXAIkdOgo1J1hkE5Lgs/cf9LyjvwBb0Pcn4dMIGNZcCNWg4siQT88PFSXlsSS
s8UFHYRYOOAFJBvKxp1k2WtusN81/Wh6Xuf8kGIE+Xz38HbIXsYIrz3a2zGJLOnVVL+Qe3Figd1s
Zsei3QenmBO6BwWdyIZLjfv+i7xbUysjJ/N/QEMrxfRDIEG61XHaHyGRsZ2YCO45sr/crrHsQN3Z
D25DC5RnlH65ob17eIKDcFPIrOUOsV65ZudLv/BfyFgNRJy0QNWDM/MslONFFc2EWNFs9CCIy6Kw
ULln9D+ZXkC+3lFsrSQ4oMH1Lye8Lom1VKSkjgj8ZE4r8gDhOxudKLdDRx8ptkwQnMBG95B7ah50
23KBn7RhN2AFGGY0KU536TB1G6InF+Zt0Izh1OWDkdnsppfmXwWNdEcGKxXBt6h3J7KdLHRNjWBK
TsqsCBDtkkKL5MxvTY1fu3p9YPWreZOxfAM3g2fRWLQEkBOsSsavBM4JQaR6IjyhQglVLc6QWL7Q
hQqYUgDQVipNy1sV0aF2VDaxYUaxTfTxuQ2OkNK/1IJBcZ67mPMfQDaiktI11F24EmCz3jTjWU0v
Hg7Y7HEIqAZFhL1g6ZnA7e9HLy/X4BH/y7YN0OksUfH43HPBmGxLhCQ8FpFA9UNPVB+mDQCTFPmJ
N5SvW6V7jxEyAUjZygqGedgFNcafld82DubjS22Ep2tmTUNOxvOB+8vGfh+/odD/Bz1sVMad8IHv
eTdHB4XyWs10E6Tu2uY7Za0WVokomCyknuJe/Cc6QjpG8kedSueFGRUARUNpuGox6TmoKyinilhb
5yccG4wc+68nPjjHDkqv+9Nk+XvLXj8p0OVznrked8mRzTWMv222lDwDe6H3H2ZLzyqr3td01o81
rlCwxZ5SyK8a7hOmFArVHxCnYTPUre/AsOJ/P5xAiwcQRKdaHCehU8dJYpWKigDfYaLIa80EBy0M
rPWZnKloJ57MdjdAIHmXlAuut6YZs1xZ96A7DiAf/3CyG8jnqJQaEil6lm+D+xGjG/YAWxUCxn2f
DXu9u/Pml1xRTzXhKvfuMsb+q580d6hSWYOwv7EZgCH6M5FWuL+xJ8hstqab9b5EFoRkXKU6KlqZ
eFmgJM2YbYVZpdmqyNBL444MaHFl9/lS0ZIA+9cSWpW8fkVug7Mx7WKIsXUaKyWFRNUw7XBiCmeF
U71Qn7/PO4I4nr1SR7iepXi6So7c7XNlnQ6vHk7iglL/tXgCPesgiKqxdH8CLQLQEXspycmbh0pc
h3Y/h9xAz882IbVaB6iHrk9nrGSBj9ims2qf4Oe/lG72whS8GMqAdpoX5PMUR2X5w1XLy5ibMI5F
TtKgWOUU9ggwxGMGRXEsuPigxfbXHxZPc+97Np5eWVmq89kqh8+9de4o0adclyl3/nRzXdJlRBFF
6Lx/gEHRA8xQGsx4gRoIa/XvTBs5DOu1rwwmThrIKCssFYMoROTU+iMiXlOgQOlCy9VnvVnZeDFY
vPy9PbBrWKDJAr32lIKOj0/xbNMRxw7qyYg2qFLjo6AaYSAR0e5uGpeP5FtdT/DDLYdQ4zKTd3Uf
OWyhqiOnhcHgzXu5HrPhr58sixX+8Ru15t4kT3L8yasK+k9G+7hIHcEahyPnMXsRHqlOZbm7dF8C
OFuIFvYNEgLoUIOqksnZYsGb7eSqKDmCklNqOlUHf0dgCoQIiPsNaT8D65Hsi+aQcC2o5veAHmlg
hvYuKCQOUn98XO7Lq3xvYpx07Y5EomwJbzQwCK1RaqMCsjjcZOUZAHT0h/C8lhEWsTdhwlVduFf3
D4lCF1mTxlEenTyMEzvatSBp0YNwFyjDL6aRnuLdKfYlBKMPzr3SbNFQWufSvhDzHwKUEkiPsxcj
lzzm5dF6l6vxMt1K5LZ2Q8vZefg5Gj0V7NdDep0u2jJBGpi++XzK4GitamxdfMtexV+AUk5StOKK
luSXlGBECk9PTHGMPwFU8EvOMVK6TUeQ5PpI4PfHfdJRekGSjeAbLCBmJYgibQ1yOjP37RXottvf
9X1Q80tCgJLfCoRy1+ISyUwiwihAdPsWXHSYghFWdyoi9sjD8d55wjeAcKUcmLGOft7kzMdEeGOt
b2QkiVEI3dYOZEVV+226U2ylgQMapEf2SdQrRNSvbe/Dvhu/p/d8pcKT+liS2fksPiWBhg9ojxcI
quu4LC8IMSTsxKrho/3fNgE7NKpxOO/PmfigM2SOwBgHy+KIO6e0eQ2ePFfruhm/A2hZ4qBS6Sjb
8IsP/j3C84jXBCzWmF9nYNhmwbmdTxmw2SDjc543IRxzE580F6WXBbuMCzLkasaiQDAQFNMvQr95
9wmBil7mo+EpiUTmG7RDlyFi4TkmnsQJZrcODsnPwD+NnuzPu3/4BKA3MomupbkQs6aMTo/ZQlZO
kRPKZSwgV3tHhjnZ9QZueqRqCFG42kWihe2dbZShHMdb12BuzVM20GFpIK8f3brpW1MzzMaOf+el
XLzL5AnNzZSoDVQS/XWPEWumpxTsKioYpXPjS46JVTOpHjweukD4y6Ex3yF02mfhZhhSzmwd1cI0
IfTbXJUD8Tcgfd0eyRcPfMgl4KOcMOY0obbP0OpLclzAvH8aty/yAi1rcYI8ifc9yxgPml84Dhl8
8gVndFVDNLqn868ga+ifn6lU2opneTXoddJwFpGoeV9fq9bU/j6wIUr4t7vIUvjUOhJd5BxybUV5
AQ9PYzVp+6/5dQHY14xhgjjUsDrN4gVM0B6iq7nlDGSitgGl/M9512TkrYjp11508gMhh6IbWnn6
wWLS2w5cy5C5aUqP5JE0z5VFOCmgpqsFbqRrqmKsjpbroPpUN3ikm0ASHWWL2zRY+0s3X+HKfp8z
0QtorYc/KGpc4MzGKELKsJLWpaD1ovv+zHUn1QqfTvwbD+5Ywzcukcsc3myXYRHypV9Lj7iTtT+Y
TJcyDg3Vv0WAKlba//nBWw34+KEM2wZPnzDHZqin4aWn7QEDFqvzLY3JVY16y22cH1Bg9ikQQssj
ChrzBrbeCI7m3CvVdh0tco5uLZczT4tdpHNYeFGCYb/F/ulF4dDOdPkr8vM/3Mh26HC4SnJitaMw
qs9sNVUTkRg5pIow9ZGNffMtXnRbA9mJVeSg1MGY/ycjrYOrh3WRwasqjfbSZ+GSOIJZAWh3YhZN
zN01qCL2jK5cmIDR1kd/pjc8WW2mcMeqJnj509ofNn1CrsBn6A9ALYFL7brQWQJFppioPYaloV/y
NWpGCtYrf3GNbJ2/EIZWTgtfGonhML6/jZjkMSRdezm68tY+fVCrZ2bsMKLXnYHhh25y7NM1gxgq
8UOPdVXTm6f7Bai2jCC4QEawk0xdrGit4EvwpgGUGpx3Z+cFeFQpbH8ttxmm6xc7QApUS+CJsewH
2aTVHg4NjvTLX41DgCIaQFZWFiRWz0U7IPMUvw0qfGFSKNtqPudCwVnYdaJGa1r1Vv+7SjjYE25K
gR41PaEENRV8LSHvqxhcJ9lgd3MRX9TBEdwm/feK2yGXdbWcHvitz4O8tQ9nrMUc+4q2GyMxB5bK
FkM7VJxg7wFL85MKE8Y9gldz/PxS7YqzV97G89prXbDemnwKrUIRwXdNDCvCxzRGeviT+cWKFjnN
hj+6W3ay5kRh+efRC51f0ludsNYQE5C6HbOfiUB3seSVMAJKKIa0LsbzGkHGDLbg8DgJRp5FkoLB
TDcNwcelLdQo98sOpg2EBdeLwLdk7J38a6E229gI5yFgW9FUf/A6b8k6hd+ascGdY4aEhcmfu3f/
ndtsz7NpRJet0o1RCdRrZKV+4KZ4HoYNFtg4jwsWz8rPz6eR1B0BZfUTgJaf5mESmy2WiBcY/9ei
xHP2B7nLuzhpUuVaoE4iTHjCLYUwQrnTRQVy+pPNhX1/0UazNPOsRaveGTitBHK7QOEbcg+E3Ep5
36kWqQjBVezUFd32TWDAXJ3jQ4nbuo9+8VPvWKvbIkxI1BaFj6R++kpL5a8uQBSg2V0/NFvDEqAJ
YZXq0X8i5VhO/lxdOEWeHz6V00mO1ceqnAb72GH2V9le5ChFC4R4SGjJ8BcKFd+SzE8uOlBubv/c
XpxI55hxYpZ2UDSU2UkmE3/HTzSYNyrVyVs7ziVTzJuz025izsVThWYw01P5meWn5TgoUYwORsBA
kXOrmUtmMb188getet3qpivftrDFM2B2oR5zdEbe/eVBBx4erZCer0xTphau5BcxbKy/SzuJrfA7
J5sLU8lqgOuHtg6jFP/etpna/35gA8z7ucQgo0YkpaIUv+rtH2tVrfA+Yhuaf/urHg9pZ53DcbXt
ZB0xAR6G/DGjwPgfRK4arLDFhxdzP7ByAFUGXlAgTUb83er+qwluqSPgwsbLiOccB6dbQ0Y8yTN6
Kvgg72Gcd4PIQGho/Yxh4YR0d+eh/lJ3Mn7rqWeu+o4BMHckplDAgiMjWoizXCIR1Vs3LEE0VCsV
5J6EPpsCV4JfMZXAiiZhmFFkTzTp+DxBN0Wfs1ZKgsXW0R2Wb+PAAE7bD0FeAa73o+bIrYD33Qih
tHoe6PaI98fiTpSGPp1pASbOAECkbD0A9U1AF4G0bFbVl4Lf0TyIMrFZjzqroHXHQhk6K2SsC1Om
0UNcKz4SSfdypu1ZrcQl6n6KCnZw44cBfs/T19Pj1uwmcHDsgF8IZtb1sYsnig/LP7nrJ3j95y2y
3SIHoTFWOyBtvBUwDGCmJdYjcoqBu1Jpeo6NBR8C9MaiAWntvZn46hjzaVSgrbammoyL+sfDn2Ll
SQ5HItyyURqpWy+tuczVp9LR1L7c6ouRiAVIVNwxz5sRjNqSaZycxXNyCkXhzAFGqMRcPIytBXt6
8CfH5gjPqcsSZTpROqdFR08tL4kbZLc2PAZbsqA7jIBWINtqC4AXcNZNnp3b7Vg13JZbmbPCSq6p
lLo1NK/2vi58/0j2FlxMoH/KASeAp5yisb6tunAhAjetgd2OEqhP4ljh8drSC8YQN/aX5CA/EdZq
EVkGEMp2CXxim0dtBZ9fDWDLW7MnDSfjGgeqYPVg/oOkt6l/FfJ6H258gSSNjbhGpUqvDrSnu1PW
rMcw/fGFlR5oyNkMbTpeasiu7cgN2u1AEkYPYU5kW2mngKBKhTF7ddADg+RjFm9KnWGYzPtq60Vn
aazcAffZXEjjMcofD7iiJqO++vZ4Vn77/2UzAk6czMrgrCYwuGyMB/E6rRQk/cOE61B5Qhs0c5T2
SBGyVm2E0dx6LFoR3IozS/ZTbC/MpDwT4/4BFABKysoXo4y4TAtPSDW9U/BUqvxtlW0Tq1kqWhuR
JVBK0lsTzjRXWEgyEty0gEpBuaFcI5v1d2SC3KejTy+HO9Zj5k+m3oq991EZ2+dbzvXcz38mOKVj
v50xgk6u201ltKGSjjbXNtWfGP0/syanXGbVcYM7Ygg2X4NOIiOkPS64SBoEiKja74XzXowYrK3A
Qu65kdbBwiWte2IuTrsurSq0ORKyAhVRnS8daq5I3PzRnVG1nj40pxxH5aND6itj22sDCTuLmzCi
bCOVG4OcjuYLFpppa3EpbEKtEZwY9aBeack7wtXz2BsI2YVmQBaiHYWJPvQS2kDBqC6HAVI8l5xu
KN7Fz59FwUdiVwlNDx82vWs3fu7x9prjJLBNwdlG1SSeuCOINTG5DEEgFva6P/du0BTpvZyVDiO3
fosln7+Qm4/nLKd9Dsrrccb3YKQF3AYhYCXCqsm5JM6kyTtasXyzGIXukPRW0osf2Ej2mO2bTBmC
jKdCYElaU/cvKPhhR5CV4Wacr86KaDsPVkB66FxSu/ilQOPHIWlQHHeJ7RT3J9rLGU4/f9TuLfsP
b4+GWv+4Bg8wYNYil6zlrlWRvzLULxPczslye2IkvTse3HROo081IfgyRgr4JTJz/+IBDV/WBmsQ
BtEBDLq0nCp3CIEUDPHnyfR0FtAU3owHTmTayzD+pdCr1p8f5QCkavtYBxLrpHV0Dm9TPfG/YWx+
K3MNcK+djxxc2gvzgazh2PGAKLQC9EwvouDSzSLq7pTY3Gg/+4id9iJbXDvJGs371j+UXKICluPs
xrXNtdGMDQohMHewpQz5VPgnuR1z9kf/KanLT934d4DhfGzyNWWh48huPWqQqLa50NSFEbSsD5PS
C5rZ5s9DtOtfPEnkRylB1gpYDEiMCXCjUClJcVM3OpAA2UIQZSnE8j9F48uGRHsCmfnhEhn1gBxX
NXJnsq5gD9nppdXUQyhspcMzoZMRWqGEJgcn+c9C5oAikHLGvYk0StiaANbYDUJdf5lfM1n54lEk
FH+Vw19DoyGLge1FeeoAAmCag5fJIT9xhfQz1C72InwAooZ6+qIJorDf3eurpFZXtuB7o/5AgF2J
COlvGJaK3EAoiptDopnuK7xSftrd+oM/DI+veFcmsvBIDshUZoYc19yOTl2UL16BAxOMPlhDYqjx
WmHqvVFE2E/s0tWPrp/PS/WezNYBT4AH/bRSTDAk4Tkni3nfcWem8bgkJ2OiLjMjdlYK0fOF5M2T
ePsaAftVMgBIOLVdjBfLqGFDFHM0gESeQHLPkf9W2okBO6NdI+KCYEuxOCZS3/gQs+8Oy6fZRJ4E
RdshDhRVZWCB4dT9Z6M2B2ChNnK73By2LLGNn7GHW1tDoRW3YKw93vlXrD3PvBzA2dGqnF26J3gZ
b/tRibXHctpoHNzwQiYDeJYop4ghUAA4i9m4RHrWmUw+Q/Th1jE0WSiYmZgUInOlsbdMG9y98HVU
YeanZu5KZpELu/i8xmHOMLJMuQpbjLkqEFZsrpzK43v9/Un6Ki+VohOkkerPkuUBcU8mgIWJBnA1
0G38rBg6Mm0LNzKNOvMeSh7+eHxomb0XH0xr+FYpmIFcmDt/7RvtTxlGgcrUKPrDCE2q+SRPUGtE
J6hBlAAScmRzrvBoPVp16NbhIOoWrmud5xbOqmV/YOATB8nXnM8DHei4kwGQ9Tha4UdftFnBTeS1
Qbkj1Ugys5RcCeqBgIUTLtvAV7/pI8NY7FtpURY8ntMmXXxbY4n+9lzrQ3a8RwM9nMjcwE9K6vC9
JbMpAG2QmQBxIrDCBt0zLHJXiMYL+yAqsof9cpRleeNcFsqooU8N3W/FdAVEztVeJ0UZcWWntoVd
MsTeVeDgrObGAFbRDNdf5oT2xB2XskKDeFIV5K6BNowyJn38DFAkqs70GoRKgXI2MDOhUbLQHxtU
FtY6Oz5WshadPeBSM3IRyOCkbiEytX7nqnpufZ0wcnBmsBQIjwcd+y9B0Jwrv7CLmEBM9Gs/Nc51
wwaYToM2RYkAnt6lyVzlQ2X3Xm1St82jfkFOTvcejATSGOPWcsFEwqfvs7Iy/u5jBkeHCQhvosXx
XaheSCb8hbCjsVmomyyvIBuy4O4aYGqAM4CDvvsi8uraBC7eHM0dfoWbXV/Qb1wBdebSCMagA3rU
5RCYm1Ms/6lWls93LCIdNGW0ekAeL4QxyxPlKdSMdpbDeLUHDANwwxNnifAyWu5X31KQXgYR1G6z
1kqN9URhN4DY8UFjKUvCtA8Lwe5e13BH27U0bmBfZct7yVkushBRpzZQP39wEu/diV7YGv7yEoVz
VhCfN4kzeLqrAZ7B5GSbRZ/ftoIfm//rqB/rfx44538EWF830ttxkas2bC8AxuZHvud+5IQzr2Y/
AVWz2qYN99QN3Ra9FqEAHssCfpHbHzDmCi93eceIclpZKAX3Nsglip6ZtU1LI+qcjXNYtYluIBy0
8KLhDCZVj6IVhgvl6eH5kfVV7VycZP7u7GVGZxxWM0dPB732vumv9MVWGB1FRnUEbGtEw7Kg9v4a
ZhOSnD6bb4Ijg6pcYkNvit2Sv/WrbbC9iYXF4EdW52hcNuL+gKnKgznyFIOxSd7DWRyOdik8/6AW
56vAg/nDRLqtS61DAG+l4wTOKaSe0k5lYo4uKyWEky7O3PbpnhbieFm8/mDnev5g7x9rmQGMef2n
Ejuko8nJiVz7Cr5RKG599vfJItcDehTs8qSSXpy763StWKihBIXh4o7v9zGOyTZdXiNLgYq/KHaa
7SKerDpnLmOkE8R7+Hwh5S+dgxK47sNHKLqUMMV8kqtOFLn1hsz7omxf3/iL885Tt2gLaI/MDbFM
M8UxQljR/0FWaZej7/n/Q1i2Gat5TjuOvI572kgMw0XoOdoOtElD0AYz+WBQxwZOOikvZQCAxP2K
9IMr19VdMToy4798tAbnQFr0BF9+bwa4e0xoiChwznIcF+RplX1vOjc3p0WnIbqYL+2mneI46gao
c7xN3IILNXXhlx+W1V47LcpdzK5ShcauD+hEGkWRJIcjv54nAIr4VC2lbZ8cPwenHT+80W+QE6Yk
qEZf7CXQBVEN64DMtQ9ixwiBE1WHJg2O2liiVOC25bb1CEI8Zk3vsFxohsVUk4WZBEEOQPmuWhv4
J19kt/gjAs9HphhWvcGWgHmtFaQ7nIufNBlUwDBC2BjWL3iQ/lWd7lSnt744eiYnOpwtc1rUiSWn
7qYooNxLh4eBA4jCTQFBRZYzlg+/5Xe5uJVV1/wVzfk7w7ozkP46haplGJjJ+tUCCm6lavyMvZmg
R7fti9809RK+g0h4lTT9FnhQKT8c1Z5WAMpP+nkyDbgz4n/i7jgGEMaem7I6gbfsxIzEK2aEYBwv
y7vvVmg2aSnmAMEpSKH1rN6Yq2r5/DN5bIHhjapG90c40uXQM/JsbZWZEMWpGjur6dDIMttfr+Um
jEwk0ORnF/MqF95jvGYub2clkNlRnCP7zqZTrPaRZ1ysTSLycjQbzxtxRrAQw5U2eV7BNIvKbarz
+UIM38Ox2PF4gt1L4/uXO/SLLKWc3/lVClL9JHa6XjvEa3S4j2HmN84zoC0lBaF/67tv0dNrIPkJ
NZTdCaGkPNm8PEviKWxMuMDVVn0vwyLcrAD/F5FYpOlANtVAvjMZSAOwpt4EflBol+lfLbFNNm17
ICc/F1YQpnRKW8qHvI4WvBTljq4Wvd57s1+BqQL3eSrTQljKBpv2izz6sxMEf4MLdmg+mNHu3dMT
DccWMG7Fi3JOob3L6onQxX66OgNModDi8IjXnE2qVKFvxrNgsSVO7fH4m6JoWrUk86RD2m6GlI/3
G6HlRt0EYUI+NyXeUkQXFyCe2BSD/AUIsCXhgTRIBS9uDcRxI9tFj7JucZmlsWg5QxV0zUIAC26r
bH5fdVEGc68K+nryWxvDvfCE0Ur9TUsGxOfToRN2Iw186qtrXV5MrVrwWTfJAPz4NHb+2IiQ7f43
p2q/wNTIKwl67wVEwWi9UQEl1PqiLWhK2znQvMDRu2XaCidnzwlCoerirjXZAnMD/cxjFckTGdTk
nkkcmeizVMNwRpwC1rKEN/x4Og2pDX8KWEYmDfXMhSJIKmWpoBPABLsajhrxr6qEU6ifn2+eB3kY
pffhtSeMxMasYewP/TM5wT/SRHEVEH09rlL4+Ae1Vb6QXdgyAIrHu3M2MkQEn2r6cj1IsOVb6PKq
fbFv8XdRqM8vIlGIrt/fE+apXkSozS/mh8cFIXck/ID/5mI6Glrxb48L2K4yOjwhjVVxPJCw1HvE
lRSdHjn7sNvxeqzNVkyNvqSEi4lL/OE5EsbuToiqMHY5QwHXQyy1H6ByetLEoyt366TT6bW3769w
NPPGMvIQySJReOqDRL9lM1ihsHm6/cZDSTU2AZ5WHNeDSyEChCIXlZGe/Oy90pdpeBqf7i5cf1J+
4yE3Cj0vLNY7WtBnKH3KqSau3rJjBDx+yR1UsEM3+/DkFO4qaldvS9EwtBFIJ3Qp4H+RJo2zFq0H
qdHHOlPjCrJiLTMsbGUA3xUBrXwTD7fCrckjs+fApfWVadYfWQZgQtjxvguuurC9PfajwF9W8NuY
SOsorPljFRIJvABi+WT+9Vx6bHWvNAMgn5MbMH3+Ude7gvSYrsNsM09426MHKNJilMtVfIssV1EZ
O147xRH0lDLJszqmrEbNbaeHXyZxiM+ttGII9WfqmdEJuet4iHFs4wrgz0i1d1IFQzDXC1Qm/knB
DkjtOzU0AnPBbBUAKOhgNMNhkRf08cyr7mbaDi1kQlDswF6qQbLJglb8RnlKoJTieAlnSqnn1x1k
FB9U1CwuCa6rvHo98weQb0EMlsElJdLsAr1OOKTE+4cZeslMlDC3E71GvrvJ5Q/GI3g0UUzAli9w
PfrYPiPXEj51IM+KXq4G4dAaMA8jZrbuWFTgwJlHeuUgmM0+ZzTNkKyFS4gbfHT5Y6+eJ+9WTrjA
X+qxa7fVcQ05t7fs/dBqrNc1KbhRuuLFokzoi+onnhcFTb7PGRKqGYcWeYyW0llW84W2NEKhGHyl
qJIDAWmvUI7HcmbOwnU3TnTW54LUmCZ/EmYKdDiqPDjmnLQTHQRNJWwkdeRPE1v9W0E8hchYA4zZ
WnE7J9OfyZONgw6z2u2z5vRMQDogA6JfSMnT9pwFIqWFcyFyfeRZXip6KQ6bQb5uZIDwCsmQ7h1a
njEaK7hw7+sszsMbABXMi9oZxEa4zg6gcZLx1OckCUtQoe2yRsy6o58WdgD7tMKtK/tAZsg3IRF3
W8PqkyxoIiBnSMdZ+uTZN/5FjDLbRx1240dOtZjbFs8NDeKQUFduJuYKo774JF0AY92FzEO1LYds
qRTdCrr4TxKLc7nQtP+y599p9HwgaVMzvNmTHz96wpAbAZECRthvbBB13ffNd+xAsXSf0oTGmDEs
grK+1NjRAYwGieKnewwMz35+Vfb/0id0uQmS2aCnMbhJgJxCLNPw2+udFDrYzHWkIw2EJ+N48Th+
T63ifJBPhPnpeyFnz2IpB6H8ScHiIrKhmkW5vwrStUu/unf67w4v86k6EsH4Zh55H8CsLY3nl/Ap
5ddNgN4ldHjlx5n0NvF76hf/VRZR6Djm11YFDb9UUlrn2FpwB4C6CnTm8BbmbBn7EZY+FOnKLLCz
kcdYB0JhsoH8KjpYRMRRUjCnaxeUSiWZtBeqGz6CLdFyaG4ymSwuPX4yF4lpPuPkl64ihvysDv1T
Brho2Ddktedjhmvnw7V4uhRf3IVSE/Xqmh++W0cXdyE9GoYhTjUMqtytdJhlsDo5N3azUe5n4qiO
BhipvCIqq5faB7QPPm1Y2sPSqeROVmfE2IN7p17Oos0CBzlv2DB5DPX3b9VECMqeRTtxe/eLg8SX
SUx6hIR0MHUPpbJWxNzLsNYZ670yGsBg7AYFqWG/Nj0b3OCDSDm9rTT/FI0DKhe2Ff9RXr84Xpjf
N750DhW3VmToY2dBXd1K+RXFyAkinsD1DV6WYhmEvCH+/lx45UCjckEgmD/V7CQb6LupSOocNImv
czLTxoQJLQ1CTeXrPqmJOTOW8zcNxLUFjBP+722KYpC20ALxC9aCjhK6QmF2ftRfSyEeW1Xphbl6
2nH/9obOq4+SZOjNJH+HjpiqYggzKA1fAmoRWLaWBiKv2zPFeenKD36uMWcyLy1yuxeXdCMVv+eG
RWrHAJRCA8A5lfGQUocOrWNljJ0sJSK25pWqJLlGHVUwo/09aqwocPrU+BrmEsp+PU5RvuI1v/d7
9m0zyk9pC3YX3BLa6cglCgjT2kF+qZ9RqFflWPIjnkjK0uyfJzSblaWjM7qFOPURxU/qCH/hUYTZ
+IVZ9tvtiGhsxTz8MEa+x3lkrT/E0fWRXXeKXDF1gMtoD/IWo1YCzykwUkF2lvB8plGFjGFR4U4l
OaXX+MmkwkZ8mQVVC/Z6STHXmSi7juhmsUjShUFo5SsUdyqQVhXNzPG0usiqBno5PNU83dpk7+PI
TNV/DmaiLPnbKiae25wBy6NT7J0kgYDQmX0RDbP/7fVzO7LyB9Y1zaMMzqMJ+p0O635bTtY9nQJS
U9LafgoOz02wjkmPkkLpnczkFnnvqD6m2XtMsuq2s7pXv2VYqg+CSXNjlyoZVjwys5rnXy/4A5vS
rEz7ThDPGuvlkz2/vKkeO6f1z8Q9DCjNiWwm2pTzx2+AnTK3umU6Akf9M4kcrHee7FG6sbZ0Q1BT
IUdJUKZ6ZeyE+z40X4Y4NA0PvaRcbxtzxXetMHcZWv5aGh0WGBiGieGWrWA0FUWi/Xo8ai1YgfHo
N2d9LTvxd+KBGnJmTKKOtHSP74elC4Eqxuu1dhpVcEkHTDMPZUE4GbOs6HxXKPadyGtodDonEzi6
qTARHF/e5KdVLX8VWoUsODPzKSVd92w79xCgoduD10Hv1LXzCymTX9vdZBKUOEMqZmHrQF70Ou8d
XcFmqr21v6Jp8LcQG0GDEDtIYtdxGarlDDXBANoRdyYW1EokL/faJNDRazjnlrOwFO604IW4JzPk
90xKQGwSgI/68ghKeNQu6SoX03ADkv3NznPU5UrkcfpC9Rh0odwC5NuHcWwLD+hMRl0wBrmPijmK
Y+wlxCz87jX4w5JmX1TKi2u3M7wOHIfDDcJ+eLMieSWOr11+VPNtuwml1dKkDvXZQDFHdQDzDVPn
s3JLDQoIOhcZXl4fFysO3Rm3T6kgDupQ08PWu8n+a4+seJCvC7FYR99LL/uIMRdj2bVd+Bq5hndx
wBYXSm3SVPXN9fzjGlAv20mT6KDE8HXUrYEUQIMOqQfARlVfGgX6y0aj5CxC9ROniICZ5cwlWuRz
9KUoYF60i4Tjjldx42RkpQAv1ADNMwDBItLXCxoXvB03cJx/SNAoMx68nKqzQx670nPYlTRaHybj
F4fxhePDxEwK/D0pvdFONohTQN6OJ9LwRTR//KGyZWlSnV43Jwcy3WEid45DjUy5gxagHkAIbnNP
cbwWAbD+YMImwrzClwCzPyagKmIoY9VJA1L1M0rx54qeDdXETqWKL1OXoV7DjMl70byudDkg8gAR
8TKpPtVNC2zcb06H/Cieu+5H0qIO/vlkHYz4PMDBllsUODGpvZ/zZzMrlOzzwhv6JyOwRfmTHefO
7oLCNqJMokLPOPPHF4jKj5/HjO9zVPQXZLWd3hqZLt5tNyDy5iqQA9tB46ExY4CDYMkoADf0WayW
yNHuZtnjqXNVkFsEyPT/OYyV7WKu6fMvK0724kSFFpv1IsiA+xQznRp1MUNASuvBt/PgsIpVWELa
VCDt5RkDP8Rx6yNt5mVbjtul1/eyTB9QVM30xKG0xtQ8X3TDPAVkebm8osPAzLRpgvC6k/2XSsNo
DAcWnS7DpFgEh7umKeebrfPoMIAofzx5vfVa9pVoyRXlXefwPXsLhOFD8ZOeyUcKgjJKyDbbrtz1
6R3KFnuY/Qmy1J9OOcIOJAvnpzPZUT7HL0CpPRA/VXr1U08Z15JIECNOZ+j9FNo2XbPJLdyd77bP
cYUnU3w21eT2H3REFQx1PzxCWANLo0qXzj9qA16+eLVTye0OMbxERb104fkrPA9iNhnbLBB4Ew7K
VHBIVyklcl0BG+My5IkcfSeTdWMZzjuCJ85IGj9+bESbQka21wVSzNGzn2Qm6E/i04JkJfwPYoI0
iKaxuwB2Z97d8LjLEqrn/i6Tq+9Da7NQytP151nGm6sd7iaRIUXaK6YZbmpzHOi2pmXHUSNaJ1HA
2VLgC7ppTu2whIHlAf2YZOq6nQIqqb1eWtUf9LSentFWBZMimyi7f5K4vfDGwRFZUg7ZzrNkZ+/A
7lntFesXXtLQ9+/fK3/k9U7g3+yoS/Tejbu1o8UobxVgNMBWJbSr3VwpRHtOE40utLrDfmuOT+Cl
vGGs/E4UamuZB+x7dGFxUUxinUYbsN2p3JWE0oXxpwnJk4qPshWI443k0yixmtF4SbksfBS2FlrP
arLqGZABJUmQORY+SrqE8DIAiZ8DoXnKQU7gucdcQKlZh7FtzwE0RbquFzNR2xlQ/NVderDkk4Cv
MnylUKp8sFy83DqA4MkEXT19029GCmfA8iWy8JZJoeJkA2q6vlIhK3NMaZm9akx2SKZUdtI7B3ZM
YnX4NkuvJcKjexL1nXZEfYMmz0OKGysw6VW6qOCS/cEN+muS3WSZoRi1IOBcnX5kIxSbFMGnANw6
R50hsWS2SWxu9oV7DfU/P4DWk4I8CkIhFgMSDx0BcuveAM9Pcvs8odSQi3GNuM9/qfGYQHs6+94B
GuzD4pl9MX76VHdQJPNZEBnnNnZnNBPIZ0txEJi7bXFUAUwYGZaQHC5tt+mwG8/i8uSI3tYUgdui
nZQA5Og011FKZUtHghy3DmArnkbtjTrX8UbmyrFhSHMkgvZVuXJPX/RqchZoX8inoFZJkq/7DohI
oB2pqLmfZqP0ypKN0fpuVOJeX+fusFAjqNZFRcFeWDVKu8dfd+CKrOJu3ZusNWyWjVJZZHfjQ0j0
o4Pr5ZVLzlmkiNr1UN7fJayV6J6CXBpCdmJ+n0Dmc0IEBf+hkZPfrvjIFfruqk0EsHQdk1flecco
Ua4p1vkZCCv46E8iDOGu9lel0AbBkFcGDASGYGT2L9nLWYUTbWS/jA7Ancj8aMJvFSWfKJAL1wvk
4sMxNDYpFHs8x6GMv5FeHYwDjKmll3o7X7SOdKeBm+GvDfWinhpQjL2bNxstNdzBVF2rkKxBCf4G
RBbykjxTufW2t1u3Q61u8NTftXNa5a6R2QrE/7wsC3NEMma8XVRrgVwZrMJBHVltEViEvdfwKMHi
TjQpyS8jKyMDz5exqyiLmOJE1T0eSqNGZf6hN81AK4S86l9f61iSnExNFTrSs6iMRaflCHEiYVUm
4IRYvzoHM62OLokdC0V4xGrcTlc4j8PA9w9osITw1WXPGYNJSiLhDfiZzDMex27jY/TsIdxdrKJ9
RPEFU/kcklCG/xV2P00rkrN9rQRjeKZ7g29NIXk5QdPHX/GW7eigNYrytLhCeNWidHtBH/BY2Xjz
D/tsQ9cxkS6wfoeQqCyWazN6odG3rwaWyHSVfd4iRji9YmI+4x71P2VARprR+0oWBIgaOwFtVRLf
e6ROPVhf15gEEo/Kz5u10b7zDqfBM+yJfCXChevkJ7gJzsyAsFdGfVNGlspV1W3mSCj8VGVTsGp0
ERcShw++VmSJJcm+Hx6kroXrNZ1Nr0p+QfLI5aGqkOItUew/f2opWzFyoWx4FeCchcPZSLue29vi
ddkniOUn0IRA5FUI+9kj7V6tHgwVDM0D3HA77203Ohj4A0a/hyY67kMimdqzInselp1eZGV+c87u
Gkg/fhlxajokyIfom2/JLTGXt80nTqVLJZ28TxV8ydQ9wTcHLsxlFaGdRaVj4Z7GaVnnFaAR9Uhm
68cQBDn0gYAaFbIRr+sAxX6gOnw1apdxgu4O+a7csfK5nG8OQPrwl96rWyeBvmr5t+49ejUAN5dE
mMBO3WNeOUy0kn9K12ppmsp4wfLmAuVFlLO5Y82Tab3DKuL+V2KoCszxEvrGVbO2ghJttB7NvqPp
N0nthMLXeomf/7lqRwBSsDdRMQCkxzqoc3Dm+u8TOY3jde9ldvxXpsGKSYY9YTWhV/WyDZ0umcwR
GrW/FCfY+iS79FE4nxnuchHkVTR5SpcyTz/BprttwJZ7WGpRxyxuN/bHJ65ZVgfbtEPx/XPd2XfY
xOE+Xk4jnK26X1bb0ypvMYoDFGwFP6QMVQ4dBuyeaKpdLn3F7tnBm9apzloDgV/1zq7TfXRzfkLS
CHt/j0RA6D5FB9EiuS2nAFkya9XrlRxfFJ4buhrpPeed6DFUWOK5ZkOFK4OV6OgSrFZEvj/9snV6
MuB2baqes9a5Fduz0EZvx0WhgSLOhZ27Sm7cR3BTux7o2e6oiOUSzrW8fXqXbOtiqRD9EifRiXWU
YS6xpt3Z1wlXaH+037l8MJp+bWmoKCKu9uYSUKUA3j5XqHb5grwUJLV7G2MNW2VKRH+fIzHp8b+k
k1vsjArIcu0UYai7GXYPuKUIB3Rp/LKEk2jQSbW3XFDqa+HC21Yl2yWBrhzAkVXspI0Kp4DWiPZ5
5gulNDPQomnrJAENVFQpaAbY89jvOI1VAMV86kfpWP7I1mkRgW5YjaXS+mTE46PKVfqBNWJmF1uD
buP481NWZlgewGsSusslADsJihq7EBtwLq1yAh69BVd3Oa7uVwvuxAx7uPZUbE2jmgZPiPhDGlf3
epgBMMqZfdObcfgPXEnsAWpxxT84pTNuzsZRFFg01enOX0LX/dZlCJciENivnxFyX1Z3NK8WtkFb
10jFpznXcWb0/U2ue4IavO9gUBolyEhjnDjrL2PHkVwG3vMhzVsPH33jljTPMlB9DZ3Iuu0H5ig/
llcJu65BnAagZK/6AO7Ji9baAkySzUGJwboctbILH1zjO7fDx72y2Erw20FYaPJf9AU0gGjipOYx
oHmIbDxnOHzD9JoJQnhIWj8l0AGtjGneMVCtNMJrPwwFGupco+rf6oe4CxY+6L6LjBP9UbuGzQ6V
lX7VSAKMrShVxZ3dAaXSSytn6JZ9wISK7ocO4128QOAFEXMRWGnPdaKZgMxp4gbg6NhomvLP5f4i
NxhC3CbnhVYSKX6QeC5Kc/mna4kRxGTjikOZqcLhYDCUJIEjku2ih8sXVzldYaZADGBc9guGcueC
cSaqgfPRovyoLosNFWnh/hCmM99SF5HzZp6quEbv5EtBmLIcetrSfJrtQzU9+MAiMmBREIHNLIva
sDNWOoE7Rm/0WH6DlQ0/Js/Rl5WVILroUEQtxzXlgldVppcWgvrKVNeoviEezZ9X+jFkv5ZOFpMx
nxqqiByDeelXmOHgnw0E0f1IQOEoYfUDJqwbw41MDQGgq/28FEdJC6/pqeA3hp4mRUCQpEW2nZbl
rANIwi1hxscPi9Tye2KlCRpHBhpNztmPRaRyo9eomSuqfZDHxwc3RH8ulL4KmEIysCpF9AoCpME2
0c8SkysMdkGavCEX43hIGsqzEsZ6Idx367DZo5zcgxY7p7tkwC5GljSB2Ed5y3DX6c7Zt9qRINQl
AI5pLxufGfqsmS4KowIg9ogzNA1O45gMgaXYOhgZt+7vdqH/7uRgzgHmAJOxdMmlG8uGnV8sS84P
5w5JgOrDXm6uTU7PtZSltKaNTRDLCga+doe60VM4MoJpwTnoesJwjRsyyDVpf3RQL6ZWRrdnYfe7
3dVIUVTl6IvUfcU4+z99xLiafnzjCb8wSn7fBVgIZ1sSQrbw6kfWXPolrnJLLgl3kEzDH2emqQh5
xCoeCJKw/6YzHB2lvQNOiIVMy5v6IQH64wla+0fQ99RH/Qniqowa+4lnio0ccfAd/LC7DFpmzuEL
lddu9ke5WI5qHDExw66tfAbi49KxV1QqJYNQ93vwfaiE/J6P8XYSiZwL7LCOtLiuM/KhXmzrKtA8
OjXB91LbyiTb2OinaILAfq25b+XpGKJlGsV7Dk1YysNEcF0fdg3LXxijFzEV3ICG+VtnMZ4ByaNu
ZO/tsgYxXB9/+eD2OuRh20j17twY5BcttjeSIARVrJcqS5zS2Zcla3tN+T956svGUh9BbyAK/bGm
O6xssGmigrWfJg7lhx0VOxTMcbFaNGCxmfYl6pCPZjVqxSuCNc+mXXmGCm+LRz+3q71zIIAVCYc7
9FhwdQ1C4bYO1bvfz2VsLUjxyiqJBFBFY36I3gMxlj25vOCS03QBAqQPzW1ql6Fh/9Zlvq6jw1XW
tD1klUXYAVH7SjuT9jXioqhJNaUyUagR+k7EI7IPpO1iKCD9ktuexRKn8Gek0HcIIwL/srzZ5wMd
iKeFNeS3ZVOARZUmxcm+0jfxGjW4SwgCWiQo3YSSVEGViCFLdi1NOC+kbYSHsW4j5U3FIDHlssmE
lyByo9OWZb+YGlQ5D2YdJx640j8e+W8/zMFY7s68QFKCY8Pyzj1hTasDaRmcx5E0hQr/CLV9D80v
89M2mwiSzWYdilmemFyO/H7eTSeV8y3ZkRlaWlpOEkpzo9QVxyK1sCgkmoG679SAKRSMYWSzCvbB
71uTcNEvLNTzZjQD+wAyXPCfa0qMJTFTc4OZIXLQRnH8Bs3oukd9p5eFLA8sjz7ysSEZscOeQVp+
H78XCv5TZrSSvrmITi5iTAjdN2R0ZmANx9wSsJ0SgGFiOmERWqFaqYdegqXaTepN5g8pdu4J4t4g
+QRMWAt0Q2yQOMbdPC5UkRv6kz4ZCIiJAlTAPOvQbv6SmOeDFRp7e6wvtfALrNH89sC1t0aaJFmp
Gb+HcnmfhyPnrCohC7lgSGUwYJXdpEZ6KuTeONZvjEXceH5cLEaQRf8bt4wK7NQt+ODVd67nmTUS
PQmdt1gCFB51uWCdLX4awXH5oZPuoDIptHwLFvBtpn1c8F7W+PF/WC5IVbmlsAfems4bohwPWdNq
Q+/BPlrglLN/aFv4bZbNzC+bh0lnAVfImxDEUlvnI5wf6Vi1vsRENV7KlDLJANnMzk/PvvbfL1mE
jx2jxQjKzOwgVcNhq0o+9yhjbZ5ZkpfdgiDaX5az6WxQM+6NT5fxjS2BQqKzJPCoI+qsG/7SH+zj
av+dVFYSWDUxAcPPl7w0scqVef/h/HCqW2p5OGLHKT8Kw2Y6BZkE+OJbBe0lNO7hxq+Z7NCFzdB+
RCbA9SoqVzVCWmWNTFu3OcFX2LKpphoeRk8k0u1pxecItUZvun9ectd0V9zVK2drhlhFS4HfmLpm
H9OOEitS2yOSYAZeLxOIZ+nePb6B3UjSQrR0AAaFdKqaqv/6Z+WrJiwpggV3w4TRjZCcQJ5+sbY6
Pr/FwRNFhVYOiVeNN7yrxPCyGaLFKj/A5TixuvTnNejRXUBxLkZyXN7Qt4uBa2ZDkxj0X8kQbPF7
jUv3XiDL5C5n9qZqDH4/kst155dlzomQ/Eu0pApdzh4Z7mD7hHtfQCxM86W66vODronAOGzT6U/c
Iv9BbNALUaaCGnokmClgk2bDmYFPtDhe4SQSj1qqT+7AdPmqZH4JPZ0eSu9/Cs6mcovhVlIOMq53
1PydCJTWZhRwsdiNxNUhR+pW8xKPyOk6axc4Zta3qbS30+Bknr58JEVAKUak59t2i3TsimmFNgbv
QsfKELXKVTH5v8kLVPy/S8SQBuWj5VYhvkkOvSV5RY+QOvN3SlcRmeIooRYy6q0dpzXiKKubAldD
tb2hbMu1i8y+7OFIS36LPS86k3XulrlSW/jyJe5rLfmYJPXGOYTFLCfYd4/prbqecfOpq5fHe0Wy
AUqbxeJ04gV1zBgnM/lVAdCz7BMpWUOxYF3eSeNINS3nQK6TNEuePs9l5EnuKpljgxDyBpLJe3dg
n4duHFgKYo38N48nHXv4+NhGgmT4tQesSUKZHnzC53wPHSvZHPTDoL/YFVFg232JqUibcxvrI3yv
aDgyIUua9STPHXeitLbQQ3o5KkNYUPkQ4fisvIlL4G1Qz69hG2vbBcHIuY3pmCD+8dt5G9lqhx8y
zVCucJPfB2Z0/Lt+g5cw+rDjwmrMtS422xf4wX7XZLfp4XQpWz8+MW2InLKUPEXkOOxJBUAbPo75
X72h2ZRtusNejurl/q2oiwAWCWk7O0Y0KlbD6P1wndpghp7Bs1TWVtbq0T8rnpVCA7njFR4cSPQY
B8q+AG5jJ/oBQgLuAqtJub33sfqr0FllpYSsmVbTkRqQAZuleXY5zI3pQFx7E8z+bxaMlD8wLBT3
BK6avFBsq16v/ptVPUlbNxTmbZrO40AMoVEj21WAL213eqOBKin+CtiYAt8hKminxhcRyjrZzSzC
9Yx7SWk8u04FDclU+Op9e+YR+Ddrp2FqRcfKTVk8PwCQvZ9GrmUJGMHQliEXsSN/Jc8d5I7q4JQc
u1cXRUFzowvF8acvq1+yJjro3HsVT2qJu1FQlDO2VIEMVCSu5TksDHz3wL+ovR1yiS+nVxOOuFFO
Sw6aPfGYdc4Vsp9PP3Y74djjIkVKsqTTzHh1+fF/TvHa9EmCT3ibp/liUR/ulrJ7mT27HFe42gSS
SRH7Fc73kWbPyp3orlAIWBHdM4lmso5V28i1S4zdErfF2yYYkRfy+tF+VI7GuNbzjOJN/pxGdgme
iQdCR+CryURhiG+7qANK8IZs9EvlpPDMWAdPWxp9H5O5YexI36LWnOPBts4cwhqsVblg30QEerez
7YLWa2frC+QQRqkAB/ZHLwSJWehZ8quWgbKN+O2OlfYmQoLo08y3NkMz8GhzjpvYuiOlTW1vQDJ9
uxrGBaXeaVWk9kxQthGE8R7Gz5q9gqLLm7FQrZeM3Y++O635kLjmfp7GVHklJkEzw5Ivz33JB22q
KZxudOTMA2GWNCRGkvD6/Y5FASVnItbatQz9T1YqJWaTrbJCJlYx1kBWAYiJLgGDxLd+0l3WYMt+
sZnUhednG8m/cwC4b/9+3G67ZA0W3nrA/aMtdkKX1N2aAENxs0A9O7hPkbJEC+hDVVMgAcfU9tN4
BVJq06AAFlWRrQGp5R0zOn0rZ5NHMjraP4JlwfpyB5VPNekvSdYFS+EB4p4HkCeIGjaWvoanCnCd
6XOiVawgnMXgW9Qo+41ncjpnorJACxecGrj+9C1pCdAWZBEOixIcAjMZxrZFNotDrmVbUfBmYEp4
OpfTHcjAkm0c/q+8bIvIrqDE2hIu3+VM4xFQMxttmC6SJZTW/8juJURBjedrrdrPQSUpXmrNwS5K
EjhIYwUiTpLG1f6zBvLXPyyzS7ApGV9hUXHPbHIy5quy8K5TOLuB41gMspo6OQpjBLgzKpXlUKD8
1tGROsmVttkrhz97wxInMNmCOyfumzMvUjde7D80ukzjAakC390Q9tXUtkBTsWTp/oRyl156H7Dr
lse4y2qxL5cJgsSlM/GC2/Jmr1fZjWLAzEi6vUtYI78Uq0GOxfibosFH+jjOeG/TexqeC4FM4cN8
+WMmuuSwCFWWbIUlUAWUiAk9Tcp6zQuZiS4hKBTeQCiFmnQTq36W7xxhQfSRxftW7qnqGNezc6PC
5kR6w0BhsxzZcfWUJpMcMRo6KcBi57VQA0MQvYf/VXE0NKgLUvTdHjUKa8xCY/dExT7EGnd7XtIY
mvda31sJh/xnzLAMgB8XPH5+mi4xM0X6HRjf6CJ+MFZVX/8dMQ44gxlnN5hqjcS8KknnOxyLDfux
5MvHVXnO+5y4s0RHGT+mSfgfV8Lg8HRfz8kOR89xUzzbGXER/b1t15SGUvH9uWe6qxw+UBqVu6sI
ak0PbsY4anFu4V0NVihLL3pncPI5AZUWVSz6kjTY1jYaCZVB9ZNm3YpZ8sJukyZ7Pzms+OnJ9kWg
GNTYlhr2hhc8osUw7Xz1inHwqRJFWcx5bGm8kqfqzajgD19bOhEWrkESAYjVg49A/c4JrlG44aZP
2EPbh4M3lzzpfVJ/irrnkt1728mrMfWpvi4aa78b/gz3GnHZYjBYWZhUnS4gStPz5ieiP3gdkhtp
H7Rb34npa5jNDVRe2k2YwzC4bZWNYBo0Nj9i7+xmlFYen9JnXtjpe8Of2mPYcJGAX+Q7h0IPhbv+
Oc1xJM51ptL4d9GfpPjDIJ3kmfIq4SJAewzZTA5yENwxNsoR8F0kz2LJuDn0ON71F2aKA+w7j0sm
jp725QsA+loQDDErND+cpFM6vLeNqdmxq0OBgT67YJAxqkUvlTC2N/ySHT6mspqteRQhOuTdq3UO
Gi7TrwXw7ATZD+Xv3D2JjGfVuex2Qh4zZI82DaC7UJCEFpVW4b/Lg+1qUGaU/wxncXjVHMLKsrPP
TK8H/xciTEAbe0T2hHbOYkLV8ktvCi6CwVJOncuZkbc+Ko+wmdffPJIdakoOiYYpFshCZgU+axgw
X5D15U55RDtQOKds8qJISq9Bb5NjuN4rFNCYhqMTzXip63nuGo+Kdaoa6fcJauZEvMBcO0Oc5fsJ
Rm6p5dNCbYwWI2Tx444yVLVYD2VBweNDUmguN630PRLOKX2Zv8KC9p7LZ8eZ3kia/S/qB39qVeY3
sk9hgvD5FHTZGADVowP4gF2nb3b/GaY1v4LVEwHznGiw/4vPoRoSak+EkgU4i/kjH1PfDKsCRkmz
zEYn27hjMurx5ICOXEP7lyYX9kNKwrV3ouKVc3DvLWRQ8p3SBw2Vwgu4Xqn8erq9YEK+ssqVo98F
HJpJpjwDKVDa+vaiaGkucZZud65NncbNtQFPtpbRjs8bmQYHQGgPdXQ7oqaJHtkVW3Gb/c9ZxY76
r2Ap/bSxM3QpvBrRsIu0AQc9vZCFbBKvNL1gSvoIvAXSP3auMcPyYl+aB+6Q5DuFH0GY5IgLZOgt
rSP6agn+qauNWCMt5O/YxKWTM/EM5NLgedF5oNRQ4KK4H0OekDZG+qAtIJh43fvwtAZdGCEQf4qL
uZC/9xn8G4dDDuEOrwCDzHFA0/PIlGkUiupt7oPdzwNd8mquexHbtYE/pZxRuIC/qT8/kjkqp+vq
IzIDTrRPt924EELWU3K+y3gSyddSGR74PyYrzZT9Z76Kjf8mJdQfSanb1Di6ZL/6uQdAi7B6oTte
ui3tgRRLT71HrxUyLkKkV6SVe7+Q1R8MfXRoorNfv9gc4NF56MCC1ukPiP7UOiNy+vAMpscDL4zj
Xy/0dPWuztiafgSYcYe6oTqeN/4hgOIN9I211IOpI0ciesHOC3Qn3rtl3ZOFDZZ4Owb/oFYQfHqy
4ninHQPvPFU8Nl7e3szc8Gqs8q4tEXIQSo1K86Xfy5Hpsg+AZ78MdOlBji9naq3bjED8K0ZqQNRB
XvxYjOcHGgDQ168GZyFd9SHB8FJN73YIq7l2q9HYb1DcrjwbvQqSaDuDaEdpiC+P9UoROth3+jj5
Z7OGpyKiW76YG6phlOTIRqj/VwtJ+GeWMFHUhUWcyp3SQqcDzG1onhyOIBGRLaONO72mfPoe9hpV
/1LfW5A40k2z9dVsR98GujL+nae3OkM4auXr18OQm8MuWdvCQQh9ekpf1sMt5/IsAZasK97zIxTR
TQ9N//MYukCDC+GNK/QzEZprWN7bLOdVPe7UgLWr5g1lxtVn11Rpd7hFVmYYJHqnF2OakP2/03j7
1gAoYYxhi2UtM+3/5Pw9A4AShKYHh/BI4WhfVaGDU7J+OndCf/IOTTRSIhwKQMpKOeiYjQwUs7H2
LkPSQNJRx8UqzL6bvrGrZzRVKt01qO6xtdR6rGNoWgboTBWEyMIgKRLwPKEu/dbjEPtURP4hsm2F
c8JN/k9bo0srmF4JAJxqKhnR07hc54cNjZOBnpQDS7iRjloGfZkF0clo+roDEzg7abydpeJ8IIBk
2/YgQEdyVXSJMXoyJjXKE1tIRofSGpI4cHY7eUfT3vqLk++7YBkuwhyB/AJcX5kb/Let1Bphr6F1
+IuhXFAvf3CMsJjtfVg4WE8gcIX1OHrurrOmTesF+Jfj7WnnrIHScKx0Y9TZocqAj3iVlwnRqBbD
KGWqss7fANOZm8QQcQkJePrNBbmsttB6Y3WMLxJ1iLgplVeoz5q+fKCk7HHzzBbKMJgBRY5whRkZ
voVMLjlDNm70ZuDZYp89UbUxoHuU1uw2vUtz1eBZJmRJUt6Ka3xHvfAeAsqcuRZuRGU1vJ6tyRAu
LAgB8OQoE93aKYGvIV2PFZlu03emOPF0esT+wFAgg/lLAkkCHoife0l0ynEVPXB508vwO4W/xhue
MQRn5aWQaHI7k7suSfN9i16wIyym3sRA7bNO2i7KUr7zH82vuDa6LxOlMjMeHmmufd2BaFDLh7eS
RNPM0V6D/fw9F+6LeGuq8W/QdSvZWk1aA/92rkaMkWIt9FW2LeAZvOa75Faz1f1UPeiThUbzNvW6
oM3kQYA0oPqT7f2eozeJpXwtr7eRocT0k31vWvKc0KzTP0zhRLL/WrElhnQHgsiH93rx90vgjki4
lmVTLbmM15hMf5BtFeEO/vZ+hKLfp0GjzmFHL8GTra9/PRlQACL/PqdSHns6bWE697WaL0WiWxcA
4Z9zeV9XfW8k0KZzN9aGzMa2AYJL84mIr1tt4hO7ZS4hg5uiGQZbTF8z6hnb2oKj/fF7DvUzAfGp
/38taSWfDQdTOfuZu+GHyJkIySdtChuY4Fq8zHNca67pWUn3QHY5EkPAX5GJ9i+L+1DKqAx/CuBS
iwbXy5OVukKcgXsEVuNFMq/LOIg612uvWtM90+NbWJAa+0qH0Hsj+TbRGajv8SdnvGxqjnlO9o02
gujaxDGslKHZZutUfu282I3xO8+HQACDLc6ScWZOrWzSScTrvtvUutZfwCaB4sHfLM0645+RISKj
NfcZIMiz/mzOy8bd/5fkxqWyEhhAnKCNCRjQ9cifMOJp2UB6KrvF5NFx9R8LhhTiTYNorxZpzplh
FVfNYpzZsxUrVOG6iertWsIVPkbdP11z5Wmsgvt3ZciPOIFiMMsyGb4m7v0TaiXc2l2BKY8gVvX3
8le4h+4Db8jiA8eBktzYY2tzcYgdB6odn56y6/lZzAK2IG7cawJRqa6XI9XcFCI1zl4t3DyIMUxv
nyN/0napW/5qjnlwlSu3xcHVoDGYHvLJ2A/L/YSGgqucF8bM2Iq1YKpuBA3/nVYzTiLYHx0asAPE
eFymXIzDaVxn8D9GKxrRavNASOtPbNuOb8fKS+LY5EQBU9JY0R1UGBdC0iP9deP+kyQ77sOw0ryP
jiJU04GY3S7wXgzX3RBNjTNAzMm5xRRoWRr0uqWUXUsnE83dXITOYoscf8xQG0Oyp2uRVTqk8Ksl
VLE0fAWnwWBXdz2H7U0InPE1X83++wU+QdyQrIpJNQNohMDICAF7YTGhIboabJPrKirE5iqd8b+v
Cu9CPnsDHFV1gEC/xAyF1+Gy95Yxrsb3wOM/bcSEhrZrr5kMcXWqvIRuTvExCc5f8FfMuQpursOO
y/LtLUlnJ7SwhY14PUuvgyjsd1wLwCp8loVv9gLHGRKL0sdYHtDWPpoEDtDUX40eyo/LIhLgKNOT
Og+zgNLeIJ+P5nfmQSwSQd2wacTbbkw5Y0yldw5PpfTvbw5nHxA4JYFTGeU8SBzjjzUte85TNsuT
iCgV82k4qMp3CliTsPQqYyEuATpv3PJruxplbTZOssUf8Mz2W4l2Psl6oUl14ZK9mcQimSh9bt5/
BmJwkd60caWlgoNBaGuRLHaW3nMCz6LMRRtED824RvSnzl9bUrrxwEsHarLJjbqvs9IKLIktA7Vm
IGyS60zEqqy3W/PxslK9YeR9IVkgueuadaBjiBZsoeS+BVnFgP7Ro9vMWEum93kypRqL/0r/YZ9n
3lKzMdIqRm0Irl9tCXEvrafWv3fc6MBpkzevjjnCFq0ob4bEnzdyg/4YWMWb6s+v+5naKy2CobQK
BokPzmLC8lp4pEP9icsXosWk+Vp8OIW5Ci0BZjmNGM4LDtTWL4/xSHUvHVZuaKJslpAFjxlO5Vod
xxx7COdljxz7FKCkKed9cCsQbW2PJTaahpdLoLMIR27XznWnzfnm1ITbnmTZsaWeviEsMC1O8xdi
4EHx644L09672FvBAeRDE+bN6VQ8et7jqSy/Tg5yVR5t+ulnti4GPD0Pt+diFAVbobUp6+XVC6bH
HafeE21tRUrMIVbH+nx4swgNkQsSqmbJWOwxOQiu7S9oM5ExAgeGT/8qrpc9ZRUwA2LKqwQLd3SO
6ufjBEdY0tkTDj+cmf9ZmgByfbNSFToQJGksH3ITwo6wkjkf7Wj7N8Usrfqhb91ErMPKtkRn/Hp8
6ExSVhiQsHJ7kw1YXXdPiY3Stk3c6nBrUpWNKPoSBj3on+UbqhnPYwfHZU9oIg1aqvVHBjpBklJC
BTzH9o17NvEHKTdStVJw/Io9Ut3TNlNT2aeaVf42srtkn4Dam3+YH8A6/HAN1zXD/SObNp/crGUd
PjloskpebOJOaSDa55UJ2EekVFdIkcr/kT8/dSBUO5dpx5no4ccTZFo5lx5pMpzNfTLoq2KlzekI
zaXsgiP+qCZPhmUJ6j6JTK+O4qq/Bbli1RNqtRjI4jw+jw8XUrpEHXeeiomimbea1HIjB2yXR0g5
kBOaRTgS2fqPeDmA+n+Guh2f+cmJ7IWh0WyEMlTGi87DSKTGPTYvaxgRzlmIZfhXk7FrGGkgv+yC
h4IYDn6CnBHv/jz8MTLJy4iI7pHzNuiIJVka/RHxVYlEbI3i60KkxQvE/WoAWTvkepRm4bm5Zsyh
h0WcMag8H3Ug2y+ifGhnHJ1tBcHFe8OyPhXa3dfuikFCxpMmUuWmQjz9yHfBBuV6f7+IZPKExQTx
84Q/uE2b1pw4MOmrMjhNbnpRYgN1G5G2wOscxjzSIfIHOqRNwLYQmGTASSGPfSIzFLeTgk5QhX6b
v6mJxHnO/z+GNT5K8nHSQ9Kx+iaeqsbuwC2jUV8SNkogKNVl5eVNs0wz5ZQpPzwiGSI2LbTZpws2
4NRirAPA79nUlZm/360uK5fcYZCUy7tcmOoOjjdtcYNaISBDrqkSRInAepOBN6uhWavfRph602lz
B44Hc4YasQ6FpoxaIuXvQx7VKCNiGdCf0JARlzkS1Ox8p5wUCtRF77fiJhr/ZuBZVPcBIpcjxUJ0
speiyHkXmjts9YxeYLPv/LQMKbO+jzuuXT6g0x5PIISFZKjjmFjv56qEBzFZW7qPXVQwIgjWlTtO
3w788Kl0d5Dlj/8bN76gmhyHo+fPkzAwKY4BMB72KbETFSfg01h7PgInhBKBJZECrjo+GCedk0Mg
sCnVwgnFomMcuAnzXNmkNZ+vSGDLMJ3kVkQfllG485BRb1CxyCn+uO4uI6QP0ureZVdRJYOktvja
CuLMjMpmR32FUWVoV1BS74ZCWAPAF9JIgOGrruUE5tVNC44XFB07TTSpMTkXAi+LEwOpFcTwsCLQ
MA/zOJFcdjfcS/Xm8/slf6YFf79wBap6GumGAYkSDvoWHM9aUmOyfmeN9taR8LPWaWRhq/wLrT8o
NRpj/Cd8U5Fc33f2DGkWIqcE/BtHueyuReBuQDD5hklfFQHp30/vlcPBmc3Fb1jdaUK37mvDq6w3
K5qAOx5EOtR6P6akzMFj7PLZCWSExWNusXrFDP86PD+jfHLvmDJZ+cLyOAUOBMWqWpPTQ5Q7gwlb
PpIKa+NTB/6XQRbyKKPzPHZsB+uUcXIdTPOp+cIBsSlmnmxNPDLeSzOtQJWNBWTuZpDXzVVkgEJb
VhO1GGvjhEp7qhJ6FcBE547VkkxiLab4bS2NT9hZp0YbsAC8eVhjHOLzFopZFk+5lyYlYhll/+tH
CDD8ShDIDOndeG2Ti+1rscFVkSZhQbnhTl5nzjC0kHzzomyR5hENXW2E4J9r4C4yG2LFe+w4yZAo
LbIwudNNNLhejGeotkNJnLlXiyDrEjiLJqeTbvhGanmuC5pshSQT3R9zWwqpUlOg2IKHR9/kXAti
XEvrugN9VdtIPK4BrqkkKjMMnswOsObSjutQmRozlwuPjmIHE/wnKbQaSrh4jCaepBaRZZ3uVSgG
DCDZlxYt5SXxFtQlL+SF9ewAMXaSFTsitUvAeH68m6m4mV1/UhoLBNElSTB9ztucsutsc3OPWpFM
RzXBdHjpQWGVOYBek8SYtPXqAbNO/JLrW3eB3Y4DsTFkN3eR6fV6FpJhb0QA39xOZKw5pDsvYLI6
j5ClxuoB7kVIXK4yKaFIr7PDVEFCCWqlfd7AenbAlYEKkFB0xOo8KBSrNthiDJ0nxguuZ2XXrwM2
M6ubJiwai+5a/3QKbWWKTZOmBL5xfe1pXV3hHUYHeJnSXapc5diUiDYvJcXExn/hOJVzvIXbTtFP
EugX9Eiv2uz0tUu9M2nHeiZBm2PmpD7vpraHePcHK7lp4c+5ywXo7o8WYmxtMKAXOs6Q+J7gjpe/
LtoFaPOC36NL8VWTndfeACeQvXwuaYM1un6aBXnWiIQFLndHFVidsTzeiIvMxk85Rvfg/XszJPlj
riuPCbrM+Lqgkl7kdRzt2IzNp6vvZyqZFMN5fXZ/74ZG6Z3gIe5Nr1wEg1SaKa2b42geod+BM6s+
OodJWXS4YcyzFH7MXvz4gSJt6mRZfQixyL/PyTyo3k937xVy9Mz4zy/yesjNA9iCTXW5M4uGdb4m
xZHwSuxE+PX3vUWQIP+dwLFyCviL1bL4E2mXu4lD1DM/Q9aJgFj6kr961LnpzaUmf7kkUpPUoeew
ZPUedAZIBOuJtaq9pysJnTtKh1SisiE0UN/GIhSBaZjp3vH4RxXDa1vYhV4rbgFTcyQw8gID0u/h
MHnyycsT8i0xL+A14tvH7kct3qIvvcyNrSrzq02HGQ86aqOYUP9DYqZCAKhLgxg0EHyslcy8DZJG
v/07yzxHFW+z2mdmhy1vFh0upKsjk4sWrU5/aNkKnNTYg+nO3fvgvqXsOs7VTVTajg4Jmi95uaeE
DZGoGiVvt6pdEByUqHnz9zXpzQhlrYaBLdGam5vqeJCjcbNgOZZ69vlr1n2k1LfSZmM+Ttcgg1Xr
3vubNIw3sOGc7n+lf9U0U5Bog8jtQ7I1Mz8mQLY3iA/eEaknXJGZ6Udry7X2jKhNzfeCNmtver22
tc4QF/XP13dFVMo+mlupQv+UPjO8PMEEIkdBvBWcMpZ31DQUvbm2H9/u/DinqUX3HH9gcPn5035J
vo3xOaVyXg11Pla2wZlScdUq98zTatisOE6V3vkTPT/Nd+69oMWYOZU4l5PGYjQwKyVRLciBnnAh
3rvxEgDKQ9VXUxoEVw9JjKwh3kLlOB6Z7Zf/+MN0eLxUlIAqg7RJKDQ36J9rfi2omMvuV8YGobSO
2Bv8luZNeiLRYwPHysy/GMTgoHy/ZNc+IdEJJUNV3mV5ZUs4uxPpqne5SgbBpKC1kfKScvWG+jz0
4L/A1PCucxTGveCPQ1zOg+l5z7jlKpD+YmAazAXgKAQo4mKYX5QaO5bcZgmfeQwvK8LNgihvHPDK
wrHBQEdX0iza5RHqbi6Je0vDSkTQKx6w3oVaxAarQOBEzJ0Ru8tP1G8jHOKefORsDaeeHXYpYWFH
0F2ZVO26lXspBsrcLmiEQwgEYc/k06xZZSSlZTTzU/8UXH5CQIrdfi4kGFpBidPnhewdrXnLTJkD
eJYKB8okxE0aIR4mqpGxrNJVBGCE6gfRf6G3LJWJ5OQ8aFFGd4rQDvnVfVPH+HJVzZ7llJtdECrG
/cvbXUA996YM2ovAFRGjD8zt0gUV/DkKAQNv+nE8UIn3dPKbbX3PevIRHoeGlyItjH1r8A2Lk1WW
A2hfSaTZFSJSTp7cjD1QRC/I9iqjkbSkzjjr93iOC7qSjlCxLgHTZzCoM3toHzQAf+OilpKDhPpR
QKV7Lzq/2iPpPhFSPSAUGzvf23pMi53WmJp2smFmxdC+4Y7SOUKo2dMHbjkTI1IrnQAw/pski4EG
7NI8rqpePLa4RMkv688U01DuYDnOtliPIuv0itLQKbnrhV9l6GW5sNkWdWRnIN6MOUlodO/UrpXs
4OFARw6WJlFTk1pj76QHMqbSQskxqZW5EAsW+kRWXJFh00Eb5Kc3ry0HNanM6LjXbnQpVqriBuF6
aerE2py8T39rRdlv9tNnTXS2sjre0oP+G3xV+rIl+ThLG9aZ4nbYTEhwJ10UebG1po31F+GFFtia
/rK2b23qSuFX76Uui6LvILrYCe8Hgo0E3iwu42fbsveGnz8mKmrrMapTLzptd3UbU0kSLbc97aOa
tyjeozhVWVhW8INUx5K41OTXKFKgikqXH28dw8dmnAVwsLh0Qe33pHURjeQ/eL+dq0ydf56UWwV+
Cf0JX04afq60uoIOaeP1Kt43xmnmh4lAZgGqp8tbYnjZQKJyJzvr5jRJT4n2Z2RRcRGhVSFh6ynn
yCsAmDzdnDaJ5mPlMSLuoAle3b1Hmr50Jmk+CCjB773DgsO5QuRD595943cImAzd1v6A3XG6QdJ3
R9ETxteypYXr7aOj99a+qG72FGh3FQjAGvdqaJBfu7dA2NMqf9f82DE9G+YeHMFu02x6w/tiFK6L
B8fWxEjCgZd+3DGljtO6BDknBG2pUxf4wIincB3S/DsDcp3WPxdSsPMy8+NlMeAA8XMm48gEQXv+
57QwRslW+CK+IoxshIdomcPmX36Flye0BzXpqKAJxVauawKE4tYiLlfPQxQRNkgD5ifhA/5KzNQn
fvOZfJvdGIL0u+H2Gko636CuqKncHB6TMBjTGtFtU7mfaY66Lgwr5fcAzj5dwFk5hBoSGEIiK8hl
HrJDAM8BfwTuwMT6NVlWkapKxtH+pn9Xx3y5aqVKSbMvqEIxc2ndjOJyv283MD3FpchaE4dLfAms
X9JG8UgIjUuFCehc0vXR80QabOujRsbK4q88mnjbK/avt+R+d2RjPX5Dn5DZPP9rFdnXm8O/TVob
i4ZsgnT5wzQgzG6SrD5vmUbgM4RLw4fv6pC/UalgZYp5WXXu1UY8reicpbwrum9V/SwjxYfwTsmA
35vXSermGzNVfATZ7idDZf1EgK9opBSTzP9qbFz8MbX+QfIfs2WHoJlnTTxCUXCrNNXi/alq+y4k
cMq0VHBYHx5Prb8xqJm9NbMwx9JJSTLVuNKTB0DuZ8h7yClG/qJ2ph4TcWJY7JcZuzjwJhWy0W+R
2MM2p1+9EFgg6mbK9RBss2I+1EIHiYfIXgfe7ESakxnO9HgvVEv/wV7bOrQRzBSUa7Sic1ulcGdW
WOJlZtKW92qBwp5hyHhI/3Y/bfqdbo/Alzx9CahzIEkMavJSMrKj+pLCqok3AKWQZsyUvPYhAxoV
ILFG1Mj460u8wT7Jlo9xa8N4mh7qTU/gS+Xju12RxNUFwucEBpkatRmpgZk3srbLn2sCGPfPwm6c
RiDYGgV+5xQwn5nyCnkGXlnnMsdVIu8n633pF2swx+4YEeLUb8BIct1OL+CvbOwuPQRdXELzMR1I
Z+vZpiPFkuAb+ope6TfVy8Usf/7C4sEBtgvkOKIgtjUFwlNZHz/srR8ve0ADF8cTfAyhq85ovnwy
sV0xCcC5VrzK1IXYK3cSVoeQVKXrYv7llPVnxe7okvxS7G5fUUJtvfZ0rgrj0YRBNMezahIGSmOd
cfiYOU9p2xy5xmfLZoR+k9ORNqlVxhkrydlgr4DyWqQoo3pQlX1veEaaNlUHjnnkkuALTuEkQDOk
J+PNxw/iCFRuyokO65jW2uQ9l0g19rYY6/hAuZ00cm99coPCxIqX0mZI/ofqMFt2ae2ympPqFARW
gdnEcHQ00LlxXV/PHvAx+OGqfMUbS3O4DXUb0eTgu8U/S4VpryRz52zM1wK7KU794cMr3Hs2V3Wl
UJ63W/cElSfP9PAjUeslrdkJgIg7Co5B4aCkhg/RPWgwfvJM50yTPlYP7Y4Z42Sx6+ysp9HHsklI
7g4pMvy+UF/WAsvmBwh3T54d+fERQzal5Qz6Ik2o/jAoa6RSYEF28dri6CvSPNL2Sbhp4vAExn72
rPdp+LGWooYZ/jQ2NTN0Cn9rmwbqTdn2lETRL0nYVL6cYSZL0Vc2Rdo+/n6r6IMWmlT9Bl2aJVyI
A7exXR+wuGc5tXzA8nsaRbcD4b4xj0bmnKVu0N4DYJuqGYycxoDtZU6Zp4TZSURq09sFvfKQM5na
xK4AKOdLL+qIOfVjh0ZkYGNBbj0sSK4U+zM2hKfBxppewpIjEC9LFu+xlY1ivQqPGhwC7frZqGKg
VX4r9sboPMiQ52LRZh+xV0ZCBVyOwFF1uxZLo8HTx7sd77LWjgK7QmqNF/omryWID+qe1S9OMAO9
xt2ZO6UspiD+LdHSq6g7JHxqGx+g7AmgLsSPtlk4Kaf/KIBB76W4oSrw4SFm56SioekQQX6cJMGO
VKJ50En1sEDMlmdQIHRF8ypcpLVSKhEGz85iK3t2SETNxkskWiPpLR02bANfaDdeRLPzNUAYkt3q
76tnidmiMWBjCHUB2tY/oFZlpNdWNah4w/4NGuf4vi5+Yb0OeiqqcoIEWXbKes2Vo2UURc6Ha/Bn
bwcAUWthTqAkwzoEKZIIhhcTElclQDh6T858LDI8nf6hwb2NOWSipVSgl4mmZvswaXw9KcNB+D6X
HluLz/Il5VCIBGj9dWUJsD/mnjYjM5L182YzKKjPvc0eDLTKiYU8CYAHUGZsQIztj0q2ndTI8qd9
+sgbiKdXBvisd2dZg16DzxmUC5E21LGZMdCvDgGS3X5Wdtvdt3JJBfE3GodXyvrNzPJ8lo/T79OM
TaCu7njMoloKehFg6V4nKL/Xrzc+/mSyQf3DKetgbQvPy2kzphIjxjMhFgQiDgmBEij2Yxs7SUNn
fpK4CibkRdriq5ZmE/gB2jo9ULoL+8F6S42UwZNeZwOaWVAvkmqpEV8M4Z5klI1ji5MCI7PkMz46
y73urunH2SccMmDb7J7LXOAbogJ2gh/SSqxrxJbElgeNRiFxITYLR7lLuV4RdjYlb7mT3+4erJ4l
SkBPlbyB0g3DBfq277JKFZOpQs6qYUm/nVsfXnafyhcRLr3GYdftiR+I0JdYnMCruxvqiOWvUtAX
d1yuhR2cLGaWG6DWyrq3UkmbwcpL2kiLBCoztKsLS8gbqiPU6q0TE2mRrWqWTzvJ4CAOzzLVLy8Z
TZUuCFVmPB0lBgc+WGND1Hiaiss46n5G973Ec0Js/Da0dn1MAOH1w0XS0D76JX31NP4aY8STM6FV
OwJxzPTidVOFQwNOiZ/3mCFSXHqFYwIVfZiVVqP6NQA43mQDNvfGr3+GBTxLKcydpuoK/blo6lxl
srn7CdAfem57iq0sitvKU1ncKAMWt7cyUZhlL5DhhkBm9hz19yiRvfneQl+Rvl2ZU9aSA8QQKxyy
nuUk4rR+YeBnaWFFxSUFXUSO1RQ0K+KY9sh/SbOpJ9W/eRAVVPOvApoN6tIb6oBrPKY8WvG9IWpD
tmEpwATpKsSKY35Qci2z/Yb1DkcGZBItKOb0W978U9FkyzRiTJvPMBHZDJAeUFyPqplKmtN4pbIc
k3q/rynX6hgWayrQoa/nMtVVFZdFdcOKJ598GgU/vi44qQsEwVF5K87IkbMIjtcpNnt8GRF753oW
lcZeFPEVh4LGPJTu0GlxwHyMlgnsk63x5CJNjlsJPgzpoW5714AE5riQ2U1N9u3k5S8TZTlVqC+J
LzbQicAT2wSjQ8eZpcBfBmkE0/Oeb+CuHOjeoEX4s7xI1YB7DGSkjYj5evdlSeq891NanX0lkXCP
ZoYLvVVhbTYdJ+YUNQSglQ0EJS3+H1zA2MLgwqomIDv3C3SYJdPgkHGRj+xcphD6Vn9YiTrrgXj6
94XRi1s9PNoys6NzzHPiZKgNhZaDY9sN0SXrbj1ZpeRhrdfpMPA84D8NCDuG/rNwBA4XR3e8P2Wu
ChppoOZRdXobOtdgxkZohBjVeC9DqQDk/NHgFXZ1nVOjQgsZDmaLAU64Cbi6OamMM8UoOfme/Lnp
/8d2hFBOfN2JF3GLr3lS+PjknoDgd6NwYO6B2S7sqECEbGSxyctClvaSJfO+nQ7larMGQwMbaCXY
p7TYaYj55NYUTwEd7lyMtF0qrtVIk/O2NrPyt+KUFUL5XncbNjEjcFzW+HJHuxMgoy4MF99Ao0C4
A94j4fhe4KDL4h2AyDtPjwTmnWOfBJt0NJhSRYrTb8Skb2xI+CpHy5fR18RitvoH6WrfcUYlJtw1
m9WGoOJUUHckQUtI96qwKTakYuxBf7Lmzc9W02hx07O67l7+7dXbKfRRqnE0IcEaR/ur24SKbPI1
dNAFG0FCCPFUNDQcjJBuuR0CxaOAzWvTfW1zpgOnw0RMeqpqlSHbuJllmTliAuzGfO1fAv1YyD5l
E45F3tS2tCeuWwhySq5jA6LL6UEh/59ZQytW4EF6FSHnGYKz3Qx6DwNI0aR380YWS1Nx9eTLe5g/
YfP/4opn65bRNMzLPU+VPcNFAqUYxF2HzkACuPgfHc+as/J3yyxuCk/lWj/cFUTc47XBCwadR3hY
tYkVCsVah/Q5tLrM0F+ERW7beXks/Rl3U3zzf9yM7UebyGwF22FS/AIhJqFaB7MJFd8/9LVta9Hr
nU25jh+VyxVg43JmmroDa0KPueWGwME8o9Ep4TYSd1V8iGv+63kp/MjM4tPXdD6ecQdm1CGiQ3YU
6ZCFD86sf6lMq39TS4Dhl7/QgoBpXaKHLr1FryTtdl/idCHrfb2JBdNdYEAnfgduQU5xR998+mG3
SRqP0sbLvj9w/c6PI9Tf9XdQrxZXn8jNNvqik8dNlFyu5tWD9YmxwRrUS7UPN8XQKs0Vt4/izY7P
mARoRIosWKsdBvndmNEsYTY+MY3H2Vrazl8kWbitLW4WyNTLksTLGKB8Vs5Ju6Wonjn9QCuaJtDY
CnvrvWT3c/tZCgDCm7tMGdiJZ1/NC8An65JCWnmFxIn00KiTLR3c5oYd2ZqSvSZwyYMi0Z3bKT1J
NpnoM2+aTiMVzvxDW6iyS7WkHu2HXFRDTknJxCMWG0NnZbysHFCUBoc1OvvNxyu3bz2CbthlAzTj
yllCzucTBR2vq20Km8hN/+DC14mw3xpPKU7jX4MnP49+zAVs8n5Lb3J5jArKlutYIiYjZt4+4zsc
R/3lhB7MD6qAHDO6QeAGljipu+zvNgiRsywRDcEEMy2LrrjTSkfRVUBEdngzqx+IQOwqWox8Rn62
Ca4NEKBtVt4zak011dsSBQX8eBc/aN5LSNikoT5R3gEDoLhYRXVxMLz9WQqwFhFPsRP8lmFWRMTC
wHjmpB3np2i9XnZ06tuhL2/guVZGNHoFTq/jy0dL5vK2QKoaRVe6ZIDbb6dt2ExqgqnHst4BnIN9
VzsnNQciN15Kzkgmv94gWdVtYioZHcWLhYN3djHTqdtmkWreulywnpJN7D9SI9y1Q1HahS/ZB+lm
MQB1yyLvtjYs4GkeFKcjNVQmUCYBCmKW5XKOk4ftAz5vSKOqC3dU2NiD7EKde2/Q7yAltJ62Jam3
zp24Kyd5xNLq0uBd5CDnUSO7opjFonVa7cO94lwhlADvJgGmaeF9qdidBL8rx3k9Ponv1TTSH5Nh
sM6HubaXVCvF/2AhztneAZnzQG/5SBhonuUoIUbAAFAkE6pjL6GQ3u4XCiJE3p9Koat/iE+gwRfu
1Lgxm4FI/o8VEssyzI1L09ZiWpGoC2e68uJUHBbvSUad31mNH1/tRAGTYZzeZI7/2Qq34wYzcWOn
Mu7FLmPZj5kN2aGdvRSeb09W4FTKaL6Alaqt1/iBYNg7wJe1KPspZirkruypJiINKCmdAe9G/3wV
pqe3ZXCqRp4B/5Jv5thqw7yFgfcemT1ZWLUnpy0MZeiqPJXhC3Rhp73kCjs4ehfUmr2uvHM4hlct
uHl2eg/gvNen0FzIxnY8Fwx67wsCMTDfUsn9DA4Jn3jjepqWIzG3D6cfYdTRpC7hSGOPlcRfWKc/
M0SVBwUbUTVT4OzBtmA9ABT/lGR6RPRiZo8rkUXPE9JdYH+VeSrpM5oTQVZ6OV10RxWPip1ci6C3
gDD8/ZNsvLrhwmz0e4gck7XDy8r2oqmcOoL/DcNtXrxl+zltbvbdfYvTvTOdvTEC7GlGY20aHKJI
CCRfCnKT2/EOS/J+me6y4qXbloiRayKzLLkr0Q6Lg8EIf3DkaceevbUTCDiBaLD7F9jufYPXgU5X
BCtefauv/0SL6VCjVwh0XBaGPR2OpdVRd25yG9lHZbzYD9Pon8wrE3FGcVRcWMD0NN1DRSxmJDcg
lCqfaCwfABWihsc/ifGZXOct57ETIqQauIUy2N4aLrPo9jwTNGk6KZ9UpxoDQDP08AwnbrkacleS
fRltfBYRpo099mo8UwvyByrZuL9aDtAKPy2VFGC4hezM/NvHNT0bRkUisTIZXVl2j4qRJSfUACy4
nPka3mtMHxJSYVmTDgdrGIo/4HayPJLNeUxxSWDH7ltaASn7URJdCKv0q1TPctJXndbNPZl+xtKy
GlrcNc69qvQpb0e1rlxiyBvGHEUCip38CAdge7W8ZYKKQ5Lf5wrMTdaID/FX6lPqCZWpxeVhLAC7
lcrf85Os8InGc/kHC4bySLtT526UZY9gaLCZ/oM9IDS0rJIWhQ9PYvm8otq3GgSwxhJADiy1eriB
qhN4T89fST0QpLumvs51f1wicmPdocBWQL6d09spmi0Z/z6hHcSKntYl9Ec0HxGrUgbcjUq2F+hB
t/vkHTDVYiSTcNlal9PhEw8/G44L8clOzNzcZ7MDtuUPxd06YrHHc4hip0zkbRTWAb1yoLH0q1Le
Q6GeFGhd93R+jofRbd/fDXWgVgwvVBaDbktSuG1mIj5dnlA2tN+Dd1gRUSmdtA5HdcBww8cZ2bvl
vHk6gVGpxIfQBJ7ztl1t8NIDWP1FNmO26nYpIbiNXF9wee2d5jvKJ95XA+FME7Wr38nsYzoh7J0d
sfBs4kFTEmrgLT5dnJwF6+T3YYHpHr07ykk0xUIZ0lHTdoy6s2wefC4nZCCWBLSeIa13Pb9++cwu
urpzryFFaKpEWiQWPHijQ6jVfD4/p8DJDGNX3+0opKtxeZnrpXTi7AJhk54sMdWNjBf8MX/gEPDQ
M0/BCbVgU3uxsIFx3I1CSSk+QsjNuud6fwjzE9NheG7Bk2C6VnqH4+mvuMU0aInmoM9GRScTr0R8
jhG6mJCJs+jkB/q7GjXp8t/sAIQm59TOzqxezZJ+X7R2HQ650ac/HONdz8VnjLByhHLkon2zOKxt
bxTN8kYxwb3QcRPS2Bwx3urTsufleD2Lex7cEEf/qqNwELyG96tXjaNoXZZA9X1aAkmSr8GNnEAk
WF9mR1RxLjHEJtCOiDygkBuus1vk0oolucq3BQ+JhnRPqq9cJw9X/aOTDi0q+M5pP6XwZ8sZbf9X
gkEg4bWViSDQtRScp1wfCE5FQnxC6GcgGFxQRIJdMc2kM+Xb5RzGKyp9jWIwqu9S3tF3G9v63wrz
KOmX9PJWM+ZQPJkoQ/ZajxFJbQYozPDvVTRmxhF58apacSI/XOvQF1nvKZti/YAjirPnPsT8j2uO
kCGLRzmouQHCng9bjX2hLOukLq5CySFdtpe0LnFoSPeHhV+ySRxnXOVYd+S/ShJ1KoBdj4ZFS2Rt
8aQ0uF94BVgcJgA0oKdNvmlVRZVp/Lpiquw0owzTojpBO2SZn8o5h1hu2bUReZiSzMFxzdz2Bplc
55L8ZI6jYuC5akbDPGPXuT56xnIxeIx/VnlunOyAFp/Gny770iliBAzXsswKiDWgiIHT67J5ZT5J
3teAFtTLnY7WKruG3xOLq+J9BWjKtlRToj6RTEf///RGuaPtl3MiBepU85zGjSNBRK7y4yN/V6KB
PpwXl9gDTaLEKGhtY7WhYaK2vAThfL/5I4nvDk0Cw2Q6SLq+Ufw94SWZnstQ5x30SmomFe0QOuIu
o9RjRtGSYj0FDYZltGTM7qLa7ibVjfsFDT9svvkWAJJVc80Q6y0TdziMnxCmNc8qcYklOiiVU2rD
rvCC6iuveJYjOEr4cGoLLA3bO3+Q7DkGokYFiJ9gICNMfSqRe8pzMiN1yXVLwPD6ASmK3MVCEvZt
jpxawyAD9fNTuEi4OgAWBMPhfuXeNKRnEKrwDh5x0CbAtRiJlMHoBPynv6ZalCgeQwK67ZEgRqm1
vSPbYTobi4AXfXXMp2J+SB5TqdAYm75lYLF7BfnmNfhyzzR7JnhbpAcquiNrbtDL/6ZTlaBfpY3N
CTLo69zOggqXzlgpWEvcdjuTmDzKHvWr0ohXjjOl+arilkpu1k9/ZbftuMS6jj1BsxvwmjIclJbu
KJB5LzzBVfwzR/qFIqKjz67x8/vFKxPuaT7/3mTLPhqSpbDa1Wewmf+LxY8jwnXjBHKF8QsVblEa
d1NbWM6RzZhmQkDVcHZYaRlwaNFvz0/u6PO7oP1jWmRr49bXnzDmT++4ABsP+VNUBJVq8+CRHDNl
nmqi3gXRBTzEyAjZX3zS/1/tTOXslopifsBBIq3i9qONPsGN67l3JPRboQJy+x457i/mTTugDYRs
EdMQX9Kg8kxj+o2ACEEjiv8Mgs62iblPrceCjuqQioHmW4BKYPT/RsIVDq59TPVdlcl0XkqfiMty
24lRIYX+R3b7h5vScFtP0wzjeKWqjkxLk9OSu6TdNUZGVrAmTPw4HmLByk8dwTexyLNbNucWsxAz
u6XGTEd55vQlWs6OtvVAnlgLfLy2nnYq0HTfuS9LSY7g5fkRmDvC5ti2O6pd11sqjLhXQI9A7/5m
IhqeZ806TfHO0/B9iMcxdHdhg56Im09Jv7kCTrVsTZMBOlU/kAYyiYQ5VlEjntkYVqZ4SOsMdI3M
c3j/nPpmtuxduFX1Kjn4kPVS52Av4OvrKianICHGC4kbzjB/1jZaGMsTfEj4Rl9yc/M8uu/cPmNr
HAyICpAKsoE+DQ2M2r0wxOUY8idXSWZT4KJotUOr3SB35q5Jhs6njcukAjO+/KZjCNcraU6nT3UB
0gcDxUmwhwCVBRTkfFsbTVNH4myhKI4NuZK7pcQzlHd9DxhaBeECRDmmEHD7NBG/F6HoRorWvJxq
CSMRXJKjl/ait20Y/4FbSRUNKyXiYdE4lzCaS36CM9rmQW0du/S4AXCujRE03vJ/a+NQhCIPsMDV
kH6nVhDys08V8E386Sk+nAO4+5HbeTVdk01hg8XmHlIizJhs6RUmvAQg5M79N8oRKY5iRQMuwxlT
lghrc9lBPmr5F2F+Fnr/VRnqyUZNONb4Obuv4ddqMn4KAxEUDyqXdZYhbwOhgBhxWmtVzXY+h7VD
QqJnmUync1G1o+VFM7lLurO6Vej/SaDiTlx+ndX1IiQRJTRkFpYsVN7LyO2S2Ywao9mP8uWAbXd8
RLgPzy06+Yvns8jszf83henVem0DvY+lWwcoubFBnlq98Yc0QtMKKBy8QezzmjnHwnvTV+l7nhVJ
fNvZKJJciRdlB+LNHJbEWxQ3V3c90alr+tZeD7ttYP9OCeR7DcIc2Hh2HyIG7gbGQhY22GW0shM+
0uLN38ZSOIcuXT8E/MydVNQ8PTO20GmvGxEdQhOwTniT+bCYwA0N4sVZzcbk0BgY2p2wMcO0iTMP
udNB5MrBMC7WaR2y6iKrn1EKewP7PQCvWsi9WSJqEqXt6gQK1GHpRBOQofAgvx8KjYKsIT0/dMQ9
NEdwCjRlN5fPlul+Kwj/G9Iyz1DIp+4UiVVsT2IQDxRSf0m3UdCbSN2V61+ItK7kWKE73FT9yjhz
PwbfGPcT/wOpDT3BsP0Whq5IjhjiTPcnUR4o4ll+NpEOe2q+tHgBczwEpADJcCE95powbUwNwiLn
UQT9HEgeX9wyfNxVxB/Y97ddBGVg9K/bOGIssx1XA9IKhZ1IoQ4D4SsEhYPrOkSDzXcLhoPX1rgF
rxvohgNu0T9d6yy8WFXhwK6J3YORhTs98nzmVtMWITzr+oFOA7DDavZe7Wo4oQoVpg0c8sn9arY4
908sTt9kSZPChpC13mR9E1oDvvGIlJaRPodK6F2wFduif77qtffKLYxp0p8U96pvbtdOQh8arY7m
T2QHDzZGKRmpaMmEsJ1pYVkGSq6QI6l+ZFwO2+EUPpRkIb2x7++zv04qiWbzkmJyr+PtVK2AXJNY
HA8mBudrYNMqRCHV+lQq5U1dvJb8ew7df+EI8kkC7DVvh6vLp5XW01q/whZQ1q/s/SDOCP5mkz7i
zNqeZ0nkxiVsH9ZQr/m/xt75VWluyAdy3BZfIV+2XB5hsJyKCchAaP+dw3yvzH260katBAM9aNhO
mzVJuDyYPX6mGca14NVhVVu/GpSrjdpifyxckglzsufSmFK5nTdTJDL0ic2gxSw+p2nAN8O5CZ7x
eBWQUu0eGRX41dYiRm/tKKBCaM51Fdm8S3EGBgnTklh4J6Ki1aCPfNuqr7GbEBi6CnIXkUrJsP9b
zrWby/JkH+a9vDs9qlNU8AGlkScz4nu03nmbDWnQsmgg65wnoyrY+Q70oYIa775iQXSaQG/wqJ56
RaaNSP2dORH1tJ+g45Y0Ji23Bvbap59Rx2szfTfcGmK1GHlGnAypYlYnn4fgKUtW7dx4AmAUlxTq
ybtbOaZHANJAR03O3nGeQ33MdgS/ghPdiRI/9mpULpRn9jTSer+gk3AlEbfoOGgMt/ND7sxJWyEU
1443flNYF4jSs3mvkEW03ILew9LpN1pz1+pVfzb5M8zL1I+L6D0ab3sdoKBjAhR49b0nkM0BTyIq
50RFWzIHfCJbUvRzVCCvDSzf2XTa9JBEObxfXFtlyvdwVCdmGh92LnviD7tncQHUhST063a9eUwx
Jy0o7s8M/mI2t4papNU4ObqctkiQ/VzvSumHbGWwlT3iQ1V2YZBeesKhJxXAITFid1VJBvDERL+O
/NOq6SjY+iIQu4uFEypAp+A9CrsmfgTbeun3UgBE0z2B70utigIPMEDdrh395ffUxP09Lfq7OWFO
MMOWu2hYh+sEe51rI8Jbpc/ghBvQMAdIhh9dw1IuOyl0+6twMntoknsJp+kMmchIPE+uF9+eaxjx
fOLBFYQpeMsZjTaP5BWx9c1vSWzNEoJ3WmgeW5KNmXRIv8BrXfGSMk7DEQP4ollw9ncXW3/RFau+
GbYWHuTudTTFdvufePYgPapfXtqrtfRpgUkuufw8Lc5ZdryMN/OkDyzUuMsXWjfolA99yrzR21we
ZgDAN/TuIQFZgJwMCm4d+qaXfDbjowEac4RcWPaNjdMbYNs4X1jZXwlzwlaCpJc3XpztwzAu4NMH
9EuScTvOlECkebYTMorFBIZvAtdIb33BXEurw3O5SWuLYVWyMXiJcVN5YX+xK1cKqDjMY6HdEaOG
AHfPdcw+O9y4WWVPxhtwQpfD2AswrKJu7LRp825g5tAN4Jzf6Di5V1a7lk8PSOKZyFkZCqoe1I2x
QhNmJU3osrZowMXjhgwldJbWqFw2mY/6qzxhrFY9bI5u2CZz/tUNmJQX/D/ESzR2L5wieA8M1ZEB
fd1m/cTMT0ogb6lO2uVQjGGXM6ToDn2QuMgfeIvylCNNpEyPxp4KB+vkjm51LE6CIX0WoukOI0iR
WsB6V6qKbzOqNuGTCHW3/DeU+1uL+BbmLyEAIbv8771jEMtC3Sw6imcbS98f/ij8HPs1ClgcnQIL
+OCpdfELvzvbQq8eaQfpROTTG9B0M/7X/6MCS4ksCwo58GI16qSZPc+0baMhtV7igYy2PrJCfJDu
DeQsDSZBiSiH4PJrXtYXOZVRes4G4w0pgUtstsj5FnLKSuV8iOPlXmXZWEi82B/PGQSlD4G32ytX
TY8t5jyMNNQrUFlpaOZXnuXlAozowH0omR/XzKtNE/LXQpXkSZN6nliPULgwea2zoe3Np2CxBqu+
6GVqTvUMRmT/54xDX73f4YIt0fxKZukFWsMAcloFksR6uo3Yh+7iF7xlVTEvl1IRbzrj45q9qAyX
Xx+2q9HHEcVHpq2tVZXqKfRITkyanMhP/PSknaYBj6ACxLndz8kgl7JSGPWN1Qi/WsVnQOAPRPGU
iusIMfadLpoxcXXWSbpimSW+7BYfAV9ntzLTW4i6tvFeHYAzfMwL5KDL/1GUoq2Ut0XDfpy+lODS
95KeT8DPolGv5zHrEARZIFfvIuAAzBGecJse1GcG3osr1ZZ9S68LDJts9TjVBVljxLKMmemXnk+L
yYv5yWivw/hT5WG61GaH/lP77Sttzs+DHklzB4jFMlWQpdnhvcFuqAjBYii9jWyLDrQKnl4+JlW3
qf6yus6uxVxVGYOXnPCxcObf17blcqJIDB7GZP/XXIeysogtTPgVkdzwaqMytrIEzKyRILxmwAJ0
gji3oFggwVT+Yy43rtIYkWFrYRNuFfBpMIKbjzvZFdVMKFtKfjI1h8hunsXC3oop4LrFewMOM2wu
fLCZ378Vpp1aDg7Opx+YmCZzy3m9xultBIfxHz8okBqa5wIEH/fXmUhR/vFk+GFRHckqEbXaNi0y
s23kam+i8z9XlZjVOK2ah+SIPFai4r8G0arVUqu1/4hPv/iVcfDeWwgxg9+VgJVRlyN2rTj47ypD
jPC9Y7NWIvmIwSBc4mzD2PmGVQTXrn8sCbEq2c0R2kjngsHA57LY7fif8sObNLsvs0rGCRwttzMl
C+amnL76/ASLJMGpqNrN/KSgyMnQ7uRc3TlHLxqH6Fdqm7R1ej4KRKJXt19IaJlbfJRSl5gm2g7J
6oj3esWw85FpP//QaUmCP+Wb3bW1KxEutxfx7bZxsvZxEsWsBvA3t0ivEpbCGShdqese3UfANKL3
+8B7Gnf0vdW0Yqop2EGXF67PC/5B3m0puvQpfxMAiQ0Is9DMeBYYBaENJEr6rIahtOltBx2L+ZVq
PMOM+Bbmr7ntrr9VPasbVq1la3q6RRisHAg0xCGvPPGdABnjzSPqCL+cElkEDWZ9XaHuBJJGMZPe
0DK7kO37Pdh/e2/rbrp1o3kJaSpLMLUVDa6FBVvpTVZJiJv3L9Xzk7sR2bmmg6uGB3EmztharGay
Q64I+b7Lk+a9tM9X+rc8VjXAmiZbws/Y9w6j1QpvHEVQhvfsOBPpeOV6KDcAwtura0XUc4fG2Qfk
34ipki0iKK0VWK5xC6PrEZN6iUCzC0rj92ItpXJrIFGmcPLjeU160AsA/lfiF8VJqsttKltqr1Pj
0QoZwxms0urg2zZ/SINfCvHYcXWSPOOTU+Sc/HF039vwIJAvDWFmn5jKr6EtRou5mYtIo7r9tWVA
Swr4cucMjawLP6WACmQLArPPa7lcpnkEua27yKfAONv8RuWpmYYwdQxlYOEc5ykAsyrjO2dzSMWN
zi8FySASz3AtS4jcqjya1JdjHrRa9sYUwR5ajeIARKa5COCY/QB2hqcCowbDWVHD4352lyBz0T42
Am3g/B4SSPpZbtVipBe2wXPj1sqS1Mf46NDhzRb6Echuz3c9zLqo0cqBQo/dBd+EN2qkoCXbAiqn
9GtkclHdygPj/asEbtueBZjlTeE8JeoH9dGNScESg0MUF2Wfc3ZBJCsV4ARKrTZt4qHjE3oB9Jks
/4A2zzfBZhKMyDldeVVc0wZYN4VOnfdqXD5+yTtBSlElCqKFIInlLsteE/gqnEW1ZANJvjiX97Dc
ghanDNab8z+/VkOZg8IRVsWUBmdOctoLrFi1/SyyUJzqEIUgf54dI8S35dLXTNkEPSYZ8ZX3BJhk
jvD3NJP00mRCF1+e3dg3pP8ismeW52ij+YWT6GUKPo4cjQ2c03XktWGgrA0vhHeIXoAuD2QH5NbR
8tZ0ZK5iJJ7Pzb7u8Jy5Gtn4Sp2nXbMevxfDbFUfsyxitOG2SPvGkwx1Eex12vGVy4Kxoy+g7m3v
R60rAXoLf5GrXWYTLiF3kL0yCdGUNl0NBUb/OuHqZGtlAY+PPqAzUhhH3RCht7oTT8/GtUw9plXy
PNqPwBWPGrR1QPwi1goBTwz4a8VHoljmGoCX74WEOoboM4t8tOefjBPPZWwqGDI/Bez8GnmwQXaf
T3egkt8oWsoRfroxop2dBsptswCw8bHznFbQ+5eoUvDNXrTBqLTbLruuI2S23xMi3MSOCZEEIFQo
FJu9eQhGqwa11CqxxcxfotBD3TddcTkmsCWXoZPEwDZDc3Opw8vhc0PYUmJpEvOd47taZxxBYaEv
PYSe+ABU1b07FrUWG7IhmCrkeFnrZcj2ABxorcoznHbk2qUSvFxHzUlsWp5jCqODQaKB51BKwDBg
D2Kzcm14SW3MHxssUsRphHf96q+zdrvfKV3G+DnR9BS41yKur1lXSv9u03YoiS8CtrruePAoDzXF
KlqVU13mZ1cqSAKPtJfH7bRsKUOh7vA1lPgDUqjSzY/obytq/WOOZ2kmtYG0B+S0wX2r8HI5PY5D
lV+IKFG5ghqCnDuOM0R6jZs63TGN9EoAGMbud3J0TI81Gh8YDvbdSSC2XYC5VgcImr0nmPQQzH1J
BRoO6aEuVsuxsQstUu9M1g20H7xIirZuUiZJvv6st3eEEXE70cI65POK1T2EflPOn3BoGpl9ku5D
CfSLu97TnTvzD/qtOCHWE7dsYtGZeOiT37eoY5G3CNhPVRqLswiLNHCC7BciAqFXXnF48Flkxwer
MvIT+X9EzalHrwoia8YMmtNqCrTwBvurprOoP9aWbSu4aFKk8HebFcIcqUJGzxBguql14+KSwaK2
dJZzSbRX29LO+z9sHjcxY2+nIB+0kopdDioRyBvXA9CXnAtt19U8k994pH72EiK+huzO6ZRk3jTq
lB8EczpNnDnQMoPw6/XWTRozHVU1+ZtpJaJI/qjd/s2QqlfTF43aada1Zwz7gmEGRWsZLnayIVxe
UjGHjFS/rQrZ9f6DhtWhLCQAaLOy5M0+oaVESzJRgNlddIeYRZpeQbFQnvc9TkmbUvjFwTPIBJ1/
JQgBb0ufEdtxl/RxN/r7GSq0j4ealF4ENxT941z6Xmu1375ou0uAnHH7ZrmsiuJbnG3cX8jrYo0k
mheVKi4AHKRd45n3ReDOR89wnRsRo/ZrgjmEW5weeRUnDaiwDcjmFjkLwWVMCrXpBBKrmxLU6mXe
ctg9WDoVRJOD+cWLQ9e/e+KIYee4C4O4ynPS/dTWkhsEVyibmDto8uzw+hf1zY0Xv2aTW+Fsf5AV
8WNaC8TwLklnfEGFpbSkOelh7QKTrw6WaiHCdLIu4d3mdszGf5sew3p2SQu8yHbOKrq3ih0hyuiM
P+/HMk6h+mPZtPF+4UYNlX797N8qUYECf1/8vMszDT7FRw4pOK64/r4LleoN08pd/NkdVTem3LeJ
NezX1ksFyGiF2f3ygvhAmM2e7vNmbw35Ay0x/7hrxDywHbQaJFPfm5x2saZjvQpWJuzAzdT08drf
vsSCZAoaBiRH1SMOf/Ijcmr1K3BjVyfoaZoj7jBFObCMY2/nI291vE5uKAsb2m8faO1HlJJGRktY
kVEAa2/VApDnIrdSZddD0aNwaWS5e/YncCNecjXPvz5Kq4yL6Sg+cNTGeLhFQa2mi7mc4c28XufE
X3dsTfHt2/HM/KSbR/GZK54GzJ6+B1qH4TsHt0XWpQYP/jEUj+Sna4nTdL731J6ZKIBEUtE/I3Xo
gY21KXrBEyVdvdv959xjGn5FtUJIEGNUe4ywtblR9mICnUeZ68mlcy7S/1v2QYcCjK8PfES89Q2e
7FQA8p4C5pdeWj1crQVgOm7vW0eLY6d0ifrDANAM4XgwY7iWsJbb76E04MDoFnm6Xjq4RWCW4USS
qzTjnAaa50X/iA0sXvborDkPN5L6+5bamLsbh2gFax9O00j7+Y0MB4yTY1x9RhQdr5F75+Kd3nlA
7bdBGVcliW5z6M4ht2mlDNNbdmWNWblD/NB6Ehq1xe2XbYkHRVNIcgfH6kXvv/tg9tyP6HgU7Xwk
X7RKta9WtEqe98DvxwwA5urdKqZJhwPbgWCogbIxcElX8IlAAaNvMhKXrJp6ZftZMrPLG905Y68+
PN+fS2MvywCMlZyKywY87VP8FI4w4l9se9jCe4OpbuoOyVgOtiEQgAucytrbPz2PPTx71G1WThxH
Pjh2SkxDTG0qIoMjOGXbTek6EKq8WHLclkviKumIjSYRDU92bxzWNAkMQHbRW/lDy5BVam+c5Q0m
ARFOUHsarGoQ05YOflCaqoilJwR2A6meIufKsu/ZhUoJBZSqAjmMrs1IdfKhetK3079ss5UAGC3A
NPTYRO1L7zNXvh4iTjx/9ziIPNHWLJUAtTnoUbFlYCWOVlRT0JsFu45srpDcUneGgchrDkxNqsep
dMYizMI+EztEvA6m4r/jrqzkWkFg5+YckARTntGTtaTQWA+jaIeBB+BNhjq9GSw3t5g8Ng8ZYDdb
Wr87ioZ2D+XMKP93zS1nqORvcwy+yEC2IleqKcQfolsYVRqoffbJEgoMVowX8mDczKezHyl8mKlR
Va1nssW42uMZofv3BhdrpA9xDs+N4tW/ajein10LSfq5m09MKAbTO36GuCuGDeUObNceojNydg4a
BOpFLruwd/2UrSdvVcEMeV1cbHn7Az/5h+2ofZR1ffDACvZTH+JDNA4G3PBWe5tsLtOPM8u8O911
OFxH7a8/nZFNM1nvmcLiIQy8dIf84rnzrBE/O5Cffoyebjyb01cY1l4Iy7myxGc1vTGB+LUKEEsY
54E61uLnCIYPB3e7n3EiND/LLeORU5Xip3TftxiAyNhDU1RiHs9wpbOaDNhHh+24hsXeFnopGQRg
EiV0Iex0atnFzlGYcsNieLX8lYLDPAtO/inUwM1o8CCNCwWGmi7PyGtZw1agIRaDvBpKDcUPJ1n0
iO5Fi67uSDvSTYQI14wKqsWvfkSmFAtJq4rpb1NnU9cUr+u5U0EVYV824MjY+U/L8K+n0HKmrdaF
4cAVAuLZ5okLs8kaOSW/uErg2tsHd95giwyf+m7tAdQ/t+vgyQnN2Ml0/BCiiT68av8nILu1Cay6
dTSzohhQ5rx2HazNfo5urFvSW4D0MO7EbqFjdhsoDOHgAfdQuCAMvlgjj7kAtSRmU3WzJzWmtXHJ
0/fCLgwFfC6/IVPwXb4gj/o35zaEcMzEeXVZGiIXoDzBd/s2Z+F9qnAJpzJ8c9bKVDC/12HGo3cC
OeDjeg2q9rL0FI15H/oOw+IhFaj0T+aXmA9Eun6rrG3UPZU2TGMeHyLhNggfbQvNuFptBAsINbSB
yqRGUQtTKcseb4Wq2BTxQ+EicJi0FQoBsWX+7Zf3DRW/Wcurgl3y7Apy3CKC3YwHzSusPPjwfWty
Oqvo/R7ayzpPmy8MCEKe0aOsSesn7btgHlCQBgQsd0lcBepaSH2wEKWjE2huP62W2J8alMJVFnhQ
yVRuhd9XpoObrWwtsU+V2foRVAJKaWML9qGfVFckiKLCoVEbfBWUce4B+qAxugoKQpVDxEAGs+hS
YzO1C+fi4f070v/DehRRr7DcYWremwYY+hV0lgRudJNw2a8P7nUcp13A2y3acGEOgyKcDgBXJrMn
Ed8KYY7P0Zg3FexggUPI/9gYfLVY0IkF9sBuzYo37xG41MqjdLMbEsr7AF++sWG6Tke3vSVIQYoL
YUC3knganKS+h5UNd3sOqxPHf5FQoySEAE/NwAd7M6xfejgVceegaDHZ7A55zASLiXVAOGxQtpS4
Y4d/3S19Zh5LhlJP53BWXNks0sNue4XxAc1k+SrV5OqtbIg+xHObKqt3K/GNb7nhsdBOrbA0nL4g
SUjq4nAqZSczDJoXbte2ITNwrPGnL741iDGU6CaEdjgQw3KD9FoKP+RfythH7i+gw4peboJFk+XI
peNoyJevkAkCJz7f0/h2ToL5CBjdQgqpjglfJldmVQO0wAw714c4FjmXryTyEoHOQ692NYDVTZ4w
Jf1H1BheMV4+2m+mLtDw28KaMvX91sJAoNSw01NLnys2rIWavkut1pxIkrLlGVSgNkeSlz81bQDS
LXeStXpabuB4Q7JBxrT00vBLrrBo9FgQqTW0FlwHPEhfPom6amsWRVzZ4Y0eUKPiXESIjdGVg40i
FKhMMB5MPZS+Mxjhp2b3TCkVQyKqTuoPff9+VVQHTGpEVFcJ4SMKJL/bscz/dfu6tN1MmoAywB/w
hN/OnAqUvJ3zaUbVrhYmBzZpNvcH2pTUp7g4It5nXsKLdD69ux/ViCuITI2yG30Mr22WEpyk5hRl
vF1CkCLbJwR3AyuQXED7ITfVAhSt7bfQ/TDDgHSabu83uMLDXWqkqPhnMRaCuHjfSHWroKniatS4
MRZMWX91LvUVKGX/1FDZOyA0CvYypYogHodQiyzkZo/YRrGrqeAvAjUILDvwSyzcSz8ie0c76/y7
L8YtkXy94Mj0U/wFHqZCVKx5cZQ0O030jo3RQk4bxMrfcoxmyrq3UGdV5u+9DQkmZXMeFT/S0fhW
eSwf2JIP4BQ83KaUmrcLnolD028UKsy15XRUovnp7iFmETMtFlBhzncny5dcH/KQaaYsAOfWkR66
S5r5N/zABsvCcZwen2k/h/P5JqaN+nvr/GQxx3WnRU81tuqqWZ+538QUEaYmLpeE/BTJ69PGj8EC
Jd6yao1rmE+h3mcBkjsdQ1QLXI8pH1izcEGd9oU53pa+2/BqKRHKGIcchKQxfa/IoN23HjfjnY1A
NznBng7+umXxn7Jcm0PSW0Ejd0+gMLGT04NKl/k0PK5dPvGOU69ED1IqnEk1xSSPMbkpX+IWkNHp
inhpBp3RQ9KX1rwV2+0P95xSNZrSxmH7IeUBvm7VkCdNybjOn5Gp9T8ocEcZMPPYTmMSZUWmS6co
9Bfp6U80IRzZxtaDxnBtZu0ldGSjrdrPRC3EoVpHGb9geA8GT2qZEuJ6gapt9lcgn4EgheoxH9hn
Z5oZEFZf4S8a6XFkgM6EwLWfLyb6yg2ovo6MxfuM9TQHMWeEu0lEF//FCgHVb4IQFwNG72STKG33
wB9pbGlaf7KSu2jA/k25u4A9CvcDnQ1NGfyJ7rDz/nF1wNOHaJUWlFM5cjEYCw6OcnFfqSMMYtei
g9pccvoMDNgC16xkzzA1v6nuue2WJohf9JopHvBZPs/nicKUbB9H3Agyy68s2qWzhoYGX4GP51I9
dCch/i7RDrNRjbdnwkQbYtLuUfxWZF+7ovZT159T4oLWDvkVV2UsCI0qGWha7AaMFSCrKy+RAbk6
Rdqxplazt0kxeOfVA9+majKxWgUJDPqUYzpNz7Myt7bDMo1Mv5bHlbeYrx0aUcg2pEf1v6PeU0Io
j2Duv3qkkoFrVyrS0YINH+VUU+ZAF/G+x1asCtrM9TycHIwh1PGrneWiGDYcVfzWSc4+8ayZfP3H
rqe72ToWyTfk1frRCq+HMbehUu1JgD1asru2rVnNv16EhoK6cCkbtMhjjBGQWstAeZdJS1oHcaIY
K2Oh84yhkW00tJ4LSsKkCDuVq9R4T0DVMDG8plu0zzp5P70ifdNLQVs5IA2MhcPwocMrzkAnd4io
feJ9cSTgY/sGE29YqbUXMkEJGEoDVWisFWuT7+iVezJ0vuzeveKdeUysqKjYRG9IbaOKvYLL5/vR
ijVX+6cu1KWZw852AFMAh2M4191hRi2OGxBgcH+qtDvVgtl1mIxJ8RW39zQh4myV7TISTdK1Pl31
4fqvfMZg7wZBQPebs7MbB93fmVabsNCszIAk0yDYn21UsYCyLDDIb32y1PVopUSulIHnqbsd/UeM
17Q8GK8Xf1x1+yzvDq2ogX02HSLoUwaLaLD1RBrsxy1xfOwF46QWN+r/Xoqex98VHWl0aVYno611
7qf5xp2jRBrWHqeOZxFSRYCdWv4iJs7dF6GXAMOR1ZlTJWIQchgicBTUgd2NLh38mmmpoZUeeuXR
JKsD9G4d9okU2O3QMgZnOgB5mkRLwmSV3ZmE/k7QGOwbgaspiEdPgGZKamwhx+GXX2PPCB0BHU34
/oH1Knm7Y3gjvkOfqcP7ubVfD48ylp3QvkH8h+shId7JrdLRQ8ONATC6glyFVVOpJr+URkJHZbcQ
bQGyGo2XLY4N/2iIdx4wx1TGONSl1EiblbRM+FUwJwEbyqEyKY5+FWEDZb/Gs1AZvxv2npy7rMyO
9lPZj3gCBzd49Jw50IcfdjIDzOTlJIjecfpJP4VTgcnTSrDyz/MA6XBnKL7TerS2E1LmIP0v3qOa
MncQ97sKlUXu0YfFB5zQsxcBIIhAEXoRcMkazX3EATGNaPdFSomtF5sZIyPlxZj65SAwb2szZtDR
OUvilEr+liu0SDlbX0qBGjhRkQqGBs6bzeLYLfDfnt2cbce+QSqw/flX4r0zCwIFrld2MFu0tXmS
YB9TbHnWmkz9LYwVTku/nkIiMsdwG5nF5nD15NxaPP26wa3syI6+gZDgZeMWXBj1WYLnZd37DQjn
UOqBhc+J3sM9GYDs3dAhBPr1bbjXNSsSAB6u+CS3cQh7c99ev9lFb135QDmu/9oh7A/O6esMsput
3Wc62evIEVYrraaenVWtuUZEJSofOiCHo1E7GjqlTIA10r6DHn+SGFB4DHnXkhbH75QX4Wd25tlf
keseaYkt96+z9pwjMzmipzh1uj8Zkl8esqtFfMX/0Nzgrzgd2x78vYP37FubFzaoAYLytdPfUNWB
58DsxXTdssL+6wPHc6x1HbvkPLZfZ4KLOg0u8YIULV0/3Dl7pMTJNgaPbwQ/O1Ew0a1S+kMHnY8o
wcaeLIAjpTxhyBw4ITomPdNqle6y1PSaFjQCJJQuCvigZHUKRsIIhbL9ZTY03TWdG0j0wvlRXd24
OFNqkG7cc/vDYVFVs1UMtcf8jp13liPssoYRdizd4d0+APK84Nsbv2hhdRKfLsQELAbJFlCJEBvw
eNvJqGScGA4ZhASzrReoy3biLhi8JHaMR363q35IDfBiLKjC4zMisf2/WVzrR68YDd5pFRh79YrF
B/vSnUs+29U084Y40kSDBhtPOSdHJAinoiXuRYakaSgQXuvfxO50cYF++JP48w6u9wpSl9Q0/LX1
A3L8uyL0J0/Nd/wnPSengzvW7+YPDgRMRXAPVUzg9PIJw7+8xlNoIeAvmvtCMuOVX3eLDFWJealo
jW1y8Yi2Cu2DpUrh2bTWx6uvMYcTJrjGItEU+ntZPqqRrHtSmuYCy+T4/hDMbnxFsaoShzduA0MJ
vYEgZ5t6mV5ftbM6ZS3jlXNYuTwrmjvX1DfCsntpQnDZcgO9RULgRJWqfxtVs0+OTpkT7h8Vq+1Y
B/5kBybN6FU7Ht78o+a54KzDXmxJ+sT3IcWKXRWFjmCVFkZyG4K6qIhKn9INQT79sayUKAo966FH
uoRSGGeKkcXLLWApgZLbuERle1d0R5EcvsGEoll6VWeux5SDS5+8qt0DCcbG39ABBUJe16Rnz5s+
W6Fc2m6K9ltSRc2K5VmmomoCJrobd18lQrP07VxV2Nz8Q4TgaXSxnTlK8N4EAc0j4WhoaWwNW2ER
4wRlat0TAn4aIs6KFJMmVUTl3Xtg9FWVFyFXwJ54MLBu52dROp1HdxBRrurd07jOZu5t/BWgmFn1
FgD4PVdu2QwwAH24W9TEQRsde3tVm49A8heG2AWXUZHEhfDuetgsy1TuUQ5o4+H0qA1wJ0CpeaUV
whAeUTImLMqIovMK3quM76V9MWB6xOaXQFEjAjhJdK5LY3O0AfelhrKs6JCpBp64wFe0QlKh4zt/
jIfNtS4M29XVeGgJVmD32IKfcEjKCsAsxMdCClST71R87HdWEXZFflCRZwHq57EO9obyki/oMinS
MyHX5FdVu1827gLq6dTr0TQzGhJN6gcYXpMlGrAzxzNlUDSmaqBMdcCLuR7CKAedypEqJO3PHeh+
R8h7y84j+2yX2/mbuiUI5r/psSU+drdBv14XJWlX07B6/klD392kXI6RMWfg1y4unVYWuTmxz1gt
uWR8mPEJ8bcGDOSToDKWka+kBgtbv7OAgdtEW5H0pXvHK/05LfJb0oN5oJ/yvMs49HdH+IhOjsfQ
mQJk1OlC7KS5AqL2VEB8SofDdNeCIj+kzDY7DqOiMqvLA2RrNjWB+B8LUqN5yJUk4Xy1uPzV0s/K
eOY/Ng/KZwOE+vmdCkFpPV+5q6E6RM3gwZ+aQlpExCX9PUe9CP71sC/uvD3uIz+oNTI5W103lEG+
kfN94yQ0BbSCjfGRE0LhE2TvQUQpXP59+IvUh7f0gy2sAasf2m9HxmNZFKz8iF6r6nXFfAMnia6O
P538uVaXR+7EWvySrYX4/sp6dU2dmh8gl8mh/I7f0TOKntENFxW9GBdxrqGuWuUlxcGQAULXu2EQ
22gDZIpzRP7Xy3Iv5BWaWJBQw/AFH+ywHSukxUpy1UbHRdvv8OeXbgHC/T5HDFP0qrDR6GQkyOqJ
EuJpH9LRQpJWij6lDDM6wig5PdQyU4xhuVm3ch+sqjAlMikgsoh6mak2ASFGcBITL//6PMN9YN8x
T5YN2Hvqq3TrOvDIliELtkmRrWob8t/fZl/5LylgQvDViNsDWEnNZTabMSwbPw//6bHNsKAaJRR7
uXEE3fJUmfPxbb8Wve8aoGvGJcLbYGz/jP/E2K4s/rQN8pOzfewaaX0ZIgGgRhoUVxpZNBqg3xng
QTDsl9uItuNS0NbH+r/7wmWVtmRXWWCcwgep/vvaZnHI+7MX4njxPlveiqL/BCWPI2VOMYzN+Dek
DGnbBDpAz9b1RcHtGEhQU3TVNjwS/p4rjhSkREVM/1g0J79qUDg5fvtsmjyKdHV8pG3tSpSxBxfp
vgFxNJO2IxVp1Tlj367BsWkPAZo0HCPKhgqd9YgqmrIu37PeoKOv1phGw1+5NsztZP449euh7k2w
+lrbh7ssfTjbeBktEuxq2CbDeXh8jEWdI0K9DVWn7REhu/0GiP40Ta9QieaH212yCrTukRh67y0y
hmhVH6yR1dV9PnkM7d4zIKhhtXAZOmKcQYQjVmy1hICrZqu0AjBDOBzgr495YfPbhWf4GXq3i1m4
VFb/tvu5XMUaMv59Kl9fjNoAEMskQIeWgO2CuR0BPYggKgwtBPqGdhBKmVDSSwezRynn3FDLCOw3
sbpZN0sotau7r9Ry/Sl5Aqs3Frf0Y/27jVS6sTKkoGTdECPfDZSybodJr+rxqbkMoJsGX+ewgurh
ce10xUM4XI0pCFZWy8f2dSSibnq2Pc0jWAeLK3PbUojeO1JGXJI/fp1hpWIUkxT4noiBV7SVftLT
N2Ttxtr8DObDUtYKUhwnIPFaj0Wr4Dm/e6gQtQSJWLm/sJoupHYyHHsGmFoTf7yzPft251nECYJl
uKMi6PGin8REA1Y/PA/dcm2cmz+BzIwo3xUH3kWfRsQ2Mv6bWsjhcIqFzhFubiS66Th0ixxJTEF9
rRMeujl5S0rbKsPNRKjPpkRye9rUhkTIqI78FGVyMIhTFre44gUQ0OYccw2bQssPc6ItF48sBma1
XSGnveDxiCANLhPkUSyPcjtdmOPHOA0zLAf9Le4poIE8+PaTe6cQxs1H3RcSTE6pOTe46S1kJtwe
TYybxmwrpVafa7RtcMVVbu38v5S8aAb94UQ+R599u23S0wDVieWhYqdquEmv0zjV66rUlm34g8sV
yE5+2gnra75IKVWX17xL0CX8SdevVPIILPdUKuHyGUf1j1DjqcjWzSCnctjwMrUPBF2CsruIGX/+
oIX0CsCjeMIac0jLzdqBTR18tAC242womkYcbFKUiaVoB3tL83HyS6NlWRq2HWuI1T9mYuXGJ1cE
ZHad3J3hllrqQJDco8BJ6bZa4B7X1CUfy0LWt77mbPYTxRgxTEwPQohxYRHOPl5BnGsH9BIEwzpp
3UPlVHaOWJv6ou2zajNEEEDBlqS3AMP7xgASvNEYqZXCer3atRa8KtEPIGg1qerpNVDRnBplu04F
3hakaWOS1tn0Ziq5apld/TDIs5K6ZjcZ7IudA1oAgqedF1/HQZGokqDdXXxSAZr3n2J3bYsVsWLU
433whUAxduSf5SLTb7smpzxSRj7ypSLdLvVdP22okq0rif4baOc0sDXVTJ8a1l+TYcsDGFcvIYGo
33AmCCwoR22WfaIlau+PCy+Wb/IeCjX7G+rmfv82WCmRKSH0p8p9vDS212mj4pRHcisRZEV1n2g5
Uk8xCoWUV815uEITFbWWUDZh4TRJHUY7H0Yajc5puBwhmUkSzS6skWdY3Ef9gZnorCLm/1rNdQiN
ASXR0N9qUVA8iQB0v52jAnqMV+NgjZv3eSSyMalj3DFsrhgOJFJ3teJKub9wd+rjUP0RheSwVUX2
iQJBZBHLGDYU5S3fSnWHMpBLcWZZVltdpLK5RoUnMIr82HgRGchNKg/ZwJoupFMgQigNvRwfBpwW
GhvVJansFsen098GdCrVYrbrQToXNfsSq+sITKhRj0vqxzaRQKQ1Z/kztU94haqAcPvEPAdtBazg
iBqKaLPgDKC/RD/wenk9huV8xVslEqp28VBkuOprqsVNY6/Qd0j+N0ZSiKevyRF/OEHnmBPgqg8q
zhccMjff3zMf9LhLPSisouD5HowZ2LRyJQPEBxAW7ISdU2JP7WljcQvNSYwJbt+zCDmpEaR0PrNX
qumGGV5tWDd0aqJSH7qPHUQjDhN0779VRaBgB+a6VEmeVji3/uKqpBuxaQI21SMqU758HQlX6MxG
MUrtG+Lxxp2LpaO3miPakdXXVoklRuAc5yS6v001LXQttopPuR7k9F3FWmzRkmP+XsSXNecLGAbV
WVVe/W5CjqkoTecOdZPihMYMtJ6qMj4Yxt12k6ncMsWqSlHOKVH3mrp0LYUWSB1e1AKrLVINKrsQ
2zAkEGshZxBBLo3gfKdWO336Gnwd1COhl2FQdciSprS4TAKJQ9HXw3uWGpPMJIK0hw4z+KWAXE9g
ciiS//qb0goPdQ4jVnCqBaL2MR1dnM2x0kvVnhS+uEHtYLQ2aeDYRN7m6ksnkrCdeROMH7uZLh5Z
ARYLv+3rb5vTU2gCjBsv/KNn7PLhWccKfOfKo+SX5X32IGc4obEOrLB8HVPl44jHIN2e7fL20xOL
76t9R80czTmU9/ZKA1zxMgRPPra93alLwZBs42Lk6QUJov4jYpq+6eETgAKhipjvh5FlKGn/Dk+A
NTeJf0aXHCTxMJzRuFe9ZnPRQHnAvxZQGB49rJmPgLgGI01eJbr8rTA3cWx6sOtAOZ1h0r8/Ky+f
wdCYWh/F69mj1QXOq2RQ3OL+B3W1iVxAvxXaOvV4Uf+RnN3KOqr6SDY5d9nH2xNrObgsFLE0IUkP
JY5KOfsCRyeKYZBpt+h32xNpTSBMGOvAgydlqcy5uBa0DLl2HCfveL42LAddHagCdx1IykqYSN+t
7f0jROb/9W0uJ2lLolnTKOHk0EhcNNIUovB5nueLixylRLvjDNPpI9Fy3Rf/iq0JpINpPL31ro2T
aVO90WbSiUELc43pR4sYx7ytRKTp82aJ8+jrnYZ9H5YIUFFyN4kmZG9xA70iwV/oTZCTrbJYPjmg
LUTusdk4WxY6Fz5aaBevrAw4INtwalDCaH1em+LAB7zU2yIIlsmgKrT9iet5eVxyg4aJYYUWU21a
ZuYVM+CaaCcSwyx2wamHrUPDCDxvnSaz/eHweYPa4iLxobeDyYRtQGbY+bmKwTHBgAtMiM+lUdDL
ims1ZbYtdVx4ZFv0WQRFLv02zlRo6Q2fgM+d6JXWqSj/2RLNeWTqccnYDBoL2RF+erPsKxs7V54s
AGnlxhdC1tR+crOhbXIMtfiHNuuQpf06BIE/okGPxzFV2ZybAD3G52B8ca0/MdHwuCLJL59pqIJF
WNyBOyibRCN2LSAsgnO3ltzUFHPAB1EmFChuLn6m2U65AxxaJlf0teSj+giKdA0BDwGrpnOnfa/V
Q/6FIEvaipE8eHl9cMX+d0k7QBZbocxiuofwmZx2n94iXQ537X/HqQlpOgRmZfgmycJj68U3D2lo
LkvL1vudf72HDX2ksy/d/gpcEk+t0hCKt2f2ND/AqT2dFE0Y0qsGiDBKAOUUfXJasamPTGG2pAI8
TH/KTPctjGs0zS8AfrDYdoJax943OoBsIiK2b6Fn7TND2majNfrwF4Ny72HR7VJG7bCksKqgRsjF
QMtFBQPtK2LAWC2iaZPRD4oNlsh0AQSD0IKle5FxYIy4RaCd8RMXkFrFTYHqn/QnUbGcAo05Coe/
6QpB7x3TWUmJibZ5eKZCloYcCmcAiQL4TUQmny5qXDnJ9lYL/FJYc20VJD+a2DzlcH0zAizoLcRH
urNiHod2g4sjqbQfHB8PtTkPDUxZlsSfkVeS65htOgEemA3+e1eO1MBqxo4DEW4k4Zu4bbQiH/6B
Usj0k2aMYrXbRlzfCnLz7xVUDV7VMvRqKFIdkdQ6EVHHUP3zAsuVjUaRuOaSMWdTZDyATcJvetFx
ZIGAG8nrJbR0Mqb9gaC4vpEpD3QpRfsarebH0+ncAaXIp2DF3xNpY78y58U675414a7R2jHVRsKe
4oqgHuxY1e+iP0/cayrTPDBJK1NbqdU73u3uArCiU4tofhP0h5HLZmBQzZ+kBQs+WWdkOJ+WVdOj
xIJETEadqhOxDbDlutvG2VxNbcuLIveEj7QLbG+AFjiZ8tMCe6j1kM7uV3v6CRoD7xCneVd5DOQ8
OySQifycqtzxJzMELuck6OD1azVc/i4+GEKGa15xrbbfJpbU2naDXe7BviQJMgpho8XY80fLK6mA
On4vzSWxd1F3X7JIyww0xelE00or4lJ/bIqrSDaV7+LY/FB35F0eK6FfCyLRH55Ef7QEkCPBXuyZ
rs+9lQ05ifKSEyPcMZdPReikrjqOh47UaJomW20ZtqUGkBy4Ip82Qm4hyBzGy20jrLb4F8p8Jq0r
+9itJbxgeIqhlXK6KEJ7fVoiAaJ/WAWUCuhf5R15w7iK1Vcj1z7iVSQdMVD/wSLhEnEurhgnMBnR
bCtQVrD4VhoIZpc35SBz/huqk/Qcs/X+jpFdkSbLM43F9RefYk34ZxyedLp4RgM+rArM9UgYYo+A
vOmDYlkOyGL5HjJijvvDZzpPPtO6ZEmaOF0V+BX68XfvAHR/9aNZhfIAXLnA/nOqVbSfYj9MHkAK
OX0qhRWK+6u5hvJkU8iTjbnyk2y/k63vdPfxJpxOg9SNkGWd7EqvjXze5PcWnG9/LJ345G+Ve0uL
G9f/hZDGPjtK45AdQl7or6XWfYuVN+VR8tXjfy7R+TQfGreOoEoYocNB+W8UOueh6znKAY8B/XIV
XbIXGry65WCdvVEnDia0n6h+WF79gbnT5AiWhXTP2k+B8U1dMY5fPtJorMedgYOTDrc81fvLXpHj
1G/EbNXD//BmFDL7cLaQuN8YW6ypHmmPtlBDxzcbrIpZruuImzP2VA3Kjoq6ppo7o8xlKVPAHTIB
SJhIRI9FYNXE9eDA8ucUJxc29YpiPMXwLQ78wKmXdbGyfyc2YbUUIhvpmrxlym3PzSXOwnTYeNeM
orPkvAPnEQ6dNYJ2RrmN3gjEiBVF95nDza2aRzeO51UAmjjhSQJA3NxYAf1DTrhC5T4t7Jhbfkx2
eSmCWzCuW6cPITk6Fe9gcawLb5daHyJl1jzEqDdmhIiTiNDn06ownUMOwv+ebbcL2iCpH52Inulq
7CjQ5IeiNke3it5lyudSpo3laX7VG1SWYLfKw9T/zqWxmExdTQmTc1mCwoyFqLwSCGwHYSlwB9RB
87W/fT+ufDfO3xMfwuEucOr1DXFlplYLRFfuO5p8nsmrw10htJ1SjG3iZCPUhHz2G72GmYRJ3rPB
qIXxDjViC13L22+eYM5eMeAT0yXtyUIiMDgjhv7M8VaxNqE6WJThuZNMwe4D4TODnfB4nOAtoVxJ
7+2GtaZrBeMQGFofnsbzhQA1RhclWTAnJf5/UPKFOB25D8bmNrJtBaSLMCnvmunQLocEmVHM2Zo2
yfF2y8z+IdteKbMvEZ8PbhWGJQx3Wntt98odEmdzWMkPTcs3pPKWjk6vsw66RabL/3hkmw5QPSCS
89ifNOMAdKEz0yPBjx7FD2SL+ygvX2RvkJ1IIlMPrRHDcbMIkQ1V/qnHHuvtE/knV2D0hOTLKIkf
7FZoRNGNYpc5eJJLrhHvkKFqOEGZo/xE2bvlt5G+B4cuFzAnP1bZ1tQFzS3RldmAp542bjbuPwl6
HRnA34IeI81oIvBSFVZmAONxRvXSZAx6ky+rjfSSOd7YmALNn23zj3iTOMRNMESaRDcsLOXG2w6I
51YziBPkc+ju6ZkCiFDy2PIYEm1TJ59wCsyCpswC72ATchjzQf/Jin2/kc4SC1g0B17KZzfozX7G
pEbxmNgPh2goVjY12t/SqEIbykte90ifELsivXD7hkseVAuKM9Jgia6yAP4d5o10id24gCO0aCrS
w8HFwY6wnZDUCk37gaFoMPMb3OsQhB9mJRIxb++/o+l4pwAeiZNiAdeQvVo6ruH+ZwIwiITYm5H0
mXjMkg7tE20Xl0Onzg47KBXVTQd9fQPFKlrst50cOFOMjMXSWrHlzAIuujgxnmH36/YbKNARo4dr
lt9AxUAeRtsBoRG5pHiTOjGQIMbI5GF6xVocbUp1u6Rcd4Nyvk3DEKdjx7rErBHFd/cWIwnegZ+p
7IfY5VW9dnqpRn5EmrsfumvdmxULgZqY6MEJHOMEHLI8ThdaQwr6VDxIBC3dTyJ1gUEcJ5jnxfUL
T27cwiD8vhf6s1lbDmeoVUQbWv5UfHwWky6gbwXdeAaltcH3GHKEnGvirhdL9QYakUSKI9a1vVgB
z8eVm/mo86vpiv1VyVSvqo8goqFhyimBpj+QxNizIqcN/o/+KH4EYDx70erRlH3066RBMVrWWn1J
SL68G3NjxHUNfwCncuecplUGeyBWSsqU42xR5O0dfUVtcwETa0WMv5O3gE32Zy7XOtLtuSuoCoMs
+6dViohPzdZ+u8K3kbTYYpVk00neKIhKRbDlJKGE37e7p3tG7piMEycL7z/ZQI8OP9Rk+2vnEBuw
XevDYyZGwBLo3fG4VJ4/oA+YO+9e7Bm8I5YEPqzC+i1BA26VMyGIN5AFL4vi9sDTY12M1zKlwCai
dQgZReSnMoM8M/2aOJa9MccKV6gG9ESNLm2LrjRnrbyVWuPt66ZQKkXotz/0lYPTaZi7P/gYm6E+
tGAtUHMolcpzR3OSoCgae+PoliJL4oYG5slTnSamMRVPKxSGEtjABpoQrHhnXo+8oOcz/KKVXQEt
oRlsbTz6cdJEku+sqss8QSAXLt1HzPCGmKa4TwHpQPjzVyDLhRRxuaGXtejqmcjNZPl2dWF2sPHV
lJ80KNhD3r4NlZW7HI7JWMuqAOOeAPSoZc1Y0P9uEt5Cml24Hs/fOeAV4BwkRASMLY5LzZlL7xdQ
CFnUUzc+UHGGChJXPrscpCmoPgp9f9ZEyf0KvLvKjitndZPFbv/jS21BRs5Xztoj0aWasQONqW7r
y5vfYabG3cb+asy6UMfZmN21tSSP72jCeRcGcrq125lTtKI3jYQn2cYjY7FA4yrPsO7K7Kacg1sh
MlL/OhKk2N8SZCWeviWMwxjZRjAdK54ZfevKFjcZmcC3iX7dZM0KluZ6gEsvaRp8ZqmTIRkTkcvN
2SDm6zoK3/a3Pxn77yDf/QjfWwKV/2RsfYMoz+wSGW6u0T2iL/iyDZ5KHeUsF4XBpEKqBhmqrcU5
ElcLvySAwKce3HFV2A7CWH2qH0lxe7j6KGv2zRn1RJo94Z0TmCkYlK7FpmFXk9sK/pJqTzBe20mS
kUuM+WRmTQ4K0TFle52snzOz3Sk37SgRAthp/whuPqBhjfdm6MJ3zS8jqwz3ZF6BpgeGx4kZE+qk
2cRy/gftzGQSh38hmMIslfhH2FkHBifYaLOzghDjD9wCfJHVxIh1GeBoI1OfbMFTBiQK0+CIX+tC
oGrrjeCTOL14y/JIGOqmR5KIsG6K+WFRgE7UmDDfDHBuOExO/MyQrBV3q+rvSz7Dc5qEc62EUoR2
jMon5Zg9/0Lvk/QHmCDWInL5XzU6CxRzgrIc3bxSf4OwOtnB1XGZPkHhCe40gOIMlvOuIOlVnSdX
+1gmLGbPvLcCzDle6RwKwbSrpOv2DA4eriY9JVWgB9yjE6dwufBOVHma0nI7O9bvuwzCSXnnU9zZ
7SdtmcrLWWacBAAwj9KkGVl+3P6jrmU8lcXCcV0/jwTqDfaudPOufDXSWZbSVk8j09evqY2qawnM
e9Mr866BEXWfjjLJ/i9dDxyk1ntPtXlUYqKxhqf9uU1PtCsI++QTA9tEeVwhdjiwY3/U/INDdk+W
FyBix8AcNL4dhrVg46d2pOpjw06FMHH+mc4h8AbEDDXtxAuP14lBoHL3pNMAauKEJ53AVS5UQewZ
MNb1fmLcxIsAwtymxIvcZ53fSduDYCisZVbuxzqaCZM5PiSZogJjfClLN2mPXkl4Gyp4WaiAwCAo
5kXYW0uU010EQSosGNBcmrr76K85JiXKrU4AUR+D2t+39FM6I5oIJOYQyUjoXDfSpXUaSDixya2o
6Mn+M7vAdBuFg1KIRPsLwZhCGUReRE9wH2WCu9enf2roJU8fiNS+WmkM3Glb3tOaEANz/FGtqrT3
wzuxJZeRw6lg00dO6hiMLSalHiFIMJMrsfA6wnUHIFAkhNl4VJLPCMH5L6SERIum/TbRFs+Vqu0F
v2cr9o2jeL2iTVOUMi8hPQXBI5G9mdsWvbwZdacnr2VRdc0nVz4zAeuAg7B6XFLDbdZZpVscwneX
/PjVTtJxRLbKBtJ1UyOQ2T2gaBp7lPgbEmRUPkWjkSXBDLHv7vDVhekxSIIhXFjbdQDivgLgA56W
7e7BiLt5EkAbjkp0xrne7QdMP/5IoHA1jl/48Ghlcge9kVfCWkpbhloTxTV9kswWD4vb+wLMkS51
XQbtcS9bDPN87+AUvJM8Fnz4QCHWChXbazL7s/cTBuanRdcg5EGUX5tBRpV9E/S9ax7p69VNEoDE
gYR0njvX6KsRMivkTeP1OxL1mL/VR23eG1fZOBgEkbBkl86BkEXspvL/wEY+ZAlfMJtnGwXxxIwS
zLq1c8KENZeszLMxSD42HaQR37Bkac8zqATSbLWkyBvupB9oT1e0Ik/P4BH4m8/uO0FausAOyOgq
Esfd1xux1bZI2LtcmJ1+EULPBsoKHvNY9U029PadSuVzS5FmotsYGumCDBV5In1TCiO8T8xE7Tr7
mfy0LEiOg2iblDanEgCt8tnBdbKNHuVccGThcng/gZtP+9OTH8FYJKeCjfYCuc24e7lTOuNCJJJj
UxNrts4QcLAR525qqfQs8y8Qa8+H9okhE4DE///1yrYt5jnzZcgozC1zI2jw2Jixm9IJTeqkDtKP
R2fSSTRw9jVm86MjLezwchwx2r7N5ncxfdVYNeHHt4dZ1FFc5epO8PPVQwcCPr3I+epaWaXYSiwV
BXRWi4IzpwR/xjGJNqqGcE6c8JOX7mfbUVfuRQEpSW86m/DfMpqPA6MqrturnvmIcPirH+q32kdN
mkOR74dL2lfyVwMJxSlHiH5ojVY2h1NhDy3uagWdZKbW3liJKnjJlHm2ds98WoLnaAhKXmeK2HE4
sNz7cye+ThPgrTWMQCsqaAaDuOtvlLyDERAvDjCL+VLc4Buh8YSG4Eg1eV4QE/TrVkrmLjOSvjRN
pMkfqtn3KqpyqhfDgEKWMy/XaJbR8Hi/WRzc6vmZ+0Y4nftMliJclcr4TX3lKRH9Lw2/ACZA/qP6
S/tKQHAGspjVXi6G3raVeQk+i1pg9Oo5g8tfdfdVNyDr4By6EFO96DXnJ2BuqN74+sZqu/cn1FyC
1x/wt6DJZT3i/NVnZ0m7gSDUmQBFaJpEmC9bAZ2r66ShpcATK8ToPZlEYMBntzbxUCQV755oaKAX
PDrbFNXXHgJ05Vv6J/JnR5k2MVCFZjudDTt1uRucBQ2I9qqOoREBQ7xUTMA/MbuCXsNotD8D2YcJ
6Xy3DjW0upaWZ+FPFxS55tHnEaggcqw1oHSLpwSTNDNem/qhl31Qq9iO9KzQgBfD8Qv8qeoWrh3P
33PI1emByeCDb2NORoOMM0nCffTqYqeOMed1WdoJQ7pg6RtcVTeYt4/Rr/N4XSbOQ3ocRGPET7gp
buzEYZ/jglhjl4s255h3mMwNDEE+grqfWnkGhe9EwI/tRnTtTqiJyglulXGVEjGsOcVpO/beVV76
NyAJjWtazxj8MMBEkBfgMkYjHkux8uUtoBjfvNALIw5l6pldVhSR68+ZPbEDZE4doUlw2mJxPJhC
cRmxNdA10o+W+BKzMM7QeLBcQF1MZxpLGZmEaz+9vOvFDk1OJmq45BSE0jiDBiZlEdnmDpnrAlvH
/V7rlVPdgdutLBHfE2MBWBlbAanRMd4CLjZy90WKjdYdimg1XUKXD+w3cb8n6YXQQvwjCcNWbL/I
DqjH0XR1vUFy4OsXY3F40hqFE0ITjApHCxp3E0yvFPhWmuLt9B6IRs7FhGlx4gu9slMvSBcDlgX1
+sHw4qB0f3dFvW93tkJN6YESdZs+ICuFzr1mrLcgLEaWpuCDhDnilAFsKhYbXITtDpAOwBny9HNN
SeyArDczUwDmUIK5h/S4FAJxzu6kSw5cZS5KDcUDWXxEHDnuhlVWzzQohSnW4+6f70C6D0TdsnWf
RQd07uPpZNsgMZ/CNb2OnSLje331c05uUj2TNaLHQFr7g7okVa7UHJNct4WqSRbHeAcW6e5UiX8d
kIMT7TGa7AHSXR29PWawHfjCdsnY3ZUKu3rhMGQujwzGzXP4hTNmWua77s0SI+gdFjweOx8qJqFm
VtG0dyM2t3Jf8xqhi2pByYFFhuoxTbK7vZqu+NHX5s/5nyfC9Pcviu+yhXGj34T5MFVMn+UFBYKr
VoTRwcPWokdlJgMTlcmTeF+YAF0SFMIzixgmiLGKQKSqs6IAUIBgjQ5Wj2Jw5shaMEAev57woD3L
+r7tRQRfHrDFn7m025ldCr1O+6I/HhUf8+Hn3FcCxn/DAMSu6fCUP2u1m7JJ/gR7GInbs1YKUucu
318/gtmv7BlV/xHo/KQHxR9FOLdTIeviXDB8N+Oh7IHFS8ujMTXG7X4pINTvT7d2fOK81uKiSL26
NwO/IsSPPqN2/R1bjhBle5OQUifylm5YATOmdC/+cfJ+CvTIL/B5iQraP2n6MiFJQqJ6qd1S4ULo
1SPupcrgzrUsnI91o8Hl66xABLsOyao1aBUGAigk4hozSEC7TP4qkl+Di8S5F9xpbaSIeiOFDLBR
8Yq9E1lzzfESipjhJstjatwC+K5csvPZW9VqPdNZ2vYPJjJ6P3MhnjluiQwm5EPcoyw4NcHJorPm
pHP3ftb7FY/S4Exzn50UxB1WfbEN/N0JpNYO0BUumfzuvegP7a3HQ88I22HnBrZm2Tm20sUNyaEs
+PqXnATxhwvLg0wuVaKfCq6D4T5mkrHk8OfdzgdwfmMSsPMiPaYKPcr/Hqtq8hfb0SyxVYR7hWPz
KBqHxvidAIWulWQfFcb8iaH19I8CXWsxjCquDX8XQXQkEi+T4VLvN4fHfcQYPu8tpTHqlv/0qJjC
fwvOj9t2yaSmUU5qhmQrqwnglfYe0CcOYuQt9bbpnNezgntep5toKeIHTkFoSm2VYbAJT+Wom4M9
xBsdDUJRvXs2fKr31GF3HAwKkdTv2I41Dorio49IwOjAY2C5ksK34H1AYM5T3fd5eUcwfcNVcNe5
J/zv01+9hFXJATTZBOBIYDqpmgUHGzcx+saL0dIGNN5tsB2t9ay+U6910WF764IEN6XwXYEIljVp
QXu4rjfnu/kHGHbpkUGmI38y0ojIpikyI8Bvk0GV7JumpA2a1DoSfOBmOU5MqFconsDEOrgTDwMc
lOR/NR9IkIQLMYID5pl6/OImJRdCCvun7hVhwFZRWz/gPNYofqO+4YKRabbJrNc0xsIV0zooUDnf
dO1QA/8AKemRUWmmAnyrJ5UZ7Xuapkd+qQeIGRoVS4hD0n6+2PwenCHYokMU1yjGEgPigP99Gx06
KCt9HKTjHbIZq7QiTrMleyZjKg+aDFE43egDxL7w5DDp7BZrsVbcPgEub+hCShtS+z0nmOVmLya5
lmo2sk6JfGfyDClM0mw0dcyutxT9URm6XEeUg6J++kSFvPUuIMwFWKs0XoGQfOXoIO1ZCnh04efK
U/hpVespsT9ps+7whYRo3UidN6aYMfJnQ8MaaORntWCkGIHlTM90qN0o4EZrFn6nM4teewmNNmtZ
BrC6+lAvPy3JkH1VtCGuouLLfX1pQHfA4Yrqd6fhndQNjyB0DPBj3MLk7DOqZzwo3XfKxXfE2X9A
gK2dpj6vrGQ8EURaKaidIkrSNbTf8wfvgoQN8HCJaXHqFf7LrlKIt12r65C6VR5QMogRA/EHhXV3
ZUOaqTpl8/PkGJo9+xk+TTfA1R16prscmKxwpa7RfTzCJTyBDEtWPWyV7ZRSRfvkeklFoJP9I39o
2cWBYFhOq1NH5G8dC0COQWZ2pseEJ2r96UBb9HP4kkYnuvHwuroe+fcE0RW07ChrTch4yQnF/qAj
co4YOmgmKlO6e1Vlnu2geqDxgrGNcLJE7BLTeN/YkXB1Hvfr6puamGtivDSEjY7j883mXhzCxFJx
zzxNHP1BWzYWkSgX+alA2tNJa5c91IFEXetARIsqiaQ4UsaJdjNEBmXcyhybseUBsT8Qq43Uxtv1
p2Y15+7X+hTTeRhPfCWR8HaxU0n+DiRmkqCrdbTWVp6JKo0xEBRjHjsixyW5+Cy/y/vgPt5zaBO/
WtOr4jMBPc6hcdB+Tylbqpto2QM6Mkbiut9S297k5ojNCWOxocWWcrmWR4tlViT8LXmry9UjdcPA
eLS87gMGTSfmqYUA+lz6P39jbu+GWzqNaZP+amOVjXIYN5DoNsq1swh0B0MGP/uKmwjKMsJJAw1I
aIHHWW4kH1Ix9TSzwqi4lcJanLwXiR0PCFWMckQk//Z/qFSiDu35YQQyM9a8BjjHtTEmBXS7xrtu
EeaGl+ACfVmmZC1C7GZotlwm4De8P8KhUt9Ke6JF9Uc/J7Zt0paeTcv4dY49vuLtsPBHmB3RazRT
foOMgmlBXQX9xcvxpXq31xWnmPTDJpwgOj/wy1sn/ymNfd2O2aT10ae4v3T2gB9T4Wwe19Z7fc7Y
ip6j95Ox+5K3oJOHW8TBxxjGxf1VVD2UA/KnV35LzCVCfIbzP6XEMd5AR9osmjhRI1qdSolIOziM
fDwWUYeAnUUi7lGAPnw20A/0LKRpjXsimzZtJo2odeOrxdxqcS6kQMIvvcVjGoxPzAFkY6+OP7x7
fDY4jwU3tfdQy5sNPUcLnDpk4ACSkTUwXDM1kAsGH9u/jgoZSwlI09wqDCI0LTU6J70oDiE6pKNp
wbEkmKgUbwHsHjKH3UIS4lpGMWaH7sz5CdaHLIi0+KrJY4U7GvPNbNc+s61HdWXiRK0U1oobnAUm
KmVuBlMPNO5ahJV0luK1W2RN+A8i6G17tlD+KYKvye2I4a49S84UU8NSBOqkeW+Q0CxuzAyYNDgV
XlHAdwKKLlokFJ2Pfi5+s1aX5V8zA6ZFDISFffUYmflB1BMsabu8WuJ2sLAnRwyyotXYS4gCumai
YseNXT5CtMSWJCZOVEVn+p0QL0+ZSfxQTewXyX9IFvAfmGwnluFkh4Zr5lFasF9SxlcnPSI92DuD
YJApNSup0K4qfJPuqGspgHC5pbab4nIFqbpWkiY1TP9orxyQm+z12Bxd6GA9cx36cDuN9tGxscvH
RBiIFedxAWmNfGbkM367GvYirFTH8pP2rmP66LRpPhRdjfEJxtvikgoPXPhWEhPdwTy9CeewoJYp
APWjLOkJVuI1evZUh1cqfRM3h0zuTkHdYyuBW9dlL1y5NGZ/7DTagkTGmG3s5Zk3mphgSS7mz2u4
dciF5X0bQCfcCcSFWatizkzV+/BqgUrAsW1b/kkXdq4St/hgqL3SX95/ijqOiFmHU2n5cIBSvSGE
oVAQhZSVTSxV9GTfwNAzZMSBhmDewq80wb11R3JBP2PINyKI9y5maMICjV61x1utMO4ArbhEH+JE
xri5GmoqEV02Ghiz7KRnnITvT83svToWSSjQRYxnynWBxXnywmPzTitqGhqHDzwYpwA9Ai9CKWu5
xVwkTPkkMY+YP9+qJu5XXQYGLgW0l02FFnubjXHrmzKsh0CVz/3Espb7i/WRDmOFwYlYaPoNx4bQ
RhMNXAKQTiKuQCwt+T8vyHTeXD/e+uf8nTUeb8yr+wU3iH44JOZMmu1tW34VKLYfMofNBfIBMXLa
ruseeMWEjASbGjQn/dP9Z2yy+Qs28nSvSoF5VX05NqCh5wU9Xc/QvZuDuDrEy06728OvKWrTRjb1
yr0Xl4YvuLPG3FiCeLKg/xqfp4fkbhlDV8jKc4vyzpr62qJUbExkJnIqq+aokFz0zPetz7W+Hkhi
vzrYsNvyh0+xZ2LQCOGSuYsloY/WqjbMvW5piBJjJcVTpG1QKIylOpdl1eeojgxhs38OnykURFBw
jZIA2OLDoMb7ydTNEz49Fnwbhz3d5HyF+ecFjfpbmMXLIFYuvG1uGQjWDsYfXVUIDxJO2m4to+mZ
lLKwH9UokFUdfyxZtPFpgbHITkoW1iDXB9bJDM1hnaPFQhXY3s9iLmug1LhNkSe7MlBMnlP5uFUn
5LhpgGdEnBCQhB7xOVOU50PJfh8yr7P+nGYCOwhJEtQVYxLkpe4zuZltAqPoTZVUF1xdGm5IMlJG
/urIJhHeaqFrYSOu2lOOXyaYoxwt/ePlEbdx6BsgYb+1ECTN5PJQICCwZWdrOlBBhFPjIRcVOYnZ
BDnWzoW8Wwg/HsouOyTOHS0yDeFmQ7HgklsWzGCcVg4qHls+dhZzSnVHmlIzhH6spla1WASSn4pi
u+z1qKibG0xxB7adqJ6V67jXXmZQ3K0iWaULLXfk2XUr7ytJYU2QNICjf7kgUiJWUlyu3AgEfK/0
z4haeO7QVd6S5rNpiChHIqj3df6j7aY5O9/k6LVqAmZyMkY79oeplqFSu3jrN8+gb6sI4weQplNZ
+wKOPc5338/0Bysig+QFZqvucBj5BEMKqN/kYbbACi3GqBIbClHNnatvvaIn4Dt3CCfHJo32QSm6
z+9W75InU23vXWMsetgaSFELVFUTHw33jMd41GNHv+LLgRnqiptLlNm4ZZ4yXnXwy9EtP50bVCrh
DQ/MA5en4KU3Dm8QdY+tLiWaEZ4X21tDA7ZCg4Kg0tlTyrrAToC2iLIppjv71NbbMPgzwDbXyBQQ
Aj8QFz59J3W+x/R2fKQyhAa5soFWK7rF/xfyqSUD1kBT5CvsL2G1TgTmO3TcjbxYMhy4X4lc8iTy
owWRi0Rnx30grS4D0hjHkDAxwOVaQFgziQD5vLfMTnO2hl4lQi3w9DQ9wzZKu2354yaoezV0wJ2a
twuSPSEyI8MF1y+DYYjuGm/BivfQijTtsI/B56yxxhuQkiSEg1VkuvMQcmzRCsId1u/eMgaIWyWD
5TOGsfjBimOUHEE8aT8JbS6yo6AUld3mvJ/MHHc11cE4QepZGfohzwGv1p4vJM2102SuhHmEPmsM
ikXCkAjs6R2X9DhjyIgUm15XKDzGqg3EXZQyzc9yU1bJGsBwC6nze98DiRwDEUGFpZ0M/s1IhtuE
ZXyL+uTYIY6Dqf+DVHoJu6m2H5nnZTXY2+xFiAEm1A+0M8UoPhXtUmZJUBLq16J6eHdz5g7zgRxe
vawRVTz6V1nwhiEYEPpYFDXVE5l6PUzE7hYf4kIsL58umCZR+MLfLpZFHhvmhAdWagL0ULqvSMQ0
hLIQgknIYxHJ+s1pWFCadCd5ddkTfXBFdAxp/eMHybP3mSjDIOC+xfDqLZOMxAZJEs6a6UkcIYCh
TrRnbDc7XWdrFy8YNR/4GjkWwdHJUsqumukAmbOZFcrpg99Rw7+FDS2gmIw4tesDNaYvTjRdXmoR
AC2nwHmgjR1pFu1JFJmxOkPLzSVOMGLjvlyx36tvSm1ruyRdNhTNkmKZjHYEFlIKoWRwoAcvFW8S
aCR2xZFB86V2pzpPe5E6gX3VkDAK1pO8+41tIHJxj4FbiyHE5QD4e1Wo8XSv0Qv4sF1WsvmQHufZ
O0yqlafr/9+/vVW7mE7gLjRFAgwHxkXxV8Z+PG4Y+h3pCZ15kSjVbibDAvINoEYokUhYBWabe1ku
84/2CdLiKoJcouGqJEWsT0d49qc2ZH5c8+/NmzUW5rb3I7sFhslqKKoU62cWXI0YtEJRjJ4QF0al
/rZlW30jyfw7U0RFG4cVEVylkbcnr0AgCWj5Jb3H1WZE23CTTUYQjOm0VN+cpW2wW1tgh+PJzzPk
6uNS+Sxco8VbqRg7GKl2oteEQDvy5C+mY6o+laUYYe5Xj6e7UldEqirjsoJWV971L4sT/irfuOlM
mMuWKrZxYaVTN/1SA092e4ri6GXNpmiKoG9FyKsX/tPvhdav4G04X/TRwJ1ssYb41qneOx7zZVNL
nTkQYcUlVyMD6D+6TssOXaZ5/DXBbMRDkf9LC1vbB9tr0IsE9J2AYsE+3aSnE10xNMnfGcD8iKqB
dwnj1pCq6upVmHETPgqfsIRrmwdO8fLYcIrJTULZlsMXAiQSfb4YxLrZp/bCLU9sa0crmu/M2iGd
UrWx7Cp8qabTIHv585BscGlEWYndWNJtF2f3ZBIL5nd8Ce2iM3Trq1wPd2trmQSjryMTGGJcOfmY
y231wbwq7wDNMuDW/xNWnI6NoKAGjALCF7hp/WFIjP9yJKZg9aQszP2xkAhYZPs+237a8rowwLNV
I4eK2YNaeuCCgNyhOGz1MkDDjEOFOlnh4XrHTTyrc4jZM6XSgxQLDCBsn2Bnh9B9bexNfVtgdqeR
eO93YTRimDSovW8VRIFtVvulr4RJ7sico1LkGoQg+7VbARo81On+x8mOLyMfrRs9XyPDjcqsqYWo
b5jNdivE7UPgLgo+hkLIsz+ZRMF1h/OkHZs6gg4FWJpRsxsNcTMH4mToGLb3T2OHzSZTxTFQ7UbX
Jz1ZNc/oNWE+sUihfA7ZnQlTepoRbUie1e3wGwGb2YDekesNTfMWgwXW+ZBILvwlXM5XJ4mt9omY
2vKteryv7uiKCpeEvjVcC05Vg9nk5/mn4EyNnq/mLzBkQAKCo1TNMlBgEHIPyXs81orl+1NBxxiG
temAywXdfEH7EDU7k6qz0eFiTVX0qpGUMR3txBPQY42qj9rLOPVV6f7GzpkUIE2Y9KOn0rYuRZKf
f0igY+MD5HkFtPxqdG7IKk1xfRxpGk7J/5V2BH1JlYb8aRWLyVhYg1elUFym2ixKYUNBfUBKPrWI
Bnop9D8qdd4EEg9YWMcjZUUIFPPa4GdS2s9rKjHSnHJbiwEtlZjGR3yuUYkvPTNikl5l9kOajXw4
qcrknG3oA3GkK5crTg4m/Z7vHF9T8ZBAN+CR08ce1MiESNjhAOr/X7yYVBIurak4chBttlycwXW0
f5IxJjaSGowwiRkGit7yyn+kir7I+rm789/4LV8DSglsN5Spz3ll25pRFWb5zNDXijn3bI5dCyWF
2lkV+0iu9EcfvfVWQXf7qOxFVjNGIngTo45rwoamQyU1K4QgpnDTla6ll5VnusM3BNBpJRfPNquC
+/Wwvs+1xC1H44UpISK5+5AiPKzpoUuavq3+cuXWheiE6wBvHgzIwe0R20S86wAd4xZVxSNsXF8S
G1jdbYYJOV19Cf70iG4puSh5oxt/YnQ5pawsPYct8Ds7lYWdIjBpDQCrnOsUE2oVWGETXQUAC1Dj
3obUvkOCbuiQkj1jwgtsVIuM87ujhsDQ/AOL7v95HRTvOgJ8UyCm8zTtpcoW4ABoTK/kcxP9+Rgh
mVVuRH0U1CF+W3pYEeRN0akTsNH1mdvtNwI8YvQlM2jkzjfxM/fvb+n3MxVG0quP2WELHDoL22cO
MiFBhDrNQm3cU7B2YdDCNe8KfDNbLo5ybr72F5hrvOkQU+HgFibIK01AJEtZj+eNMquuGQulBR2h
X5itR3vn8NzI62uZqb26j+ERs3cNSUZqZ+JZaRyuS/3vwYNu5S22XF23P1+L+iv+Kihn7gT494lK
7VmMuABbR+4Prdww1gxietVIEKnFC+PP3tVlfY0KW0oZ0NC2pPlwcQumXSUIATBcwBD/gxIcDl12
Xw5rF9N0MBLkP6FxJRy/sgEY5NkX8tlEFLRTEtlKf7COpKBiK6mMLJXtq5EWdU0MNS1C5Hm5xAzE
8Pk9PMc3pz5iC02VPAuvCuVmtOGqilQDz1q2bnriLI6HWj6x8W1tb0OorGFErGqPOUAiden2C++W
IJCnicvgHjF8iuNrs3bLvJHkckVabQkdOmZMhGze8gWOqzasogYTLNcF0JY/Sj5lDPZUcVkjFiVm
SNjqHk6FMjvqw8636gQ9xOb2P//lTWzPwrGmK7qAuLXi2UkzZ3ynkPEL/AIMFZkMHmSdqrKglCgG
zeYm1UKMZiTNbowGKSXp2iKpp+QCs0c9ZEtyZ3KwMZU+Z8O5zQ3+akxL3QqA6H46DAFdK/whVVwe
cgykGeuXfO1rx8vt4/R6es1jO4RBGyvNeDP5zr8gdRWadHXx1y/BEDm3LuYiWshqs9y6uy7ZAl4p
YE50vR376Nj0HWaXC4DEfpunb7+DJYqGQeD6R5foSalzlieqaadslH4WT9zxZkd/BAMyaQcoSVkl
hwCUtdsAqOiCsqijiDNrGY7TNNzf6rDyn+jSqT6RPEzI6B1eALJxpjY6wofzQR9yKtgpQFfxHcV7
FpREoUwBhpT9hWMtce7chfZ0s2JS2qxXyxc7curpdFp/KpMRjH8NsF60Ymdo+YP/wx89bMYoSVua
ytX1/qcyiT6AIoIgEakHDxlDe4VcxEw5ZKsgb0t8//G+53KjnZwCBckhkJXxGckrvkqBr6MdH1/B
dRkW2hNCDNwkzEe/1EDWSwnMHEpEYRbHEib1DCpp7k7BVzg6bj0Chr3HFHVk8Z09/s28i1GWRMM0
BVwAh+4ASFQpGCV3G9ICt0amcCc/mUNdCny1TLCUmrX6j0LsSwvZQvUGxwOY6jEe8Dnu1xUG7Dpd
qnx+tXrJJV8i5/lBbxX8sS9ZbhpGtoD+tdPlIeg28SvfigKJ1IPDrTEj3Q2cWFcX9a8gpYRbWCFP
h4PT3T71P3dNBuYI98imOnhDQpw1+OkZWD16SHf+xwEbanSoZxKhIH94AP3w2Npx3iy2/Yj5/G8P
cfZsEZ5WPnsuJwvxIpReM+0yVurxowEq1VdhIzHcvozIQmj1hYDqOPV4L4DwhT7UN3zyEwggMovh
UpPQCryI/xNZZx9tYhYfzPaDHUBfNqFILwkxOG7Wucl2K5CxVykaC7dQYRym2TN4AyKlw6CBeG92
1cVLcsxf5LFSdDqV6zBO80hl5JmbTpDWJ3a2ubUg+n5ggLjezocYXONOxY/Pd3Q45stxlKOs53fs
gUQKjdlqpLHArlmf8F7H/yYY2nqdCFFp4jY3O2ISI/nZmriWMmiVYR6Gbkr7ztsTQL+LS423oaTb
+GSP0xDrpjeDnlsjBMdJPJ8EXW4uD9uVSyVEjcSun88MlZvkPhVZmTpaf20Z0JrqseSBF1ZjepEK
Okg9bISGol2W4RSOB4UcayVzBlR6Lb8DZEX5miowxdivRR+hhKkuHmK76T+LyEA3/+tHxfS3dh3W
YnzUF2mA5etUcffyK9qi3xi7P3PzuQbNBcw9ZSQeqvi3ockN2dTswZeuUhHTlGu5ybewnN+TAriI
krt38LNwvzANHjJlSQblZnlnXkhp92YcCXgDnLxaZf4csrTwuwnUBREr0vZ3iZCdM0nXN0Qlx8wN
1HlNMZCCqgUkIeBdMfP4Lw7CjnoOL1hXqQwLbOq0bK2a8BnVfRrFdjbr1JDkKB9CKXrCX7TSEEPG
dk56bhvBK4vovpLg3LtmPVarynNpbsjnuToE3HmwXmkWc/FFRPCF8AGaAKJqQVlZ7XUV/criCO30
quB3bThlaOVCye0bhxxOR4Zm1RD9cDWHJUIek7ZixPYWS1nLAb1Euc60Ckrht9A7oF2V1VyudPGp
NbI27PIpvZ9Ilc+QbC6GZ3B07o4SeiAIrZJSjRhg/iLmBS7W0gffLnwQ4eGRVK1veoZQJD9TlU0/
o5ULJBuQYHFGG+fAXPr1cpbVuuywp1K+1oheD/nLyQX4y9NjdRr1vX8sTv0gIl17ox3eur6tqMXM
h/bUvZ8lOu1eIVL8k1vKyJEpqU0L3kCvBM/Yh/vXyBwdU8I8eeOWojq2KlkAg5QA+baDXGgdu7Mw
K+EOjwKaUBUn+avU9e9bXRd7fgsd70a/JsLc8ADvF0E15oY3ln2p6vZstjq0BSFLetUg3T5fqQKM
8ERuYUsElLnq9m02WHUXVe9GoocZB1GuJetjPgeEHaqXbAewkEIDTASSBXkMwZN3FCopjSFpaaae
as2DMmjqQugwqQNseg4jVf2tD5Sk+cK6jdYiO9YHq+azaJdhLtKU5Q8Tfrf1lAjDY5KP7Nc+eREI
GAuG0UC8t6xLbctlZQT/6HAm+sLVqmIpA2+RUTxQJbpBhpO60QW9BZno6mpFXe4V6GV7Xl8NoQip
ZKBOOk6Rw3LIL4g/eBNixhyBCyAl7tfOApW8pFnNGTzLpksaANbV2og8GpkAafO7CGBpS86ZwITk
awJEdOdCYEYpC0phUj4hSExd3f24aqBGtfCXUIkM9zVaVazfQqfL0keaqaMyBE+ms+H6OHAy+Lfu
oi7td5LzUYXbN9tQg5eRYb0PPFupZA26E/P+K5YsAaw9nCrA7YeJVVtko8e+BcWTbhbecyJTJS19
P9le/YkOZUUMXqdSk6FTzNsVafKZrki4RvVAVDqb77H1Sc+pSByblDeg+hZjKDU7YGFkYgL1o6D2
6ecqVovKusq8JqCg0+8Hcxy9V0bLkfTa/iVcP9bqLc78FpPvHfvxjbMe+w7Pxo1X06/UeNT7T8kt
i5LEltBD0b/cKomaaNZr/IosdR0G9WIwooZ59krVqsD8sNAhsJaJH8oZDYT9Q/co7xrNWvrWMUOM
LBQZk65St1YeKvzxa0b+CKbvNoNOvJxYjezIId3XZYO1qgnBkEQWymkqwNfRjjVJ7Pqi32kFOKze
O4vxxFVEob1trqEFc39v+kMu8L7+3E0O1P03OvQLuCpKjPkUKCLrGAxjn6UJ1QSBUHxxUXZ5HZgf
8IGShwhN5cjXOgAaYiAuEHePSf5cIdUOoNuRTA8YXBlWy76aSSQAYGnvuZSfea9GlbOVzFRexvWV
n8roup5nCPDLixjSyfUti5umll84j1dscRMy1/7tuVQx/Nvl8ZuagWbGccQDxbC+jp7kPczSJS+T
tVtyYb5dV57+NAiz7v83bczjz0d1g5/BVjltZoWzq/IdF8VHcMbOjaDJ3eEyhzAJpZ/DFdN+snS2
Gs7M9xjRFNLohTT6spjdIB5y/0+swltb/WZUnvQnWrAp3iNTK+66k5Znq18d23CBRsz0oO7GYMfy
g7gf2ua4dpIEdk2w4LW/GVIV5TA61COHGiRw7tm83bT3DP67SmL75g+2nC5LvxH/tMu5W6id5djn
FONEVr2TdA0TfZdI+TkXCIhYVHIry4N2f4m8k6OGNcF6dZZuAODDTe5fvNLY8PGkPfYP7fu3aVW6
J00KkwxajYLTwsnrmvUlqeIUO2zQif/8BUXVHuaxV0RK2WkUfTZhC0BvqVmN7Bu5TMytytdiOn/4
e7Pf/m/y76FFZvmKGc6qYt3IR2/Cgh+z9eOpKTdLNgPAUtlwKRr3d9xLMKf8rhidTAihYZcCefil
rlFW4wPww+1ghmFQ4XrahWxxQKZLAjsYruDtO2ayAehTRi0VJNPeGaE6HMqTfD+/K9R21FllhU9U
zSQeMVm4F0mUXpKB6Bu14gd1fAlMXedrBAPfQf0XTTRyP2dPPlm3EIqfWtuRCrKeoKfgWHRcUz+c
WA2X9P9MkG15BN8//JhDLVxH16qLUYawblltgJh19h/tqPRrlLWScAavwWHbbxDf58+rw7eQqbe+
gR2X16yQv1DD6YG/euOcpP+eYsQixOloxn+HHyvpU+OCPzKWcEsHihqYCwV4zsiHTktIfhT4V2Mb
wLFZHMa3HsXnAxGON5+YQCbtA7JKOXhi5nBPX8LpoPy/eufhTx9soTIg/wzkrVAtwBUo8pKQQpc/
/S8Xj6uT7NfhTpb8Imp3JGkqbK8nR5XZGrMPyJYtE0YMGNCMIxRqxIMqaDE7kaBwkYreGBveUP8w
6/2/mKcCC40mlSmkDJAMzoO57BRl6iY231/P1cGD7l2YoAGV2pSxWwuuAU3r/1Z/nCtZAxXVoVrc
od9StD1yPaMMy28h8sovoFnBn8eAZNt5/q2heVULMMFvXl//G1lj/EubG6JViiBepM+jKTs9+9tA
OJ7V70BbPApNwvaygQ1Hm4K8sYq4psZxJ+2OrvznJOu7QYXKsfQs4VXRx2MNwgA3Zx0BiL+62SFm
ZPHMpFQ1fepkaKyt46TBR+CncDWk80S2mfaHVtSvzbTff08XzVPMmvdHNn+k2xIj6bzPDvLh+Q4m
2FGMI7Zaflem5bdK8Ch+g/9MzwZNiWFhnCrKMrh3/rnZEgu7ry3xYh3cngGseUx9FLfqurW+Xn4w
aBUJbcB1h7DjxgJW5LNcq2Z5YM2OBCSlBKBGbNSvTs0UhEJIzhicHPSJLfg36y26PWw4bW8rcTGe
I8SZ8ennbpSFjf2LuqJZrKBO+MSGJ/iskm9Wx7THo0JMhBKClQUF7gKWt3oRvwRaMbNsRoNzuq14
ax5A19hGhDwyKoo2HgduySmweyRCkI6BS+ugjyLeXZLy7xzbgalPVkKKSg2uYj5bOTD+m4ZTf3Ld
zpS89spz3eZONahnLlN5YXOMAupYArJQlJeKEgfS6p9XR2G5tZM1nuk9GYa7q9ZvaPkalOXGILPX
TK6HSbHILSDVaH2lga5ART06HDuU2XgvR/m6zofQwmw3FydM8xt8tXBApClFMCno6e1ggJLCUS0d
UqcIRSyey1Zyj8Go3Pur7Ey3eGTJyKrzffOfH40tHEow0Cg5rMDGp5mutf8fVKCnTwDOSV0t/WCh
9KTYLJjLIkEBLDi3kz0k3qIP+jVuQwTPaTfut8MjXv1mHjrpLE0GFE1hJtd+4NRK3eryKzYkd39+
AZ1OdcJ7ZOtxABQ24G+LyLtWpnEAh+jJZ1vX/UGXoQxZKizMaqlMbK3N//MWCnumYSLe61dpmvEc
QlAYo+n1N//cm0KK4IlfFTkeoaSu3g+NXwUgx8zmWdY69Y2H9UhwmrR9kDhNFnBa/vvJvdbTHgVF
JdZEBZaRG5ePMrmOzVO8XSZHKw8fFhp2uPTvbLUVubhVzquT12daxw0qKeTc/eVf2yhKYQr+9ZmS
YmU6c8kxkKt9iK/P+KNI4msMKkEmEemWw7Mn+/Hf5bACszyBdNRa0BWhQQSf2WxQsUsfkAyrPDxz
ulyN9mvhrAv2qBHctmcUokvlyD0rIeDeDSE+yrAGU3nUkL8CAVabnZrwIE13bGmgP2RnmprPbBIX
9RFop9E4RjZQ/XfNwGeD1LJQOWKMSz5ODksa0HlskFb3ddO+hi1C150LLOMP8/w9n2DTm5D5UFW0
4w+pmpnGQjKk8uV1bTJAamlBKH/gTA7KUCo/B8qNGUzVy99FGA/5PU1iJ0gNobiX7wc9/qkLX38G
yIr6qtmHL2utazhKC4v60gcZHsGG+bzGHZmOW6fxL5EAS1T9HOiBtrss7ox1DMSyf+g1ULSGDfpi
v53d59vmxyy2f46yq9dPGmCsijfdGPyn1zwFm3HbNdzyi6Q5ztxV8EQHyHDeOc3jUVRZz/hm2/Py
/9hBB0DxfjeWD13z9gA8655xVvcS9trOKWFj9gIn+u9ZYQa1SQvnpmUv2hSTJ72MtfJdmzz+vpu5
E666scy2fTM5Px5iqzSQY4kAOHQ1I8L0lgOYVJFikeKiu21rn7wQ1J2gh+Ec6M8pR5/Uxm6pnM4H
A4Og+QrlwuONROt3bduQ/5ou1KkwzK1egdba1l28oVArfQ8Gv5yaFezMBrZ3le8hz9IgPRV/tK7u
t7bRmqKaP6ob4PdoiTI09M9hGEf+SQ95G58JNzqHftvJW0t7Z1b84WFkFNa12j9lcblyhzlZkT5p
IA4+gapnl2gCoBGiLCbyLvSelb3wnNzUenvczOeJ8FRFvH8FWZ4l5z8eycggaLXg/ypatfG/l1yO
i8KXQHpPHpu+2uLEMazJ5NUZGObUklV+jY2E3taVDn+C593paIbRPWJt+JpPm9L0/slzqCW9TL1w
T8pKw/HC6h2gfHLR08V1KqjPrE/ZtBOXsBPdZU5fC4/sWWxJLnjbfccALcwF9G7qeGOWxfx1I1tL
43cryVlbKSawizM6FFKYRsBkz1UadN6vWlQIjSdv8zEq/tASbnSSL7DD0fz4j6bi0LbFAahKDv2E
jJCWTnVAYOZmTVUG+jfIqNOg4/jzwQDTvQgDfKlq9nrqeehHdGqRaZjl4NQY8yoXNlzxE+MHG/gB
KtfkTIQFoZUpkQA9l5ydMlitzslSdM17I5dU7f4JAR+IFlupOUz2wFZaDPQQJjqbDLxeKTAD7UGD
REiAuoehhDPpFgZBBMa4hjUhDRN6dMt2Svt1MGSGDzgz/l16hAgkEDzMnlRlkYYm45vYH94/zRF8
iw4d8Y9bHyC+67q5VkBlO5RMGh6kJonCboTDglkfkve5LcO6UXwX9Z9li7MN8x+ReAD/FhJb7pDQ
mUtKITrxyc6a6EtBgKqy3UYfqlCOODhicGwY8+pgWedCUqhYV6S9S2HyVkSZ/mfZKUBU/AsIAQE/
W6jiciIXBxabuFAUYgl6G24R3RCulUBeVIunD2KMSxO4QKsbMJbNAiWzBfm0ovl4N2dj/NmQw/xW
TUIf+WMQbaR9XCnqmOrR8VmqFO9hlzE4w2Y2eR/G+Q28dd2CRYV5XbdgCn2MJwIXMfL6dt/2lqAY
XiuPZcveWbhq7ppvYNMa4Mf/rH9kTWAspXsiV0rq+PnaBeTkCIWsLKv990MNaR7qyW79gobBSbU0
JXAuPhfzIEqmJWLMLQE6ivYi0CNxYwmi05POt0gyiMzbIXmqn1CMkcbbqy7MazkFWTT4y/GbFDkU
yuzmSIcgLEP7jGMBhiEJR1GSzBOqXvwq1fVy+R0zIHghLrM1gHNhbpQGeP4aIdleDIDFZlq4Q8/X
oSu5bGWCR/CQKqsAqjOQrJmBYq6Ro4eBBp2Bh8wcHSbSgi93rVkCyCkuvgVt1iY3nbfMrNWyRmgj
/d+y/tEJelP6yMBsCKgLa3c46uPQ00V5JGNdTtMZP72yllzhD5be7qasRPvv/eaYaYONt8dUG8Jd
M/soMAsZJPSgP93b9Gvcp8EOCrZTiyANdIQMt/ozsNXlT6msi4pVh/RrqSJ9mny1LShqurGrXNTk
Ey2SEOI/oh0HqdatF6/sWWwWOwqm/tJzzyA4Ax9eN9Rr7DReQmpPWWLa9PU/9REguZ6gV2rzo55W
NhMMzypS3KLkbumq4WfTnOzRjYqTehdw9PD+yM2EbqFpeEo7+2WYhFzEa4N+wQnjJ98ot6entbrh
ETJPt4Ug1vJssSO+YyLxQoKafJZiSrI8c5T0JXqyHraiirhrT54hIHUR4Wrn+JPolNugRgiaRxg/
Ak9KVCn8iJ3mZWakuyXMe0nJDIZXvMbxQHQr+npiZ1bBsjafchJi89j4Yo4NOftWdl0tKzfisbc/
P+8qgmKkvPpptRoip5ZGPWspTK2Yct3sbUNym8xpf/ncXG2WruHp50MTSSaAaaSsfm1eMMi0x/7O
klLe0hhm5xEXusDeIBnYhsrmJpzxDh3Cgth/s2bhqd+VC5iUaojGZ+CPMivA+62kAdCRjdDDimRT
JJzfqBX1bDQePjIYReK6FVH97CuhDM48ivE4PkwZHQ51sgEJ+o8vlmWQhpstgsnjIfgTA5ReGogO
l/joSI+5mrrwEjp3Vcf5m6EbgLIy3twa831DRjmFfNH6ihz8ZdSjXpio5AKNJP0fyNN630b6hwQx
fN39JcBpCcecgabQsHGkyDLJLWx9BZrDvkrLlQu6GOTKOqvTYcshBFT3BfbvBS+Z7m62MT5JX0eo
/8taihYd5j/089GyR/r+fzCcNmAEF64bMtp5XnSHH86Ha0hczFSEOqXCNSMy7o4kmpaw5ZEZQndE
YLiz4+XedRMIA/bnppcvH7N5IfBNowddxAkhZWp6xP783WEc5uImhDvhfee/9xfy/U3i8yfNxSzo
QjMZdnuWB/MmQGUDKEtJcf7q0PgAIoWD4XUFfqFIX7xx3fGgKSgnyq5JJjOL3jHXa1/REZyYUau3
8DTRVMA4YKBE8U19jf/mvis0fxWpqWjpiOR3ALYHNoYfBBoyf0TvKX1CqntUyyQrCmF3tguZUl5k
5fNlrBz+OxmUIjfyfI7Vyztf09ehWEB4LtYE5c7118vtMnCfZgNILVHg7xaK7+3rNNlGUpS+uCZv
bLmCsEF0dGnf7kMFfGgUYJVddHVWlme96/SCTE3dHNqpbUDee812RNmbM54LaSKVGYGTIlUrV6nx
ernxV6l01JAV6f3x/ITg9pvhksqBU1J3SK6/dEVHtoUWhAxprnOMw/XNmIF10ArLNcpF6qasG9/X
6e8NAZGZ5tPSFKiygGoNJxAKs/tR9414YignvQgoWtnijtMeqUtE4pnuowLn6/sGiSG8EMCrwbRO
otMgMR3rGi4mnd3WnQnJrR+N+A4elWjGsxFy0MbFoZ01sZ7n4Mlo+whVD7nMA0CUBX7AaJcT9SH7
lgnw1dgK4Qa/FeSH3QOo43cdrFdkp4Atj/wJFRtps2YHsbsfhC7okj2mose4279PXAv/xLRtp8Oi
RTJXKqbcWCQ4XvBSxMugH0SGMCSn1WiXOmQ7XXJxTNRJaZMQ/GzKujo+Ln3VyBG16WeURuZn1CCs
hUVWbbWvRpHGe8WHgrH2XCAUFc/Msix2XBdJUdcXei716TlavMmyVjotJNqlgwoV1ryZUlL4LIFK
ZwTPoLQ5Qc1LHAY9GQIGoiFcHOVUCtnROuUmgJg6+QYo3wgT78j+IAkwL9tzHh1u3e94o9vQUYRA
otWVE0lOUZv5VNxnBfi/RQPC6GfkX8Ced3f7iixRcskTNtRU5Q5A8RMbs8v4NeKmhNRVlbkG+T4N
jpp/YzWqkM0GmFJAxCxQTIM6ZcC5J9AjvnL6kDVB8xL2gMeyfQSmrQpREXojX1Ul7xeicinywqgA
CgA8Fglgy0h3YbpDn81zTBY+teV345c+nmxc2KKqHHwCnxd7Pvla5pQTJyIQ1TxYG7SN10d2TRDp
YYHGWRwP2IbK1XsJv6aqlcQm5H7/H/o9VW0Lj/dh5WDAZAR40bZZylW1Zmw0L6WOqYPeDUgL1bPk
c2wzGohzIieGUemaF9GbdqGcIneuL3a/gT3zu5/kThKw6/lHhmneuBRJzSGsUPwineAY6vTABRbl
MD5RJ3nrQfGzVH4oculvBrzetQRlFoEwerwRqfSaBg21Ir48f4FrcRDKxMWqIo+h6AIBurbijeA+
XzktyW8yFPPW1E1Nou0Aapx7JIPynI682gGR78I1chQDS9hN2xKfuJxjtOFRweTazSVPXpDE+NRZ
5SsQ4UpxYPNXVI0G1JOKG2DTYtMCo/iA15VkA3aiXRs0jnoIotqWII7JfzUV3xVTvJHhP7fF1LK0
KGlh80ci6WXERKDpal2DhGM30lYiR1c0eRAfylBe/fLfQw2JSU14qf0h/joPU97YFUfQzf6UFn1/
uL2c+VkQ0+5VxHZ53Mpbkrh7BbpGkBs/MCzpR+RZl4TNLfSstBGlBbrEvJETAFbzfkVRIC1wJ3gI
kCNP0JCxpTTRjScN3WRzCAKyZLphJceC+vFATN7xZwavafkMUG4yvwKWPpHW99p+sov23Dygfm7U
VSkqwkqptjnTCyPHBV0PdTe1mBh8/KdV0K5CysEReSNhVmfsLPUlBjmwpdy2tCv9aKmZIK3IV01y
qQ4kHXSiU3hNTF2ak3NV3KVBCzfV+RxHneyOrfIicssxbe0pdXLMrU7PTiAJ2pyIzoJSZzmUgC3F
ebLmUjwbkGN3uUy0gwoeBWwI0tKNe+KAHSHRj5EQG9qe6Fb51IIygXignE9HFGtYdyg8BVLSjmMM
qnMuziLW1rsAAuC7itQYA+5b7rLsyGaGLy0kSF8fG2cx8Pd+GV4kbCVWrGrr0JzlXoBwZhuHVrUX
4Pd+jXIFhDm5aJzJNVeU/Q2Sr8m3Ve5YNc2ORKVo96Avp7CMP9C6eoeRLUz0uaQYVhKmmBvaI0XY
ahqpanv5pQY1O+E4voofQ0Acf9sE/QP7bZnDuWKSrRRBy0obSsl479scT3CPGdDznxIHrt42zpCp
nIWICR2t/miwtCXaMGqzm68YXbcj6Kf9ACwgIR8kayFB+hvOwFNq7MhA7Ihen/p0Nb6p1nEb/4GP
iO5bdhcN4hN6xdcxYyUDMv48GRgUL7KsMOsgU/pjTf37t/MQ7YkYkO19ToOJJED51U82EGxArdID
W2yAm8A13URYtZOXBWBDZM+T6Jqe/vx3aOqRkkMyizEDDoLMcuHhXW1FYttuI1orQWcN7cVTxUr4
KaKGAKFjVeTiKv+vcrNl89AzEfO7R79cJ6gsD/09FPt3VnD8+N2UkC30ashafK1PA8LWUtAyOHz6
vwr1psRUtcxhzvdVlpRbpORVaoJqkmPw6WEeEjTFuv2FTWvdE7hYAP5K7hGyU6l+mTEeTdblpw9K
DPddIziC4TpFL0plaSd/ogJf8nVAVmCOEjUl7OR9Jb1LjJQFtbU4f62l3PKwf9oE6B5zSbYENEps
l1g5OER37TvE84Pruk6yBjSKkTK1tMV1QzjQcNnxcYRroSMfIw457mBj8j69bYlLhOpnI5LbiGSx
zyOAspFYGw9JXB9vXEr5r0o/O+dIsTgx1chbuDL2zoXBwPdwdE5bLbrMUCOQgh9q2D6A5Dcc8Ljx
qeWj6TkfqoLPCi8Zy6B7F8jiDxFYBE2CXHGnbcKGswFMctfSd6uSpHKNFuRX/b3gGAwD3ub1LXgT
y6g4+GWCIi6mDN7FPqr27vMhOHhkzqQEdXwxIZJoua+7bxHmtZzMqa1JF1lXKFQGwGRvAXCuibMR
X6zteOWuLPXGUK3PE330zR4y12fDY1Q5c2JwUgrkuMLsR+BEnlL7YnQqsMGxcjb8Z3dwCOrpZ5s/
yqe7B/bCKk7QeTTEY74pXmiqmqSbBZ/Nxn0nN/TGji99wJrQf3sHbtvLzAQVXBDgovWVCPNAd7Lg
3KmUErheuRGKLxDxdBCi0xuKxzl+W5bwheJPuHdZpnBduiF02js54zlUHBfJTnQqvQ8Nih89LUU4
0yLWRn5B+0tq8uzVXGqVDcg9p7VPoqirYmIM/ISSG6TIISXoqnJPPJ9c6ZX05Elx43xULwmCYGSQ
eRW3HnuUkbWDTpuTICJ1frd/4oFJQf9ltCMD97aTPDjJT0+IGIWn0Qd7vj2u2v3ey80MSGfKTBSm
uuQlm9KAZNrEqBFMenNq9x8HZBvbcJwtt2ujkfaoOUcPhYYZ672KCHTMk+8uY0BRyK4UfZsiWygj
THtfX8KzVf6//+aIN6/yZTkUO67Pa1w5kZazhArinrP6ZxECqSpA34lPHYEWzurWGxZy1OxQENvp
algXXZbIkza8CrdBHvEYwKeRxJfiCYjwRf6RMIYyr+J9gNl9rgSLP11ssf3YFPMVHgN8FkZL+P3u
2o+YsWyBZJ4Es4flaS/+WZJ1GyIp1iTLsIEw7PCyVame3lRfK5oq3JDfNp4X8kbBic+Du1Zp1vZv
ri4mKYndcCmY3qSJJOv6blSoRlUm12ShzilMWcHIME5vx9n/18szDuDX/I6pRIm9/+P3Mwpl2wVa
5odSH1GEK0Pc85pr1jBeqAK77/Eswsz29bhUwzLlpbl9EdJBVYC9PxVzC1o8+Rv7T9vslI33vWut
kncBPQnA5mVsLvXgSaaDmlCJkxjh/+8S1jDrNj49h4dcYTDeqQwedhEXMwuDejQzx9MFB3Nzx9IK
YcCuxcFp2jF4mvhzyUXFxDsmBhnbtgXQPCN6ag+s/L82aX3TN2eDfY3Z/ZrnZBSntO972b0jPwjE
YxnB4KrQMh8tvQvBKHkltGeGvIcq0v+QeBqmQXxYTQpkK71ggPGTmuK1rfXkpSd2zaHTl0dUUeQy
LMBrTG/Z+581R/B0MUzL6E13mHMbmrHIg3UU27W5DUs+tka+TVl8xTMYbg+NTJGMqSN+yHka2u7f
tZ8JyIvgAOyZEGrdiEPiCZqfJbyKZsuWtJPKK9LgJyAZTH2300xnfS3hCortDVBCAkb4LG28eaNI
ZW7Iyig2cqocNbwVFW37eGXSu5I7eeeJ3wgNAnutPzo4XyyG8ZzVtMqvQUtVYLUkhPi0imMI44vj
0Z9SSr+x35jBPyIz6U1lzv9ich4L+LNip/ICwUEEvxCt7f9Ft1sZoG2etJtjVYeDAVwE5ofPxhyl
aAhRU3YtEwaAtXciU9n6L8f76bV7G4VI5fyVIL8f87Gr4v3ZDJP3a7u76nAvhAkFLz7q+V/eieeY
vHUn3hOWfZCiW1mEmAfHPPbiPIPJ+hzqIgh9J8TC3ymW+VhBp98SQq4gaZrLvFGk3PpGn/WI42Rp
AbzmekS75k6ch8QQqjqpTO3/iqkfrrEa0fwSJ66dKDRW0mjR5Rxs3zyDUht3rNqpu0vENpfmqsTs
NyvebQxfRuK5+R74Mg0JKKSabbfi9AcgRYvLIBEt/G+cVDbsoz6MsiFZknjpW6LD4WKUtjDsrJyR
951QrvsPVliC25nZ5EZxtAxt9Gzmqw9acUP/gI/EgG6ptb7h+KKpVrapuaB62PGd8XYv8hd7d7j7
e1hmEUwQaBpYfhUKON8xsXY4EEY/2arwTvwqceBIAsqnxemvK82PMpFFXx0Uf7kKDxq9XCnCV7TW
MyFVq53vcT8216ologrpLs/2vCYLeOlQgM8LBer48dwJgA/Ac7epJPMS6VJ2T8ZLEzWe+5woQbKz
mUxG06s96mnGUEKHqxyqlwLeOXnMw9dU3zve6huGeijK8B3tGWB7hH9s7N/3Q6vhAkon1kyHW29X
9BgAStzioxGDnGA00P+SI1exCsPj6o0PPaCXTIJ7O1COnz4/4efaQP3B1DtxhWem7KEosH7SBjSL
3ksxs1XrvMOtlmmfljHdsxms5lVi4YqtVkt/y0HSmldbBld6HEkisJWOwlak3n32tyWms/BBIkxz
eI9XxyZD2xAKj5NOcTTKeqwjsiGhl0E2V7sTk09jvu+CtNv3Zk78Xl5E6u7CmmEG3iAXUFc8gWoF
lLI6Jcr8e+AKt+HSlW4cUMVMZtvJxm7BILdPBkVXWV2xMF9WhfuLxG4ep/TeU8cbgG7enErr6/e/
CYahdYQBI8HqT7RFQhnn91G+FZfBHlCbpzATn5bEUrCfWXeTV9JnGv1ECfaxks8yLchbL8ZRLydB
PVPYx/Yx0QGGAYwAj0wKk6SsjiJnlxtR0LWA+ZGtbL6BMp/TY3YLYuGxMCij99x3xUA16WvV5+3g
PkbcJS9LSRKjOosyjCSlsLr7fDtmfmAYNVpUMBroOSQ21WFD2iTLmsJHkwI1ibz7gquzQmTG2LN5
AQf7y0hCMZrWU9VzFWVqyG/pqI8isVhzECuDW+a7rRxPySwTpTxsk43Z53CR0D6hAYseKggDM/KU
5L4GWVVqiX/lKLuYyFmKED7EbNDxzK4zs8K1eA+ycR1tqTPlrJs24tFnRZf1CuFmSg3h9ovDCD/H
lfSc2T1fJ2d+EETAjKzJ6TR553gGM9GYfXcPEU0/He1eY5/FmdlY+KzsSDUIZATnpYIE/yLrRR7l
su993LF5hxOL+eRKrSQp8aYpbfM59CaDEQIXTbJ4UNJsB45Zf4ve6Xvnjltn2XlV9Pn/AJtyDyc0
U1T2hztKfZJXfWUBwwto1OL6FU+TtN6JcWsfwomoQZ7SmNviNKDcOoshycZNJD2K/PHtbbU1c9QX
bSqZzsnTU4aNtncNqjb/lDaQsdnv50kCfGRfBDzQQfK8/8XkZivgpNkrgxJkCp+AZcv1+I3cs8jm
Q4kTJrkKmue9KbuSZjHqx1DkshOU1Rl3xOY+P+tNilpRCs9lFEuwv+S1l42JYuAiygZGhAov0/Yj
BVEQMTQ4IGFRxBGeqKMhWQ1I5rkfEQR7c06oCpwOv1+bgS6c1G+/Fg+AgEc2muvijqW6x0dRBYfr
xH8YKr3wEIkiMJfL4nq/ODJseFglwgFoTGPSuXzrT57lNlqQv0M5ov137yUjW6pFK7r985IqIFJZ
3XB8Db9P0D59BpnAnM+BrNbfh7yo3U02+9FDnDPtLhVVyRJqyHgQ2PaMONbklhpNE7RV7qM/6zuR
LjnTGtOQTu+rC20BUS5B5DFE1/dNxQFB580AgS7kIPPhmN/0k+WWaWsb2BAXQzMQjbS0QLkcJokE
3tKFNknhLrcwSSSR7r5iTXVuK18ibtLIkc3mliVjwOarxLdCzrryDWf6n8nQ3uHA9uL0wmRf7Ust
mTHhz5S4Pm62jIWNKXUjfKzrR2f910PtPtSJGwvbfJPJfvcmXMdItcHIYwwP+gzq5tJqBukst1xb
8HQIvHGBWSXGJmoxPjGDZxXvByMHF2bMVvS3JItNXXX/GkAeCaRcxGCf3GEHJwVrdQPo033PYEUC
byUsoCZNigBdoy/jyivrqUb4mNmqS3UZdcwygcqyn1ZFTvq5kCah1rkgEPITH+pOvLs9m6xG5gQZ
Jrbbw2O5xX8inDTI3+hftCVNL7LxDLaOX589bhPpeaybIBRDmaiqExaZs6Rumz758SlgRp6VDXnZ
OlhLfmUUmAO++ZGdJsJne/MTcjSzA37e3mf2x1k4F7fFXCjMUbfYG8b5qsqOrUlKgO81M+9rsLN+
qr9dQZB/7eWPpxsAERzNlmmEHYOcrGrT4UTqh6ZSpljZ9D+qy0ubXKZwHKfHoitrGHjNwfKv2dcu
yE0ujb7oXv2PRpdUlR/hS92Fx8EU50EKYBThzCKDUBPojsffXJOuK7P3uNy4wjNIaYak1mT1UP6h
MiOaFPXTL7Cc+SHT33mJ+RLZem0WsJFI/2e6DCHkyD3CDKbfoGB9xFSmGJGa2em0srZhi7Ik8KLO
5wdDkn0Tb4qBPI5fHt7SW3EYWba4uwv75CBsf5zhC8VpnmvWC8DGjxZV+YsfQTbUgzp+r62NhQIS
I27MnjT/Kt/hqJ8apWvvUQVDnhs6j+y9+i+YOcIivRBDqFWig3je44A3bvxka0KBkR81/iO77Es9
EX5D1LFDVnWisgGH6hgGY00yOHLT1eiqhKITqtBvgTEIVUMr/BSgAMP2y8Yo0MU/LKCOXK4Fhb+H
tOcjOZVFsJzpqUvKsneFXUZOvyEscwiFsigNIQp+Wwy7L/LzU/Db+yBDyEEwdbI+cGQCrXU/1DkA
ckx1dCGfFYE41uf7Iq8Q76msfWDnzP+K5ibituPYhm8dnzTI/zmUgborNTFLNKJjqs98ig2s5PWo
soi9wE2JO8rqNsZhg1K/CkNecpIG5SHM8kjq55X+zcEDarPJ2+t4BasU6H5hJ0Wu1EAYn4iB+w7N
aOHm0kPqTeYStpn+AJlFTjIaknv+My63HCjQRJqvNAPZeWed2t7oPGfukyvEb/IgQ9P/hxG2/lOr
egFiTEKT4tQA7057+2vmH59uj+rLMrWIIKGt8AemNcEyKqAJFvOwHwbE8RYc1gmfGvhL8Wi+9Wub
nUKFAJaxd9j9yIDd058nWSf9yp2VViIVBJDNaw9eWpu+TbXWiVoFTs/V8FETOOVqfEZuvkXrvvRi
J57eGW7p2rS7BxY8enVvUWai7BjKF99KSDgwirDKi0Q0CVaEZZquodhV9Z/x/eN9p53uiASscNGz
rITA8gHYUMfoDjYHXOChakBTlcOGVDU3S3UpgXOSQtiqCQ9UtAzbSheWG/JeuOngvu4PBzWz+Y1w
DD5lQwwvAQv/wsn2Bch/GFZ8021Ebh1NFGuIr8R0xyuZ1Ys9X7FB3YfYCAn1kgxDmeIaNm1nh46M
UMqBXOLF2T9c2H27rn5KC2qy7dzxNs8JdO4Sn/+LEKO8GdwlseSf9tKDNBNDHIoDcQuNECOkhX+6
EOxaisPi4OVISGF1iGyNKVCEPZagNqb0DeKM/f0nZL/gCZsbrbQuqgDs+IZdKJCeoMBJNS3cFgpH
U01PCINCWQTGrR+apjjZV/bjkkILZiFK3A/pkl/AvxJSYN6vZ4PZh3spOmP4F2Sugv0z5aAhLtFx
ZUAW6JLxiOlExiKlZvVIorMpnh4uSwSKdcK1g/rNHcvF+b/l11YXqynpBEPoKJATZlwhy+SITl11
YRjVz2l4P45Ry8vTXy8EcS521vSOzoVt8PJX/+N0Amb9fI+qJOHgXCTxWKLqOH+uGf4MuGw3IqWR
68MmCuIisNopSmbnNmATJEcDLp6XuT2D4QfrUxTqDcf3sD+flkQQyO3FvdZD543xh4pzwTF7nFu1
C9aFSRem02ACV8zXFD7ilGggzaAnxlic2bWJ+oxS5/YX2/wPwmZhO70HqV5MoJaEvRCrA5sxfq8S
wdSN4C1dNX/nysCklhnMn4CubrFQZK6gisvjIUL0MIVV3Lvw+GcSiUyViGygq4rRyAeY/LZsBr5r
O1HpDzmdhA8wtZE5UUV/xJOi9YQ63PyXAB7uv1IL1XkhmFrz6K24It2dNipfhjIvZilDhflrpxbq
UrS0A72hjylVd0/lrJSVat9yzX5MzIA5rwa8MlFTwdyRgEoAz2PsBu8A0FzCDbYe5+7vzfyCqmcN
fAzF+n/sjNo5DHBzzht+IMDIjqRc3VOg8SNRNtlkfKrCuL5VwnMs9F/hSWhPzds2v4mTsydy9F1D
Amq6niQNpgmv9mBL0wqVPJxvGJdQe3kHBBMmYZlugXWY9XyBOqL17OPLRnhBBBWIjspV2JX6riVw
HsrX63KfFVzPWjAQtKkBAkMqk8+c2Ncp6Eb0hu1eHCqDcRFpXaQ07Zz/G5E7CXAtJQF8RxmYZNEr
LOePUkhV+zlDEtzsTsU4qRnTCg0b+n/CniIVmDuJqqHanDfV1nkgBec4iQWfnFOMJC31vxXJYs2u
WfPvbsGSzcD7E9zmc3JJtq0EIWAsxLyNeI9itKia758/ZfGpn0ts7mE/S2lXbZsbq01PZ4H45o9h
6EWKvCvh98H6IvmpnSMT5uoWAZrI2kXZ/oKJ7Urzl+S5yQQOeU2W0roQB23MgTi+FMcVwCG7O/XP
bh07kHGliyuRqqs9wZE2sUPgpfzxPU8XyIfZ8B/LC8RCLgqVwa3PmJGFBmn2qyzOBwdvKKvJzqc/
KlMKoUYtojzutoBHYxGN4XbJrwQDjPTkGfA5OpySd2IxvdmXAULwdpXVBMmeBDqCXgEMdqbgn+VC
mL5szpFX6mxTNmzdIRqub7CtTrIquv0ttbeZkEzJ+u3i+Lu5FMyfZ141SZ5uXoPSdvxxci0+s4BT
MCE1axhRthLKNdVyl8u2TC9YvSS5Boov2ozrWHdkVUpQpHbWOn/wFDJqFHbYBMibqNJuaZE71riP
cxZZZgvnXAQOujOAu4oCkC8oOtrviUkVrkZRRYh9CfGfFPu/Mc3PB2kbmwGwzkmrfDyv2S5cVXPv
10DiX9Qs9TpXLuaLQHiucRnaVTKNoFMs2FnvMR/y7eZGmroVsWk1QfIUFfIwUWAi5i2s36HyPAlz
W4aYW/co1psv35ZndXbT+ia0kiAb9RdjOHuZzbCga3dwhY8MjWvG2KtHbfj/DahE8CIVxiXBpfOm
J/Juu+ad6ui3uxy4PtTNNLqUhOw32WlE2b3BLMRqMkGDo3D9uTLvMNHHa8Ck9C8O/vLYmxmilaHV
oNVt2XeugvGrFPCmSxFrJ6mxU1syjPGwCI7GhvOEnazP0zVqAsilI0gJCLQi/UdYLSLoRkfOvnpx
l4x7ELBEFvNqcFmgu5uAIu0x57GsghVoZBrUJOeN32p6BU5LqiS6TnIXObggci6W1i0p4FXFOwXD
WMGkchW+eUBpG9y+KOYyQ1iCseaovq/+NuoFkQPv4o5PoprJ9xG8M5orWo/Kl4dEwB8MeeWqEMd8
E0UICnB0ui5WjeQ+cecCMNtunw6cq2mxGyXZl6QZPau6m4ToyD+zW/o9VjYxk65EPxd2CQg9yCol
YGiDuhgD6YC5FgGdEsEHV+NHBo97iOgTd10AUxIa++M7fqfL7bfddhoFLsTXy2E128SlpRQ/1Is/
dx4uQJQF2FOGGK0FAm0Q2uRs+lcQ1BOcGAztNMdkKsly/K5v6tQuz0qpDA9LO1/wLQBLdNLqBkUs
1NOSPO15DRp+L9mdMm8NfAjISEaoHQN5nuedorlfGKFWwBVqmpSdpJ/iikqOFsx+G691EE/Qebtd
Cf9/6b09dtS8BZMtM1XMGRfkqmEUtu9tUt0qNpAzvUUOFqsYdx4qOWhFCbGsUNK26ETXD8fqlPRQ
+dh7w/0Fq+5MYBaamzsDyfi00Ez2HtKCOz2V+ZNqfy8yb/NZokJM3sKIYwCxg+kx9DRLUWQYUqcC
AKa8sfMSckbzqbrb+0vOreoPtXm5uvb5oav1+lYmgoKkOeM0A545QuDjkM3252ZBEAUrMBPxnoNz
d7wsUcytIBejrhps6hto/LQTvSs2fur9OZlPkuqtK9HC63kJVa85w86GkRZEd3CozT/hn0PL70he
7fKDgR3r3VsjD32UOfOpH98ivt3GJU4eKK5taIME7+jpCVKqkjIUqtqRbk3GSh87FJCLUOZwSubD
px8fhvE/IHWzb/rjJ+qOBcub82pYefG8om2hnLmteSy8kKKkCyO9RCKCkXV0zozkmA1KHkzYvLQu
stoPWbqm4RCRXksT4XFLDNz6Z1zvzJKF97bL89KrrWfKz8bN3CJA9xCInWig7A9GxQdAnmDXrbvy
6paxiDgK3y2B/873yC/pcOkum1NqYw/KpeFOit+qQaTEAfu4kUHT5rOk8l4PQ7AGTi7fQZ2AIuRP
xHNdQiQva3pBosB+P4GlVDBM2RhdGEjHp0AJ3K7k15vaCe0Bk/blciIgr4fdJg7wBlcokUapRtuL
rOyhzKaip6EKMDHK2tzrj/hXIkgq3LZEWOs2WyKqa+xpnCP8myHUp+o/a2XPFM+Ztw/SV8h4ZIkk
xvMOkJSv043P325titBRyD6LO5fjX/63FlaGDbLkTg6i5Xc2FFXYtmcucjF7lLzUWWv7SdLu+mlm
60x2JzkSJxDcQsfrHkEjPcB/qAsM1LPYmzV6bS+ElEEFYZ/tfaQLoi12KgDmG6mWwDC5QjxZwIk2
4nb9WYcWNHSM1lhU6mAhSzKm45Uhdh7N2h5n3ngj2DjJ1UimqorX/4voRbFz1SQS6sjiCtyvn9ab
WjK3arX1zqveeaKw/zBURfEMIAq5nsmRn64oAw9JSW17Cgtkd/tBlFWXhLNHCXXEVKb7YSFJCwga
f+CSl0dnn7dt8DOmUTPdPLiRtFKY56pJG53nBWLJCAtiqhs01vjYe7NPZnqH23EK19ZugkI8msRM
89IUDMm3EkBFxjxjw3bld1kOWjYTtbcrVoDNO3gzrGn0WKq0A4UHx12XTTtqsIXlKLtIbd+2Doj/
W7dYq/t+Q6IUFmi8hzN0uXAQqO9kcfZO/PinV03hs1w6+K/eL90zOYLa7jKxcrbDitKrnwVkO38V
ZBzYTyivKWlvMKsdX3eXlUHTg5eR/FBkwjutVu//wZNuQNyJ6Z1bMTToSt5hQ+/cZaNtPvLaSfoA
4NpRJ+szP/t1L+jQl0L2V9ZhrBxgbJEk2RpnSUF0I9/RjjR5N/AiMhdS1Htlku8UgM2W4DD7ycf+
lNIh6EQsMoCEdT6ndpCPXZGImaM3PWhEmyeRX3458QyDQz2ap7e7BhXypZW0j/zdjlpIYJI/W6wb
9AG5e91jnmQRe+FrHaZNZML3I7YtYQmt985GZoMMaQTHagpgeBNZzchPp2PijfNz6aJnajr7WXfq
BnkEXC4Yl2jqaLlivkbZYa78d0n8VYSsqk+8qF5aRY3FS5buf6gofTyMv966KwqDjYr6YvvzDzHM
I5GwbMCxF0BgCwqztvutUj4RkNgCIpq/ioQb2m++xeHO3VBxxXKSykSh0CSrsCKGePSnU7HoMbYz
viIvfWax3OV9SXJBlri7G8tsfDqnR9muIiEElD83exDXVnhZ6i0lY/JcHux/tEZqRFqgDUIGX9Py
Y8xe8PXo3dAhzIn2/Boq/7ILNP/XjPnNCFdCLwY8QYniL/3X0qVAsHi4bCAr7CiAhOxY/QyNe+FV
tnb2/68/MGEb49Kpf5j65mZLNaO6JP3haCqQYr71cltCkM2aYJg9cirZ8MWr+Nw/1jHscOAge4Sr
ITIE0gvdGqqeK/p93CE9eUT/j9+2d71iwA97CPnKXrHWHAON4r0NJWe3x1c6EVMXxuZNjoY837sO
i9iV0oTaXCeO2LGSGo6J8+ZI6sQkLnjMFs+LDpXbULEbBFPiPz3TIWyioxofGN7NpcunDMIOURUy
LMPAQQsBX3LVQXkUEUzsKKf4MbbTOOPPB/Fkvt24KzP7du3NQ0XUaD7xCyGPNx2xw7u3Wz50yzeY
Sn/iQovG8AZnbn905ou1pZaN0u7Z4VpKUz7bqxpc80Ja6ul2sOZgbMLQR0Cth1nQB4o7yMzYGvVb
y4C7xna2GLSlDYxyfK9yHVywXDgBmTziJ7V/GjCY2dnfE37R3fmGCaZLdMgRNHu7O/KFXCefyaYG
ywzD66HUCi3GUIm+GBwanmBXXAmdvm3Cq2owkWrJYirmCLb2nQsxfU0CfXi0EsR7DeG4gZiSuQGb
MOqvBYuq4tG3qIjqWh+oVLYdiDXaVLUC/HnrItGqMPBZQMgVDHCO12XD3dcjK2WVVE9aVNgYs4TF
1Zq7EJoL0VGFMjNgILly9sFGdtZ8PZdPXBuKg5W954toVwTOa1WdSFRiuq6wUj2/ROVBS2wYMWvC
FYRL9DKhLpikkdV3wV/Vb39yMaf0e6VIEejEVEpefxFO4JprWXbM2NPWRAyGZBOKHJR8kfs0n46T
IXj7apr7OsP2WolmrPG5dd3GZx7nhEjEqcbCzYoMTrAvrwBaITWg0flXu8zNT5Eft676nxZe5o33
d8ZzAcSEfxDG5c32EIvCnsEvdFaZXSLtR9gkQ0kpNiKKN/o8CpA5Mx5i+/DN8Koy8okVRJxYlVh/
bLNrwv3zWL1r+fYnhJv8hvfjvc2MLPKrUFWgu37LO5Y0f+VaVt2THC8crw2+CGhsO5AXA/UemTWc
0OXGGUz1RWVHyhjfA/wtfwIU6Af5MPrRaCxUzacWcUw9HAiVfJH3n2cLrv0u2918MHGOu1PqvCeK
2F/EPKg5hp0YeNpuOtO/ajL0Y5mInC1FGmjJ+fMVwlanySxlJKuiG7oMLZG1zyRe+vDh2KGUiMTK
39YkmFKya69dhYSiSytpTCVVbUbehjOo91+FZhIuL3ad0Aj64mCYVycGF5AL2iynS9kUJyFaqG9F
gwLfH6+pprvsxVSKVG9K6Q1CVBlsZLWY3k/wBLwKC0GKIq1dmYwDHYicErZXxmhu2quhNPoFuaOs
LNmOeD5BHQGgnJpFe1ZsisX2gS8Tyd5du5ZGCPRcD6cJNq9oYI/ZFsY6cBGvxM5q3NKN4rr1afb9
sMkeFpBa3M+wY8vGd/4czhUpit7KotqMZD4aCoC33Ocf20sqxnPQq/IKk15wPW3axp+8rveTIO2Z
7Pt1kAX3k+Tq5IbY25qsyL6S1fxiLLWYCutA2HiFAfK5FNENt/E73Se5Qz/xwE0e6FJxWjrk7kck
uXptCdFUjx9g1/1tw4DIcXxLs8UiHrT47rQzuoWlUtEl6T2PX1kHUuRLEjA5tpSi9YyqUFu8/nHq
BsSARMl0j/Yjhr9f210cMtMwtKGhLS0RDWXQJIJnvtMR1dkKv2McmcFeNz//ROZ4bpypTBlyHp7V
vO9L4NpHqc8tHQkbk6bh3xdsaRM70ePNaP1jcyYv4IBINmHYl/lG4t2J3gY6TqgWud5q9kv+lBdg
S/pTPNhZalRFKBSttUQWyzont+soKSizZJzQgqvNkv6V2okCDtEFGVwqBYHH8IznfimfmNoDND6p
8MZPpZPNfWWhXR49cCSKjMPmd/96vfvWUWS6S2R5qshZjcVtIzBqOMTS7Ukj8gTvkUQLOnUJpdUl
Th+qegj3dXN+Hv/hvIdQ79cFLHmAf0/hPohqFsxOVt9YSPF5Xujpb2NbccUUtaVGpNftnCHu9yFn
QyLM8rdw4wBkl9F5ICevsQEwUH6i8PYKcEp0JOaad6y4ZTCSsBaJS5Rjm3VSfhHPn8K+E/3IqPIB
9xAp6WRtJvC5J0/yedSHu2zsZcToYCoUAzm9GNHkjlahh67YWnBha9Qy3DEMkIpyy3NQFX3a2y/H
Q3b7X43cWaXPMecX/JhcB3ng/ellMjSv9wFlt5E0rP28OnmLjhwALIGjNJK/quk0kD64Ksj1mEA5
rLOCsUu9r518/u/lhbt1ji2usjOdP9JCBo/hNuDjUG6kp8Yt0yuYuFed77savkHL8S0orIuBkj4+
mJJxeCY+LZTG7rqNbDC7xeCF84v+inrvrE7feBdt0h/YfvwN7euKf72eLiOoaaKAXPvsptFYfmAJ
gK8ApkJUMumxz8u4HOkkK6GIDH46xb7zsLC+DWXsXPfYC51QJxjsyQGG/d1lQm2a/iDGSdlWMALp
w1kQuuK0Bm46t3syV5+4pOHZfKHbq2ANcUHGSx2h+7ggxmGTHzssBA9AkRvKhbQIaXfWi/D+pEMB
HZVdqmtEOEIaqdhL4rY/tT69c6MLfLeJX2d9AduS/PzQ/3Dk9zy12MIJzL7ks/W6SkmlJn1EgmZU
e5cO81v0OFdoHE2hZ24Sw2R0t9UEnbs9u5goLJVM2gpeSY7oT9UxMmBal5bBxXf2Udo7avRnWF0U
OnVg99++HpFSqHXd7ZRhzThd9Y06hbR4bvUD5GCHv/H3zq8pH+mHjAEvdk3ZlYOi8emciZgRO+Dq
wgMugMs/YIQd22n9TW+sD4P7BYJmx/jvQxxiOKad6prdBrpTl3dvkkHWOifVzAHafEZO1gmYangl
Xv8GIiMPFukYLUnWQt03e0kIP3ePl5fE7kLbmdGSwZs+709pSAiee5bQY9e8Gi/ss6vICE0ttMWQ
KSJxUw5Biq6C+IOAiNmVHI0cOWispt8AGclOxC4t33FZa0v9WZjcYekyw0IsijN16hUDp09dPvxq
kIyuLLiBDn46uN+lPdr+EhbSLIAsbvDnJ1cZ4qAHALdNgpeHQ37pbeJxYM4qtkE9z4bS/NNTV7Lu
R2JW4K1ay4W1Dl9glgFUTxmqn2tA7ug+AgbFWV083smMaY2AuiSgoEj2Ri6XbKilN6BhLVtHJl2u
azPj0Pblmxh/pJYynIiholCQBVU/3tBFWAiXFvhsjdm1UkjLrPflSbmGydhm7xSc6PDwKX5oW1ro
fAO9WxQMikLlM4JaFcyPEWin3Ma+fWSMZYVrM0gNUC1jPiM3keyyw1CdpZLmQi+hd7Zx2v5UdY98
kT/yznV+FrjiesZnty3C7Cmckd8sBCHKqDeDw0kAtqx2pRWNSIFjlXmhDNkOZS9Z0nYSerT1kASi
YUYbAk79CWKIvLNFGKH58BiY9tKTY6UmLg74L9aNbBQM5+D9fXS389Ic7zrfAsZGMzoP34+zSlvI
F8Rc6LasazfdSiU8T1LSmy2E+SozMXrTANS1rQVT7Qzi0a1ZaRwsjtRUtKZdciXiNMqFpv31ReX1
2MCjtSElYAamcksOmneWE5cL2gR8KF8TSTZVRe7k4Maydt6IY/6dujvJs0mRnGEu9/ge6GGKxaZk
QwpKErl7FMCMFpaG1Nuj0RoEVWBw1dE7NREU/eAaNoBMdx0T4Xc8kJF2SYotozzxtv/kSXdd02Jr
StQpq7CtRimgXc88Kkj7NTuZ6ExD1txAgXQSWUbLsdzSEpb94zYQuw2loHPmPSEX04FCUinrY+76
dQ+yNc6t86rsyv9eEhUlDgPdhJ1nJNZmJATxYrmLAGVJDWKpwFZx5k9grlwIi7qyJV8nmdGVUGbO
W0F4TsvbVo6EENFOUfeTCgN2PhlXe6JCfw213Na1UXMgUgypaMYyvuz2qqlVqGKT1JqmL+GVJkKN
KrSzwkmgSGLtK/r/nNpAI3dPgW3NR8bYxH0u4FnMfX/IQ3TE2nI9IC7wcnBe/a4jeA5jaH5IaLt5
RcOeTQlvL316LCX5w3aZ7xEDjT5lQBF0GF9SaXRg/A+65JpPXullNKKwLV2KthgkPVciEQ6d8xn0
HWM3x5YevBkyk3wcL73EQTN+zluND0tclGaV1cjFyhntsWg4VCGslrG6oi2bKbQd4oSi69v/ULXp
p3tLRQjjIxB7k1Y+L2Xhm4dFNjYUtc6IhkB3NQXr2ww06msdcFiaHB6QxzvEfhlXS8H/Dmo0INMt
677RdyK7HOta5GVVgSVmc1UzY8uWQypFZ/N+ysd45z9vzoooi4LSm5pQjmoKraQfeQUNLpy7xyg7
vBXzgJ2FfEE8OXRwPRpSDtmpmf2gsT9/2b+pcE/acThvmhfxxJGAACAnQUC71HMTXpsxgKhJT3J8
PcUMEC6Zt17YrUE5VtVz2OVsUUdCNAT7Dwl99sPTZtUUdH8gV2gxi85knm2UTgCEBsc+wdJaHFN8
so0PeMqbfVgovxZdJw5KqB1c7lkokk3KuSz5gfg5WWEcibGMENo3KFxFARPum3JhUx5TKncbdjwO
9XOrxB9tsg+51aBJvmvhwzwqg6GYXCCxh+VW0Zuy+waqY9YCrSbrxAAfClIFqezAg7yJzeaLaCK+
J7tcjDgK/OS4CSVU2D4iuWl0kVFP1Zg0zzwx//G5j4N+ujUS2l8BYS8o199IOxrk1W5+o9NkZW5m
C39OVNFPELTCJ0JPacE3k4WCwPhfVh7HecBsU7iE9NWWVigc3xabvnPPrGGNCO01byLoaI0Jxru/
NoZIjpEIOl45MfxrckM5jT4NESWwNtmyxCumEsywXZhfd6y7+MXRiT0F1P1U9UGnAFNgNwdNue9v
jkSIBCliYBft8mAdau83CGcWEUANUMUmr3u25Jhbw7JFMFRG7+pjkJkZBapvHLOl1UZUE3kPTUvA
NHhHJCZtUAALPlsPlqQ4l31+CurYPXOr3wASH9xCPvguREc8Rp9xfBCf4xoxkJw6mznqVOqt8LwA
LefFMxdEi/hv64LGr1UPp2Z7snfZeVn80W3tDq48zWh24UpiKZsJGr1qh5OcuViN9Wia/qRAKxJI
czx6LUabSsqdtMQLg0Bs3o9KEadvXTTRZEasl7r2VN1AaoPBPd/4hctu40XOD+uap+4iqbWEklFA
3/BnlB3VkteWzI9kcAv0jUdIHyktKBOv8En2+jtJNYdL1sCJDOYnyS5GfeR4uh4iyjV8j+sLhZN6
W2lRSA15yGfPLjbIMdQg9MTQRB1S8tyiLGo2LJcYJ5x5/cKip5PxeSf0K7+0Xtx3rU9vzaLVvFJw
VkSeLsrMFH3DLeHZp6ZHZ23nfDI+sCrntbAIleu2P2ZEsF4Agvq27vqPkdst5TQDvJCtf13b/nuH
JOCdhnaLYRq5tIDWhQ64iYC+zwfGk6IUmpsitrXqZVM2PZaBDF6mLJ+MmoIfAwBk1RD7VdihvGBi
I5g09/lfpRtptJ/l3yPY1BAJ9EcYgXFN/8rdlKb/wHHpukcw99u1w4j3R4+9VUdoyXMvfJ6e4qXh
Bnjq6zGeFjAhkNBGM2a4vz2C1nZtp3Gnv36gtba+cysrAt5jKJrpEE295GznRVlp3ET/IeV0OQhy
0IXq7zlTYxp8UmWJLoyBYr1axu/rCADbxSEVjLuUSwqFbt/7tVhjHWzFH+LbWOmTUQv7UKJb0YsY
RllM/mi8lJU/R/bc7hBMNgvbZ+aM3IwCjgx7rXlLpG3v+m8L+Qfrtv7N3kojkpjIiUs4J2Jcs1g+
nyMIZ+IBnR5GkHFGrOlo9ke/uutFzIC/4WcN1unw+FvlyAmvHMKGOxIk94uXUxrIq33EYxy060Sv
xSemioC/G6oFYwQ/7B4KD9vZ0H6jumMCWiiTZYYarh0NN8f4rEEfTFbdcfmLMIUm3R+yJRc8T47/
QbWxAZav3po/hxwew9oaITPC5+jFrMkAWEjrwFnaH7Ikhi0qhdIarL6aIF0JXhzigTjrKoUD99Jw
XgJGjjF3xOIuFdvcUwm1UGLr5glTtn6xxf/K5j2QC2tAkmbvsHcXeZ+QvLBWcAVttjwQLvlz9cf7
KMzMWE3OqSDLSqVtWXhF/+7vC/s2RfCOy/dJ4HLnTzhOx+7eF3Ha3bufMFkcI45m6DXrUiPoGSc/
SccL0qPZdgRNwNbcGA243CDhzNivKbHEOtfRoI8S2VlhSbmH8oTYpkrjgLXPEYagHf6Ww8EvZ+yQ
7OxMDmrVffPtk3UH7zPaQC6dBH+DqS1sUzMBK5ifxYX0w/jhmY2yyqxnHSmx6YU71yw+0cPyJ4hM
LHVuE/f8fxL/FwSFI672xJJRdPwsdHk3HIrfpt53eKalVMIzQWr6zeuwFiApSvbNV/ohatOqMwD+
afjHQ30lGPn0MmB4wk/lApSg79swUAtMP23iOfsngGQ6HS4GTJWYmiWqVMSVF5yeiNojpxpdTaU4
Je5zVM6JuRwBhJk/HQ3rwT2G+qcd8wCK5ji80x/0ggaIb8nW4/yic90Mw3+s378LP0ej4hmqBmyS
Juk6Q32OEVhyKO0G/s625p681jI7zKxZiAPj9ZPSvBmEZkHzhTYMfiP6Su6OUq/gm0HpKapvI5z5
HXqDXOofoYlrCXi0n3wxMKgw/TB4w7yWcvo59yhtHHDXyey5zVflK5qkdYOjfk+Sj2SHmHosF62G
KGBMN1VnBmnccU3J4LZYXWR3uVtwvJnFp8DzVvh2HulLk1TTRZuMZ76truYIaP+qShJc0Ls+v5Lk
8PNjJMJUy1GDVBSfYYaN0xNeP2QmjDEUlaCOAg+Q9vp4LuD+3sZZ6jfG/OODy4LGEYccFEG1QfOi
2RqG5SsplO5RuWA2aMLPCh9ySGWJ01KWjC4FRFLJrs0j5ODuOp9lZpI4rCy7Kl6uBC418ZUgmJ7G
XKz47/JUKvkdC+0M5mURR4QoudiG7jV1N6hGtNs45toch7LFHsuZA/JMcOaA1kkSuQgjYbHRzJxS
yUuOZFmoyZOj8pqgEn36cDDgqUMw9a7hZFDHQa59BBgA5ckkKMHCLv1e6rgMlHSFeUhcz2oZgrGQ
wdAo3V5qTnRgFeih8iqdVt4p/7VUD1vkPEzKPL80KgL/ydjxmTqVqZitAqtcE3JRz0101TVr5fxx
xMz9C7K4wke0ywsuanbyUewJBo3oqINBM1Q4SrAdL0t2C1W7rOi6FkD2aSNMM12qF3AIQmNY1c3Q
d12GGSPRVjK8LHmzX8V5e5eqW6n2aUoEu20BfbnOxwXz9EFHy1EuT3pvgkxLWBj/kz+7WVyzn6JX
k8Mu5KQN6ynhZfCwxfW8kjaMOVNqgriYFhSAjBIMddh6iCf1998OHGsxDLp9DfmxlawPEgKWS98/
CjBhlDzXkk3k/KM4n02W50mTaTJf75tc/LOUJ5d8kMpvgLUt+ZH9PFErHPUt0KHg3j03tUEuNMaW
mxUR29JnYQIW9NoJJF3+TeKdKMEkw5zYPkR8oohCEIXY4Z3aLOC54nZ8S5bXoWNzTbEsLH8spFCo
69ww7adqo1Tp/TWNwkXFrNVX8+CxBUpg3SBFNK3gjU3ljhDWhrkjIXhbrnTT7hF5ZCvpghcmliz5
9mFH99+ZwSuU7DtgXe3toMfHAPXZeK5S029GeD6aPvQ9EEJqRETzWpTKG1GVwTcqwlg2N70U9gtz
6MHsEBYc8TWQUiBW5v9d39/i2u5lFXCMOgVYS3ePYJGkFQkKqbgQxXpDkZZzKFAOZo78J7v6hIMA
HcthfoTUVNCXy6AGo/iVwkphM0VCxaEg130JZpVTNIyNTAiqfk/EnqoJZ1j8ziLjeyTEaXPE6quF
jxXpOFtHhppTYduSvXLj0/tq1eNDZXg1DQFy4Q9eC3OvVp/3R4fRm/MOXm+nETxlmvTDF2yoqHJ+
a3YTl/rst0FP5QiU7D7MYD7km8GyMOPKYfmu+5aNr6gD+wYdOz5/TBFRpFE4rgl4OCK5dQOL0XIZ
aoWhd5dY14lNpLUik46XbiK+7ud0b62a7CZcDEz4paeE0j0eeVd3EvUCFfjqYgTZYV9JB4bA27Hg
+NgVxM1FWhHEtd0NzWoVL8rE4j5k/rxiwQbYBOM9dJuQxZC4FJFD293RGqtBSz2bshxLciadkc9v
7V7jYFfQKvCz40RwdXgdMbfX1iZmM94B0O5uqfN1dM1XBAiGk/I+PoVh/AVEsbIAiRHb10hZFdPQ
igfUBaTqaibpQq+50OHtqUQ6xcyGxdv2wKDrFNwJ31WbKcLSY7OdZQi9sTVyUKCkq/j67mKJSFD6
tcDyJRr0hQdzlABqRvu+HN6f3gR6yOOMrBbTCauX6AGKriedOt6mDuZR1mlHDf0WrgK5of0P49UP
UZrxzUTdfy4OEMJf5tscCrsT1s+lkE46pjhD816TYGhsz/QkYw/+mrvXFwACd5as4uqE6GPT7Lxu
iRLOqcI+8F9WN3fApu+kwTMi8zeNRiwJcGYSue+1JCSRZof0be3XCIIisr2g38GzOYyYt9UeOP1o
lHzFlqX++CO5rW/nJedUpeDzZpR8mn91pclTSTuKhOqIImKRgw9HDNi0c7BK3ei6lS6kxQvVvDZI
rg+lZweeKSRZe1EMU0RDuXjo5NZ86wHuWopIp4OElFE4z3ZBrvN3Cyzw64x+itIy1RoKTCOMPIb2
oQmlrNIai2xYt0pCpHKVbV+ecymxy3W4BhrRtOOTf4+ntmLNHI5MTaHThQ1uxopkU3LmihsIgg5D
+mWku5YYP8zyK7sVfgOjYoS9OGlNYv26RLaI4u3ycsh1m/X/mDagahE1Th7M6VNNzWGVScAn7OP0
PIXFBZs4yapTGXsiDQ/iUrc/MQdbnvLpUhqIrzfHtv/cMfS9O5gpgO2E3T/3Ub8bQReR5O4mJL1q
yjq2jY0P6cWe0ig+4pmfPAwRZKU3QWRhOSBHXptrRGDcMw5Hk/0yx0YWs9ALz7P69VPfo57D6VoQ
F7tAnVymbdoaIsL+9K5lTME1JkWv2j9sm6ZWVsFD7dv+UPxsgYzAiQl+ruf8d/Jr7WkoLWadqT5m
tcwqh6KXpgfolvOMLKDEazowfs1jDMwiaEaiL391hwEZLD4nBHw7ek2NeVTHHoG1yisxcYMKWkOT
eNVRNqfwYDXjB+YTeb5LQtxZIixtOmjKajPMho8LpmNG2bSV5e5qA2uo/zsA7IuwQ/EBtdpIXerJ
oMVQy27La4SWRxoJ/SgkoLVlLI3oMbkF/itQqKRRLABxd+eVW+8n07vMW+af9INISDxPhyo2EDCw
h32z4XSVbVRXgyeKOgmyA3/SJaBN1Lc/cVCMfINAzibbzHa8M8RPrRcx7WkyVIde+HRJYA24CMKp
Nb7Q5hHXOd0EUojRBQJd5Wo49uNGJZ2JhxKQc5I9JnVnF8g0D/BZh/7qVOq2IoQiLeXoM+ouS0ob
3caGLxzPOqdQbCreSCgfk6CRudk9JJYLZUTtyPQhB6U4NZV0SE+Y0UWXXYZbTOf3P7PQiDyh8dBu
J8v++eALTwnGDkc5jQXKeo3boZpoN9G6GZogJcwLUFAfwG7CXVcx1GeMvlpE2HyfMssI9dY3NU1l
VVOvY6kqqVCQukKBS7FJrft8pVi4G5R3fUHg3zetJ/SY3epyg9x55stMbDsIQkLNw5W0pt7TkyO7
7nYyYOPBvYR9mFZWbqq2mm00U0TL7A9MUHNDh+Zd6vWffVbOX6GpMxozoVy3Zf5tSheqWtJmCOSP
JvwV+P8IQs9ECuSc4mtqqRT6nD0DGv5DbHkaq9R89qj8yfR+bTrZna8r/FaWuVBBFF5Fu4Gnub30
qbWFltFye0Y8xViiu7Q6fyVqluqOroijLs1opJ6e4pJB7dHHn4nKqY3CJaSCYNIl+KIY5WjSxRen
nSjmNo1NLfB3LVnSSg7lFuRmXDoqkcZcMwU/JXXbaV6sxyaa7J+aUks4HoCXBcgab78irJzCgjGH
M0chjFK6EJVt8LUIjf8LCwheh/xvV/cLCMYU0FaxtBWrJmn75k4ienlxuCBEH2TbrUWcpqn0BLV9
HJAloSLZ9eU72ynV9U8/WTdpKHMh2hto0ym4G+7Of3p/wW5oEJim42xEqpMvDwgSiT+Ob/OHsWBL
AkD5+SvIPYa/apwMYgq/uYauqdhVMP1h0svxPTz1v2+oU/z/1dq5jcDh6akFTXA9vIhzTyCxZzFW
dY00J8S0FpUFvGNw1RbmqpM3KPS00RzXO55AHKzFy/8UuAeV64pZoU7a3NXN9jIJpv9Rnc0rtRSK
Vc98miEVI3ZSS10L7V+6R6kZOyDaQLuW1y2UrA6DsYS3h6K5YxvndpGt9qKPXLo0gNjVmFcErLbL
iFDOp3v9ioH0ul53ejxv58G4f065jB80GvFP6VksV0MHPXZLpFdSDHQlh7AtG0tbF8UiKb7F8ZBm
ieu6uQKnCxZT6W8zUrcckY/+3E5CvTCaG4xjg9XmupL769jOjVlPQrvogSkHNIesq/37jMmhiEP0
/JHKQThi6gLObEmKFFmCFuNWbSwkUap4vMtgZq6iEydyJ0Ad8/dRRyjCxAQPGepfGnmMSBnQHZOc
WosALNPam0BDB0e2+9kICnm/13abO/z1v3VFDvb3hynoyprF5reYIfYR92ZXIP8+ZR3z7yMsL4qn
L/p+VE+KyTPGSa36wh1aScgJ82OIVzFAQBclv+/7cmB93yYuju6VA3XTnCeXAfmo1pXqcDZm8U6S
w+7/sZRxeNVLT03EhlLFWTbf0vB3Scmiw9mPczdzGprQ/W0599/OTyK832UcKLp45/dwFx6hgXKq
gx562vm2Cc4M8x2I5Ot8Zo0Zgu9PiFroASh5yd19+yLi1cZNm1QJJPmPajkbut8dLBgvY80Y6DZv
jA0yOZqAiunYrwszAf16Zni4HVEfVUxL4l2rbx+nglL3Tkk9Dw45XhY/DTsOUi+tPomrLJcjdDU8
ZryoA0nkS/B/pWIp7n70aXxQsXgthomVkjvKguksmJyTDLSunZiWBRFg+/m0rz5xlmQ9PiGJeAUu
wGATiuSr83qEO9GkoDdMADNSMH/UIg5BeChe4lO2gEPqNqvM1KTo/Zux9c1zfHr1JpYaWdvYgtD5
v4p1e0Hy0UPcLzfjlzqVVcLCphKkFUjHIehsxA2VcPF/aM7LS0jqkcsghBehE73ktB1HY6Dv1Ovo
ICc3MmTkseWS9KwG0TWJejECWAKDbZ/RDYirqfJh/mLXe5xYdsOR0Qw224a5eB/Acf7lkpQfSiwt
XJNwBpVGRJBB1DQNNZN3AcFMLREv9piMepT8xiBtImJK+rpqdA7N8rIsbAlU7coQ2J5+cWE6h5+X
+rbKDlBxNUdzJMJ3bhmvHmvcoI9hJTwaYEsarJywTk3z7wQRR556X+W/eZ7AVjd3qy+skrFxuUUH
FdhRNV/d8D25BAo/teDLahq2rGP81CYLXV2GfkFrhgEUlLUO0smjNhnJ79Gh/aeOujis4aKBPl0X
/RFxCQ+nT3xi3VSh5qQMmCKygnfI443sfeklrKskb4pgBuSSHZKnCsQfpiW6sx6HZlmGbaa/Jflj
lDa2S4WvmOuddtD+dHXqa5vCPmqgtCYGH97WctxyvOGB2cVIuiiZFQE51XynpG/OJNW7W17U7/xE
moXd8PXngfP2+G+0ROXHDht6svoxOgqMzEn00DhPyDt2H1QOoP4H96KL8gt/shmhCo/LlyKlC31t
cfCY1AHTHG9kDf4+XSKDMRA0L2mU0bFJ7xLtNCDhw5e/QrtF2gghnrKwKuDGV0dc//823037kBgx
dGuJIvCUEBv1CCrq6JEDhAY1e3QnkP7TkbsJwykBTb7MWwx+GAhhRB0DD+B/tAh9GDAdSFW0+h4Y
dR7AIG5PjjQl3uaOTJcxQf3e3SGSb5qBIZZ7OWBsDh5zgwMSWgaGlEcZDEvRHeKAUuZ44HeoGETa
q68zuVR5hcKbkr2Z8uMvxiZd/R1hODSePANaciPDtJKu3LEYkXsAB18hV3i8whZWeoAIWoFeGFFK
VNUBEd5ctkelbEa0+Fj0IEpPXJ/FgWQA82XtEDijiyHtJhqBOJi72sY5fUjL8LPJg2Tujh5NWZSE
FUXLcua9lrza6rCEO2mkRv5+IGJ/bl2nTuJtuspfOiPF3ffca07Z3XLflqnwWwHfyP6HbdcA9oWa
wFLo6oAdGtkwz9jAcUCYChL4iFjkhEt5Yy5bGTEZGxy3mW6LD7hV3F81AbN1StXtqkdvBY5UBkR4
hdBAeT5U3KbbFBRuzHkq7eVQ/Wk3kdGsvwotZA9kvCjBcpZ6Q4dihILnfe8G3nlLF6+9b5bQuO//
qHkYoSDOOPdEHUcPKnqbB0yKWp9plyDZk+eK8NZM3w5NsD521cYPEIrKwjKSbB8ynNMl73sn/ZIO
2bM6UnFvafo95/IH6UMm6RKNrAqisjZCrp1jQd3zgKdCdldVFpMFqWMAfx/kCLSI6OGab4H49G3m
9jfhaYMA9YUnZQVPB5uh/CscYbIA7efpfEGgeTBXbNdcdUcirsvlYYmQ5MtawDJSHjY5x+RAjrl9
g/ydfw5KZN2CVVQOiYfeE4uhaLm/a0jihO4ySZCnP9x4cL1e4ySDS8GevEnGxnI5UqPYYmn5vu2N
RytsXIJklAj1vGz1jQvxg2hYHymfwWph7tsBb2bRD3exy48zUspq9Ae0DgmRD2Urq0IN9mWCsmhZ
5YMMChUBxT5xExSRJ1WsyCWP6BPCZyuhntqdOD5bYXbvfuhjF4ddq9+HnI11CNGyvuI8rF+fI0J+
+fvEdj1xca+nggJa+MNvupX0Um72sweIVt3B1eT6WGJz0a/W6zuB5oKo1hjeYjeGnIIL+XdfQumA
FbZnZbn8lLhultND1o2muWE9C5qFm4LXFTo6m08dVCWueMJ6AOMH5Rn7wakoIA56TbHwJpGcT4Vz
kwUeintlSe1v4Wh+SHJqu8pwVbM/s+1vhThD09JlhjkNZxgoIn/mVfJlSHbEtHgeULVy2quGwsm6
xhT2q9fNu6DNxC9DmgpHR/J3mxyd8C6R3vXLOuSYx6qdy+WRiXEtPSjxJcR1CQYIxfAwJoWtdemh
68bflLOOVZZyD6JF7EY9J/0FjGCzgWxwKWW9PR/+m2Uy1JjRDxNdboHAnu2rSNGJH7kg66NzLB9Y
EREOfzMOaIzmdYCAtwLcXz5O/1amu0FkGN3sUes9zMM4p9HsCqUUp1rNciJQzOh5p23kWz7TN3qo
U75niWW2msna4cM/qiT8M45Qd/5bfgWuyd4E7GkbvKXcmq3+uWLV3MGvJhAAidtG6uXi/U7Cl15R
GBxLBFN+sf7ALOu4b/B3CyRNFiwGwJVeRcjLftj0zhQc84J43KypOAsnyGbKhSYf1GpQFQLbNS/x
/kZuKOglv8lWspJvWzKgpnLfi14YgtQPYzGVQwWk0a1wgrsw9Ni0BSDBkkNdKvwoSN/GSoswDNsw
8BiSIjmp9QYFsC3FyJomLlH6TbQ6BaPPnftXd32ptd3j5FqW6ooF4YI2YJNmnzzYue5rXpYi0QIS
4NIo+9lrLnRoeuamPJIqpj0cxXhiqQOoPiGIzGG+g8ZXybsawYU4+9EbXuTM76BGjWcEP2noC82V
/Djn9a60uZW0AYujZQfhxT+oL3gIw6tTwqxCGLvKJYnt7/JzPMhgk5+/n0DpVtV9jWU7O212ugrE
vufiYT00fJwf2YSNsg2JotQfKe5TosuQ0qdrvXoljaWqNRcV3nPW8pdkAXRZLDQRBHIkOsA2E7cB
SiXvmeROABCB63QoAcx2BKtmavNQEQpB7r7nBIyXD+2s5JKQYcI3KwpmbQxdDP3ek2CJ24Opux8a
cXc4cnqB3t5DGNj9xsBPmnMnVr33vq9GN8vkEcMP5ni4eyI8Hn5E5odFOYPqdhstYcoZgDDlIP4/
mnU3x9FTxfv6Y/OiMVygIqD2Rqc2juLWdEVADeBIelNijBJNaoi1YvWaEbbypL//7Kl1Cc4cDffv
RvyviOLaHR45j3Ra1WjYtvFPl+QeJwNWcOLpecQYEVntV2tdvRt/oY2RfY52A/90mE3BlaO9EQfL
zD4bIkTTkAX/2pwpdPkBUv9TCy/WKi7tiBiY73ZysIgxghiBKaqUsorVrHY/KGqXkVcgDmDaKBMj
eS5Flaod0RW3s/Lw0NEp/XS7OvJz0NcF0hfTj7nB1QEYlrN7TXtLdJPon8Tbju0MIkmHfQgCya4p
Da8ZPMTntd3/9IiwKxyscEPI7JnTHdpWfhG5ZdRt1CDDtXLcChD4XpT7lVhiQDrds6xFcw968Hv/
Cx+Z5y7jreQuLq0t76MCPk9JadUM0ANa1nIKd9jT9ovEVM0EhxDv0YHFlN197o6HMLedKH/U7HYS
ZeJBt2cZNvhey6ksDoJkCIpstxUI/xb1MdWRuhrngmszUSdu5xKQ6/Zh7RUzm5dV2pphnzWwrS3l
zJkz2SUGp3BEwzyLaAXVzux/l7hc9qIAb+xYEmwzc7SFL4B0buu6ZtuxDX9uzG79RGakxk6N9hC8
NdU4WB4jHYjm2G/0G1pZGFwaxWv+cwJFJRoteK2whjG8M/gqmay07a5htywMiBncC7TkxTytoy7X
7TyRmjKoUcTzYWUVlRZpKXEd9mdjx9JTbf2dHmU6M96Q/lLSXZJVabOwYx2dnszVDc9QY5RbD37S
tHEYg1wVIuMksDXBly8/a0Td897dnT8QRt2OiTqq6Gzy9idPW51koQQeb4TvH5zYdjx0fawcBLVS
WbNh4kbbbixs/Cun9QadESourCGF1lHEzjMS617j00fqb/Gimgolq06up95inekkdIavrE6H74gA
9ASL+AyDIO1Uusv63xjjQl43dqEDxCT2ALQceRUOFuYvb5vSAZK0Zi6EcC/601V2WRX6BdQpAU5i
3oG0XgQ3giaaQ433NcKqIy2/+9F7xByypZ8hXQWZUMllaywocy0f4TfRTGXUGEUEk0jHFvFAV/OI
4caM+9+hRRKqoTnoe7uoMnnyP3YAwRt/0rCdk4hAhrdpBkFXbPcYoEdQjRI0Qha5ljd/wuQ8qrvr
N+so35lwYa5qQ8iuc3Ur44G9vWP/qSzaIPhvIGvivIsWJec+W2r6Ny/s2LhjP7lPvEEMiApRMk7c
cDaYOyM5VA+mldLJbtqcnf+uMobIM+14+2wh7UZKYqyFKibRZi9c6weBseNooQ8yBKmJdUCzK9F8
q/4v68Uee6v+rDo9SN5uomebRVFYVTtF4ZGq85Mn4fBQ4zo04Cv2Yy+A5yrz4izh0rO+v9wfVkyg
1HVvWwZ2gS6wJNC+KC1WPzYRkkba7CaVeaEh2eh6xXpTRYAG+QqST5posgVR8RMw6Hgz19BLXULM
6EA03zR7qo4yzTGJKmsl3C6H+SlG/bdvEk6NJ8KN+kYb9WywLQeoJf/266Zse4CWJ8jmblOJKZLX
66BcIIyQ1jgFbSg/9htnTHuiEhYCU/+yRQpJuvH/BaceOclOOVthgtPsVAUe0c2VFRZJ46u0URMC
rGJdlbA2rdO4qe+Crqt6okAWpKuxrueNzNEp87sLoK3Cdw/OGDB1ZVXNsYXMmVY1yQyiEJczeLGS
Zqg1Silx3oRTHzTfaX5WC/65Co4nhqWVgvWQW2dI1gc9Z34z399+5sbrixkEb1SvzZ0OS4Fz66SU
CqGl2KnBx0apMuOD5+vjETP8rBqsuzIcShBuTT+iqOxtWi9mATJe1fXQOgufKyhuj/h1TFB6wGxB
fwAJ89KQMFtd372lR4E4CYGnfrW1xxDqUmJm3zNOnyeQAZsBKHCYu5oNcY74ftbkCGNbWwBX7rqQ
PZpsEEx88lnj7TXeO2/0N8E/qLOW3zIEZenpAKdBruHamUJrGz+3GQY7396pqWtVP3EoiIEXTFxF
l+OTE7P8nYarwOwAkTFX28+jToX+vhEoRUaW15KJ9orvuQZXPoxRBDZBbXWhHbkt+uX5rFY8Q/bB
hotSZwKDP9sb0FGAWLGaFiOj68PTavfsFSGxP/wpS78dx1ItYTDcBf04ZCSogGtC1h/8Hvt4Qbba
PwV0AbQVm0XoZfTvOgSGuzMBkIzsa15r8JKxNN27RwbWikC1ZDYru+DorCtnFBBiCVUWz0ESrGCm
0TkcBvLc3cOLM4Sqrv/qHg3K0J0ode2uH8HeoB9OokgHB6Y63eEEAjFGrURnyqUeWMZo2MQ15PVM
5Sar57xRWvp+qw2E+oEHkAcWsWovd/qLd3VbG8GOPAkuz14g6BrAugeTXqRHfBuBu0GE99abgeu7
OzYVU2KUd52cBHM+nmiXeeIjTYyWfPREoDHwY5vk4XEWXahPAjdX5fUWWxvEKjVdbxVJrL8XLzzM
1FRGaRF03eqPB8xvqtoDjnPD4ZqZIj7wb8N4hT1BrfzOHpovdSnMWvwMqzjTBYArqvONYc8OC+OC
9XUwsU7stMc4H5B6MWaW5SThTbDxXgI+rOrRdtOlbv+1Bq8PcR/mkTJQKOpSUDUJj7QCR7h/nnYd
dbu/Q94waYVquVzX7KBGKmAgMbnmy2eEbkxJmJTPCk7AJTXGHBtVgnbPyWH/bB+kHqWYvpcoIqFS
DSD93wAyIgfTvpujAmMryzzotWS1mrNvGQoeQJ84HEeBO8BmaqEJ0CPIHJN+sSB18xuanLNFaBQO
DCwTMui7YOmhDg32PJBoFZKGK//uITPsRdp8yrCT0CXyFhc7YOToOf1dajMt1U47Q/hU8x9Ucru4
O0MPhXkOxgmyRtDLWL6qinv0JGRDlOwxMk0qcnKTPlch1CDIzZF4rq8EGAwppcxGudUZaNcojCV0
b6hFPtvsrxC3FueyGR9HybcyYgAOqbNm2zcF10KVWGemeRL0vdcXVWeGBjLIdty6z1NgooGckek6
XOLqs9OQBWLq1ws1rFxQghbdx+u9QuSqP9ih/7driABOVqDtGqunT3aAtNvEnGG1ENptAWJ+fBsq
7SKBX04xJqYV09JselXMHQypIWRInLBTTO6dfX2fk0iAH8HDRjQfirn/VOa1zUcW+bVEhnNyz1MV
XETxwGlJnGzZzs6UKVLSCCAGwbYocr8gGvPXNBB6AR2xa9EvxjzDuWq7lYpnQHL3E6k4ndquI0ER
HxL7PWN4oj47G58QvAF7Xg/ObicraCRYSK8GhPrtc+NwveltIufWs2z0/e3XylKudqKWUnDvVHpi
jIDFBty2zx+Z/6iA2AQb9p7F2NuD0HTaLmo3MhowTwxUNz7WbhzcFtmUFM+lvKYeZtnp7sl371EO
3MEE+ZeK/qZw/SgFxC+4IujrWzc9n6IGAsS7n5vc/XhdhI6ncEVHUCwaNRcaVFMvXBVTdnmuhsay
5TToDH9ZSEFbWAsM2VE9arBj7nkLrs4XbKvKvUXD6xHsj38truwki5vG/gNRbyd7pS7xnpwrd8Ly
Fxip47oBLiFxa3uN+mjHddoa1n6pj6F+j/xfEAk0OAm+gmLpDaCa8M46XUUXYFVPqIrOLlD68ET3
LHKxhRI8E16Nr3TLwUjyW0I/SMybKvCrid3sGQIoIxXO+fTDHhCq3ZfwBBTr3mEBfuQd5FpTxe3S
e8EvuTylZ1mdNlTcZZVda9vjFR2BB/iS8qLuEBKNfr33H6EXubfRx+WuOe5klrV/LmWKyVh/epKD
LMOW4gj8Mfp5J7MrOhhjKGyFsdMm9FMQTfpSA1v6s2ZQOUAC0NkQYTJcR0vOr8cJsh8GUx/9+ITw
9m/zXuAvHVd1XNZOM1Od/F/2OUoZviytKty0mGgeftiyclnnc54CdOSFszwgUo7BB4oKOt9T/fgC
5aB3jZmSArmCicCVtb0m90s0I6bYn+I6jLaA98zQhU+EAkHjz7ApzuOqqUNVO+Oj3g36MCqjCFQK
75fPm+j/eSZyc7CZ4lP22igbTCg9kl4rEwSqDpqJEyjUao1k6pg9UdcTY4kdBPmEHTII9/LHobhV
g/yXoLpC6e1rTazAaZNmouxrn0cmExMyTH7fKX5hfDjncYoFmzGf3Gy2qOKuvaPJZAhZNdCmWX1j
YNNR9D8vD4S2bP/2YtbhhF78aRF9VAMP76qx4YqdW+0Uw2Bzaiw+b1CxhDHbgLNmhRYCmt/EGC3d
+cM4ch2gscmfMdiTSTx9MpCrgg5MBODZtKD8EwTypDQKbnN6J356CerD7h5e3wYhwQHgEh6ydZ2U
pM6QyfnOrJKA4FDA6BKDnZLd8VoCfl5uecEV1/4AE4s9mruxBbBbyOlqaV9ZdJSt0qmAK4ccay8S
M7dtdcQLy54k5Vyr3uCnCRmPqZaEvAk06CuvLwQcDfh6Hs5siDQnSFtnW5wIWuEQQwpkp0TnHjR0
hd9kDTWYK8QlLny0U3tnQxoMLXWh/KDKcET1GmF7v4DF8LcGR1bWxsyyX/aVMMbBXdKzPs+8eBsE
0M5QzUWvEYOswTXHQuv/DI2dTE4WoljCq3/KC16I2NLmhyLCOndfr/B5jWnt+G8DXGJi/7igPUm4
HMt3V2CTxsWQuvlzoAOdLH4F1v+bKZEkaHszS8nCzf266kpCJP4he1J1sdheNn6gfotu1O9aPZX5
DD1TlG/ZhrXecFjVHE7IjPVH7SueD/7ERhHWtVpi73cHXUUc/6YW6tep6hFY0a16sN7976hutoa2
ziMu4qMNp6FA3MrX8UMe5pHVEwe6J7u3dMQ9WlZjpXzYuSuiGaUIPDsfDoMx6TZ08hWTEe0PBZFc
/4TvYPcHwoyzGLYNCOHcIogrZMSR+z5lDHI/xc9YKyMbhksJDFiaJ9OuFJqWr9oF8aeQYopA+3qz
7Muzb0MGBgmVzPy7vtdMqrff2UORvgs+3Hpj31yOKjJ59fn1SCemWwcj3peZ2oEaxTOrYlBfF0Z3
FuDGxhVn+7ANRrZPw7kYaY8Ox0Lk8gYwj2+5PKINZhvXSLxPKPdcV2rqCWgMOCGhSn63k+LDtN2Y
4ZyKVaqRDyejsi+rOJfuvQ7Kui4YV5Mz3rYdIfZrTNE2kgMCftoSl57CC++3ibjGvDWcqKfY+kZ2
mFqFGAYv9aeFUCbxeXrZ6cglQ1yzzCBvr9P1uqGGlA4oVAWbJ3DWnv8wbsEdE/91FkumgxLJFTIP
8nfEY5LkxoquW0TzCb9NpUmhDwWMTgTp5iihlbQlI8bUnibVkZqThBSGWIIcc6IepyDHqBkyyQk3
1UM2K0XuWEsZtpXaHBAUN+QhZlMGWVEh+RQvAtHarJjjmayjFwynLxH0Zatu3ubc69mBOHEFaKQv
S4foyti6gXbkye/cXPVIfsw9D5Gp9jeDquzbO3im8jOgRC7HjRIdlik4qyel8PQNC4tjK954yAND
oRsLrZXGPyTGpCpNwC2XHHLdKcTKzzbzLDStJ5PwVePGi/wDEDuqzAnRg7fkx9+41pt18m1cO7Cr
Djqgn22JZxwLDDYGLEwaTkktAZgOhPJ1L+nuAK4XuelEZPZlUtep7J+/ETRjIRTLRBCQAi5oVeOR
eCfOspteZDZRNHAE91Kre7kfZlwpJ+Q6f+3NAcU9aztfZG3AkAX+Dy1X+bwI8OTuKMoOc5sZLsbc
/fWcLo4Qw1HGXDW8B05QF+JyY54O7kRv7MIYMqkCiEdK8s4GKN7Ip4DD4DNihZByJbm2cHrDvDK+
SNucWg2jL32UPWe+CuWSfYa93cvpD7wawYiGJLozMyuiCnT5JcBjq6aRROz1SPUIQk7FZfWRxmWC
lGrWYn8HOErjsNskMuoEwgTX0D5dZeU/zjHjtvxDFLYdUI2GNV2iIlkf9e7DOuFs4eHHJtg047TR
2+TckIqruizQmaNQsDZ2edk5cRNKGZbQvgKDUcv9o58ysSiqQRnJOhAta/rsHqUEF8tBeCnbHf6S
x67T3+SZ3ZlXwrAD8V/yrHg0FhX//vqabXI5vlMOojlsAdv3Y+1Z+GpdSUrQptvI7kUxms/pgNmx
niKiRhNAt23JHeqIFvhAGf3PjESYElKdYDvU1lYQPMNqOu9zk/Uzpn7n7XZl/xe2MRIzpuxFrafC
9yxDrOok+Kz/JkrOIOarOQMIRuTN2vhxe62qiCkeNztO+/CHbI+8tcbxVdQTtBWqtTgFNMrSdfN+
F4b7N2jgK/Lq1myG1fvtOv2qg9sQCgbpRMSi+KCL3ZP7+Yg8mmtKVEnwVTDzgyeAj2vXioAtb02m
HMvDr5YE58duwbTh4MvhWJ1mimyepn7i5TJC7Elba0mrB/eWj9hjf8TvtuOavZKsvkO0aiisiTz+
MEhYSE5M4FdgfNpawT3nQcevVTmwd1qNSc+X87XtM+kkX5UnsjLTgVW618+ijZ7v6L5rDVRznQRH
e9Evts+YwfDpOdwAX2iFzOxNfBlBqAMINF65RG6vn7HBW/hb5beBaqeFj5fMtWDF8OT41TN6jVuW
WwUQA+6RwIlrnhdqppasSB/hz5yvY1cGRVrq/wdr97jA2WSD+tWtD5IgNq7GqwRfEzY/PqbaiGUo
MDoMWTaQlACGdvBrLpaeEoDka78r8RJ5tfxQ9ZEvHljkumWE3ozfk78i1zhdmqimGSrCpQYFSJr9
mdM755+fviyM3djFAp8bP3HtXnaBw0V72lgeuZeZEhdnP4Kd94FdTz7eWLHJMh8ktUIHttPi5Gv7
qg1fUSrWNgKEbJrURMlZlvf235lNAcgah2v/P06aJ0b2OiCwP3r1r4dzfBEKA3AMi24RMkSs/Kyt
AGGxZNQWr/ctBOmL+cmTxk8fQ6QOZno68MpmWhl4TWN0AB/BqsfVX4T3C7MboN1ArB1UeyKBP3BM
PIRDZ2/xTADx2FyHcgIucXhiqW32GR1RbSLa3TK5mSSoZPvfjhiygQ/nFMrqYyu89LfjcUGAvtLW
3k18lPZ7TdyWFf6gx2sity7EIlQDLxi3tOz6oqPWblJLxvsFf7libzJfC+boHeV0iHutZ3ho6Rv9
q7OsIiY1i45RRYtGv7rRmKq1pg+bSS5mLw8C/nmNsPUSn5/FzoxEtGJ86qmeX+0aIqFVejfS01U2
gyIwlMy1Lf7PnOFtqbcfW05CQeEIBogYe8tRiLqViiNGXNn0+oGPERSfN7WTS7RC0CoXVUCYc4aP
7nZAhOpBzjZMySFFfPk5QpZ0oDNst/hnK/YuvHG6/iIqymDepSUBa7SodN5arrwLaTBnulprSWOI
Omm42ARjXGUXs8OFiqZzPSU+FmrvEqwFW36xq2RuV5SRCcpFzGGv0HkkW9D3SSzvihN+RMEsW+IP
gXnOUbgD1VZ5egXsTLnwE26JAjGyyTR8xvrsp/TTaFfkjVJb0XRb6Zm0TaLmeZt69Pm7Ua5ERQhA
ERe+uFt71F1S1EnBLPoNI/U53E6vEPqvl0AAJj/xDlbVugAF18AVObZ0KtO7cRn4g7UgvBNhvejX
8io5z7ik23TATVqnBeHr/Pj9wUnZr+6sPOHW8eHqbD+mg4nL5eYY/CxXunmpY28/7hi35UvwrNeS
Uai6vSls4m9tPR4xxUgIYITvIx9sxJ8bnn9LTlGjrel3wWIWpaPcUFFxdJju16ymaBf3B2ekLkT9
YCk5uqYv3bSrzY7l5cY3tQ7eCEhx8t30IXjjPndNXCuYvbHNgpXlZIG/QuEtuUCgXL9o0Djm6diw
x8YDJnInP80RFp+TvKyeDNL2nyy9eHDD4R32FduqJppbXJ1ZLNJR0ippvelbfWCbwEcmP5DrAbjF
+jQBhyz0qUIF0v7o+1YLGNmoObQ45N0qjvd5d64/Tlub1rgpNDuoNOsqwJ0tUFf5g+DZzCa8XMhU
X8MZPSsdPf7KdjFWkv/7SI4r29EJPDdBG+6UfGAIEp8DYYbC9jfyFEFHUTucbnpBOspzt1XNwDUP
kUEqifRICKoCFFaLY+0QdRR1ZD+YG4b+V/wSHtxYKl2iYdfEX6uW77S1qzV/PQyY0rFAsptSkVEM
XFkhTqvzOOOYaqHnW/NGqHkYAoEvF3yPovOyg0uudN9rjFF41felHMcbywQiY7iqD4sjZQFj+UKS
XjDgCvpwHrZoKTAW/yZTvREvwPCcVFcVVqMbs08NDFgMQY/jVX70YRMWtQzPRk7LhRoTVA73GXQr
Zm9I9Cae+j82a9kGPLv2nWJ+CdNccQgIpHr1VcYBqz/sutzlq6d6CPmX7oR7QSaThGIoL1/mpks+
eU6qvdtHPx5bxXKfZ60naMNbPSjop2KAb2hKo84Mr9PDgUvr7JPRAAeiSq+7HOSb1AkJopO96EqU
wJvSBVAeKOwAffY+p6XS4pCCwaTvVt6NIHERPRwWrSxnHWqGPrge61cfTXs2G4F/uCeQuHu0Mj09
03HeR6hutTvfy0hsTEwU4RJ+SE5gFRbiqg+jggleQi2qVm5+ibn8gru8/2V9uMFp9ZzOXpDAaXGc
t5u1fnOq4krM5RXy0M/jFtKLRsU+NLC/hF4nzos2ob/KGv+c9FSETJ9fUeaujEAMds5o8KJK26KJ
Kua0zUxOSOgsplKKs8Qu6537pnDxkIcxVB+MZBUNkDcoTxRMb+Uxc6jEa6V09q5gJ69pUM17Uo0p
afXsAvVXXVmghC0iE1hpKzRJcNHjgMpFOB5ld82F9DZga+kIGemVD/IJUsKbc2F6dtf0oQy4VAHF
4nhyznZQh/Vp/Bv/JUqIBX5msWfb+ONGVhssZ6o9SkxNxu09vyIL7PNtAl7qzoxtxcCVbnVLSZwu
WRPg/FdzPOFoVe94QyrfUA6g2TBPL7B++KPxl13xioKM4dGT7ytHGFlXLW0nySsCEAhpVzO8Xmxp
Q3wFXmUJoSbTZUB7j4W34VMROSt0s0TOj1LI1zo/Jdg3DcNzLheu3/ECVoF7slP7SRgo58+5FW6O
BdDznaTT1wBvRyyMXLheyWDZLs6bHZBagbe/et8ajE+JqBdOU42j5Rlah1X501BagJxutFYZEQL4
UmqmyTKCYSi93AUu7NEKiSxAFT2GBvyTSQ01NRqGzCHBhaROQccKOnCf70AVg7Tn367i8bfxUFLE
S17rJ6hqE0vEAvIq8asfLB6sDVwhn41vaUw/CqAtep2NdU8pn4mpMcB+cQxtoftejbj3/m/vN2CJ
1AMVSzAGLLFY3KkS77AZCfK2sSdWPYzLP8UACPsI+4EOUNQoGxhFHrO2ypQ5VSPs7OvmRpWz1XQl
DYhR2ujy1jy75FNXvCxhiotJR1Ep+Rj7hei2mam8H094+pPQgSFqDI1ywuJwA6zi5n6zPRLUhpvS
huG7dTGS3pr/dWlPgfQ9v17m2mm2JIYqvvrk91Ft3zV+lm8nMCOo/izJhbhGTMJXPFx4dGkpZF2g
sXh6Ifqwz8bSKSYR8C7SCE3lam72ED18kxdgS8QMhzWZ03dYnzmTixNU6TiwLx8f+dT1SZVsYE35
UWGkYFMaXdKZi4dlpaw6Vv152jx/XnxOZ35F6Lu0A7ZU0dgPwblCBXm5c5ndegz/5+lpdZz0Kg9U
PcQ2TkNYXAP90Xuk8HRFgup2gfzfpRkGsWMWm7AiGO4P+/0TkPWb3FEI6+pZF19DN3Jq/RLHyUM/
F4kW3DIcD/aHNXj6tmTkyLguAnDJUX+5xFItsFuEvoMF2x7OQuNFbFJI1NWWSb+2cdRy0hQcjmeT
Uyx+E4au0zRUd/YqDYuOO3Qocs91913chGT0+U6XCTW3p6Wg5bhm0Rxh9BoLCBMp0rMsVVxHLJ9j
BCi+YTVKNZ5lUlR0+/dYUQ+2rfnF3r7hxcsDe50YtqZQMLt+2Dt5a7UZNJSreGQCPjyzdFrMaevG
dr5ie8OYlxSZa+NJiW5qn//JIJNE+/+7le28V7J094P/RD7a7nFc5m8M2td2edG/Fx84lmgPdM0m
YM4md/cdH5yUaq43Gb9C0WwsPZNbQhVEhy+xxf/5aMRLcTmK60UsYtbAfIhZDdcljnAuU+5Mrszi
uQgRT/A7PDsmcuMddJUZFwwZYIOWXlno7k6epqXS6JOmSVPjD1Dgh9d+adOJKM2/pkkUZ+a9+DAZ
f7itNTb0FgH3n+2aC4R4dffUMAy10lGElIQIQWjlsTnXIIVjZQhTG+TvId0QYj59gA/oM5TxjZgs
gBzqmyBXp28ManWCKIYt25xU2KcUWrJ6UcdWjEItM9m6SQ9Hq+jzldR/nlPJ8cE2G3xyCOboBnpp
ZkvW7FJHOtPKSQEkMEfqrpExjqJG62UHtEnzoeF214+kQ9wXQSyM4MsqrrTEOFheCNMga8uFjTSy
ICagh7dDTguV9PMVbkMmZXIEHKZNjNleSeCxZcsbapjr5iDocCdUj6PVhCTb9icBQKQ68YNOBvhN
zEiHS691aZ/yFGy1gddWXREPflbxeLBf7bU8iJDAoIP+kGsLnvNyMngLoMVs3er0oFlKAxzCTaPd
e4AInPUsCnwlFJPiIAGrFM/8mjHYxTmW0Xa7ZvXbPVgCiRX+tlSuOME9bBpjuPFcxRs77lJKyChu
EtllQRxY+olgSsaUhkAQgAwyWApPwlZJ1EOWFA5GMRQmBEdSC3rND4Ngp/JBiPELcwBmva9Tdtnw
iIt6LfVNN2QEDDzxayliDCQaPoHgJ6GIFuwW38qp+hCpAWBdI1NgJ8bWHVOd4YETqAhSzp4GxM5X
kjaCsHYn5V7H8ZFt6Uyv9x6yW8OLaxQzgw8Mt9aBc5R3uZxAT7i03OOIn9XMgYCgBAx6sOQnoqkQ
dien5WAYTQlhSH4WeWFk7KxKiXTRUW5GWv9wRQGnOBFCJ/TwaAV4z0g7jMLncRQyF3MIsfgW4QFs
joSZitIERWtjy3Oce0IqKERgS5sb5SdAoloZSz7KCtB3ciplJKqk/+2QM7jNUbUCI2hsUCx8VJ4O
2F2LK974IENAV9Y7dptEyuRkUAlhj4rM1zZ55I3CW47OmwMEzXPrzLlrZgbS8BMkyS9KBf3wyTxq
HxRGxAclDcHVarfDDXi/oYFxM7WcGJX0ba5/Z1iOYlCtN+XxyD54S5VDjgY2eX6vUMe0v51e4neh
O7IupUy+5nxBvhZ57J2BtEIiygnQU2gRjyAfouSWkikgMleQ6mQguh91dyRLDvwybw4eZNk4hOrZ
KwF/8jxXg5U+oPlJ2u/gnXQwxU1z8+jXsnVoHo6/qUaeaNrJ7cezCIlbdoIZULM1RM378z6zlWz+
fYzsBsDnx4PmrTfOORDU1cyhch5nQyVcuj0z1c/yl061vREyJjOhGsNVmMErYEw0PSIwhyyopd6U
SL6XtIA2rno11ZF0oYqA+15QGUkcp7O46CgOQqGo8qsClhYVKYjpcSR2ZvES0cTfhu9ZB8yG93o3
rcKTXTv5AI7eEBJnzeq2GFVeLZ6LI5F3/bxZGr7+dPXiwN5P2n/mWKIaQm00wmNnIlVdSSDCXI66
P3jpxvOj5+P6cU7dZrQISM74G5WjghjQkezJFNLsLGU8WFcOePepUEkuzdxjaPeAG5YOlymqno53
bYLbdx63TQY4/UqOvorsfxHv2fb+06p5hCXficjruz9HDwJwveJ0OQt1T5m0UgpYx9+ymK0sJVGN
VzZy5un2h22WF98hlOn0Vd9ARGuHJe/WDyTBkgwXwP6aa1s7poSqOW9pwR0/w1RQ6T0CAp/ZIcGR
ZjQiUbQLvoKIMsJ8Mnnsst4BlohWjyvlBNH/cB6ckNaOywF09PbhOIbhcVgKzNwasUyabmjK+0iQ
K/t1SPgcmtH7VNl8eddJKawITUKPsH8cmuaS4dWMxhJlXqKJR9TYCngBJvGr71j8myLDRTq7YZOW
eC2nvIIs8wgTjGV/aLYsYgXBHP9gYpJm1d3LMFiasEfKCLIpVD2lIAxRMkOcVvtAj6T3d6fBJJta
xmQUkR1mcP1+dqF/XkNVcLcCCboo3BE3xX9OGqMDce373AONLL6MThZ3DmWStMuS91oGokItALab
Ly0nz4JnpDISmby6zEZnD723sVnM8Rf10CYq+yY6t7DxK3mixwF2IxsNgPVUmkNmay+E0LMyHtMO
lEzch7JjN8hwDpkjNe6/EPWzQ4v96eO8IYx972fcD7Q+16TuVOiZ31EpSMkL+XJf3D2fYxiWQ6XZ
LlvvR/G+O7o6jsz7cWcV66NbVwdXOb3w4HT7rnUCVZWwz1/ZHbhJ3OvF1d2lksC9SdY/ERTyomCp
dvi4VVuWwD6zWB7JEkBAxOr+RX40dp5TlizLrkMCBsht8voNYBeEjNEO/yYaV81OrpL+c2o8jzpP
3IjgZ8DXUQDAsPMujwwulJLb+cn2jF/gtdzN6zWBvh7rLwrjgvVEVbWuliFDeT/IGQ124jBfkVeb
+1xEBpPNHBQCEKnPEURlGPkFfVom3JJxlkxjRY5FrxM80bHsnvZNAn6lFBLY2yj2OfyjnaGNNjz2
arYrFQ1RuBJ7T1uCzzerwnxpOPSQkK/l6Zkg8x49kBSMPOaKE3S9L9EJ0Fgf17vGkJfSo6rt89V5
mwMq09uNTcNKs/PQY3Vp6Ph1mIhJPRVSvedEiiOJnZWO5C2BcjavWvCYVN4oELjv3zC3PN8UOlIm
sw7+V3qcjjCbBPhQdgFKfba1DBHtj5mXZyg8WYmAMT77AeBpekrk0DDSqm1J6FeOwFSKc92plpEj
y8RiMfHi1ldaW0J4eyJVvbWCrhD0OLyvHBGxcqGTLhjEDFmAxz+txdbwLFFaEi3jwHZz+W6XOn2s
nMCVC+bK4ogs+lLmfYzVsVT/7UCqTI30nNur+MQWr2fvE45mrDHd4f+2PRvWOpM7U3jE9+jJwx6n
++mf5aumpmZzPZuVpKdWoSz9ePAgmXHqErcVxLB1j/PrDqkAFzFp2af8oJSBXRuvyGCam4JubmYD
kjKiegjUdGLCh25HjtDtQVxe1ewqX1oRr2zqSyS3X0dGU5U82TZF+Qsezx+3bYQxjMw9We2Eg4Ql
wt6tnpmGgUHiKyawGUym1BlGaqPXy/YW6+ZXvtfaktu6DMyAZorvO38ARZGLCAxD8oerYZ6Zf4Y9
VPA1gvaAveWjFKXPRugFeaL6iUN3bWr7vFicBnCq+iAc2zFCl34UY+hW26P+0xLDxJW4346oBWxd
rYhoDsspzGGIb1Cl+sfS2+Dqx4fDeUrX9o9d5AylNOxcM/ZCYCXzSJI8Dbp7DVmYXbovi4FUVF/G
ul5AGpFr/gOXQtmaxmHV33hMKHzBSv/LflzkUDXD1ft+3XmSRF7/o3R173gjKkum3Um1b3c3uUjz
Iq9mTO0NndhyiKfhFXoBJklnzH8zJWJnZES/twZ5tdI+gWNnHgsLsX/n9stVLNi0dLYt0X0AoyRS
vOjyG8KjCZvvdFJE+G8pR/4IP1wjMb/XMQgNt2bkpzxT++M0B0mcGOYOcHn0GcERD3N7mqFL64FO
f77b45X0mZwA68Lg495k9wiAcZYk52VoFkC2zoBid1FO/UddSJf/bz+DBye071NcMwoSIQx/YNp6
1V+j2MYJZjEWLSlq5X7Jq5JERW1UHOnXJncNw8Iv0UxXYI/Y5QoyGMMS4miMKihIIfJqDwLjU+ZQ
jkyTrHUIZX/f36c46NrOLuK8qzIVeRaGyJGgO0Up7XtRFouzjKLtSsKSMDzyPtxXu2k5QCAzusj6
q9fsMJhZwiVBtk0woWoaANzcSrhNmoG639p1GaCH4YDwsVHzMd5q3Md4hRsjjWRz8eEk5fASsMSE
xO3bMDWLu/DmMCDThvxqoh7aaPk22x2vJGzxLx8lzdsXU01hRnM9FjdOC3zrXRq7K67QeYHoDlRs
81P3DsvFC82edWYKXXVLaasnUdtTBQn+hWc0obSRGcBeC2TOVbEda8bHcBfyuxbTe+kfWwLG/DIo
a3LmgKkLBW6xk7KvOUvipIJQnZ2pmiHFFVlZJ2zLRFP6XtTe+4LYHLtwnKwH6+bBPELB4uioLScC
4PRDtvdmwO1giLHYT+1JS9fKAwM34FZznFOKr2zxEHiDrptoddzz4PcpX78zM7V7udVUjLoEWSnf
9bgClBBEoeHFrhI29uO6KkmNMpYQOraW5USBjD1jAe47PfV2/o6SozTIPw3Cfey/eV/KZ6d3pOze
LT3NkUcQtkAiVTO/IEog/BXLLlNVlcUN52iOGA0mZKb3/VwTD7YrNLilIApJTZeHjeatRrIPyM5u
BY+MJLAItD+u+BXryokxVr6Nw/X5wDl3ou+ebJbkqSIN0nib+CkKe3jpcqDfBa6Oy4TKGoySpA0e
xg7tiOoWCqSTk0SZC/zi5Y/T+t/X5DGlsAJjNaE8SL3DA2VzrU5KFmNHBmkcsrM24j1Varcsy6eJ
wXS9VKuhiHdbhvsASL6Db8639qHVil6ROpwEbokZP8oILh6dwj5riE2HYv+y45RYUdstZMSnxi4E
nq6KQJufqYuWkVFp4BwPn68E4O9NVWFAmk3EJeyMxMKl/4bu0IhLo256xwraOhzSET7jot4jDbUM
4joJlbTzkIYGdCWT0/R1vSGaUkBORakTwx3p89qy4PDMxLotKkgnfNwMRYJwFWxC2YrTxA8X0QWx
lVEGtgrJHWy9NJVG8GO/xuprqWVVDbGXkbUqP9RXB3bk74hoeg+mSIB7ZY2kZgxNsRvAD68c9PaE
BoNZ0dyHfyX84gsIRHSKMfiGSlEY2XXE7G2YdEGjRjNcyNNLlz55+HG/GXSXZtPYnZ0rcEPW9yNE
eRqxDAJOkcdJ4oPHxzecdSE3wvR6YfCvMTfnYpRdDN+1KL+s54cc8dSm13yRUjAb/LgWzjupLnMc
yQzEiqz0pHmZa/4YL+eHzoz0ajSCkU5B1wCQhdvntvl55+5m0J9XHU6bghsP4CwaerF72Q3I+a0C
kGVd9XK7lDrcgXBThrz8+KBcsP/elEXdEUYXZOD4W2FtXIIDyz6odFIaFL/TFhhiDrfc1IFDKMF+
zNSSr6PnNPgVpDcgtNuXDILCyPRZa7wx6v+oT5p6RmeRqjhLKZI+xJatA2uwQV9nJOop2V2m2D40
1a/V/3tbC6BfBSln77x7G73ruyvq/tI68U1kyJfnxEd1frsoCcbEJ41gAr4X3AMedMa7fpPCBWW9
6lD/FOD3quhdm0FVFE0hQ+70L7DXQLNNd/B4NyM4Ai9wrD7CCen3uO4m+1mxyDUbWJ1W2aQFxysF
ABXJWC/FiTlK13jNoRsz0QyL3m0dU8k0XfPumylO4EOfkqjaVSPeSf4Tkge//MIx5K4z+qsOEKUd
TJyTN8uQwo9U4MQoG+cCSyBDyE2wlONXX+Sh+rdRm27zlJ2clEC10Ijzj2zQl51OehT6bUizjRvL
vnp0biNrKVN1GsHo9gCwNDHcUJ0GabmK4t/A3H88LllZsCeu/3se3gAEm93qcxpvlXCNzjohFoqZ
HylT05pGdtXrmo4ghMvFf9TRlDbls3lMLKMS+UYR80L44w6K9Dtmfv9aHKCC23ogGAFx2MZkhl6e
cEdfiHZA2utwTuXgJPh00snHo9AgMI28JBhZR/H9CiePUmmxC6noBj8jISjgzsFGjPpym/t4Zvge
OuLOMFVWuygur2nkLME4QqiBXzf8baeM5ziMATfv+PcW7ruCOcVBN84BiOKJX8xDdR6uZ3cn5Azo
HLAu0k4IieCk02dIAbhJfLn0vPnx5bGypc0Wa9nAgmJ2VxxJGT874Pp0QdjxuxABydXFfkeBX7iJ
HgQcgGmjs1vMdgBxpvEJspBd9pPH56DPepjs/NnVZDK0rlTiPCikEB50X8uhqgXXJ+hkADd7nfjg
WyXEJHk4XLeuH1Tvw+wtbYwWijgIExc+Bs6shxAean5tSmWObdTq0yvJvE3CmJ5HLWdjossX96MU
aJzLMi/5myLvJRLUI2b3xMUpLE5S5Ft7Tu2C0Cp7KoAhH6vDYX6eE0iqiSmDg0B1hJ4PUgHSwaNq
8PtCXb0P6hKCJ00lRULEFQF4be0Mu67OWKL2q31eQXhjwZnbP9kjIhlj4Xf1CX6J+eNj+WHto4E4
zfAhhM0CObhZ4Vyaf97HAOqr31wTdtCVHe6XzvcJxePP8i+9VxdD6KZr1k5PqADiZPYN02WpV6+H
u9FIgLeMCAwK6obAHUWKhH5R/ZYgiQMKn7VOQ4aM8Pr/ylPBbXNeEJRpRKV8xzjwV0BIeLvY2plh
WPoigvWfOD/GlIZDCkwlAP6CnsSyvaWdaNokJrA/Qy6yWIzv9sSZn1W9xcUOyqtYBwA8Oh12dVxS
egqc7fFtJXfotKJRyjdVkZRVdMNHP/YpNc2UynO6J31pVYH9arVkDBqfL1gbeWHgCvjeCcHFSlNd
LgCum+85+NCXg0X8RSIPFz9Ec+xBg6Tgu1rmNuvzWkvO/YNBHNCbiGz10y398YHxGSchROIQPH3g
rhNFQJmap9dtDCUDtEOViw7Ijn3Mo6kWgBffOtpkxX5LeBm7LF4m2s49I/wNe6pxtCfTBgfUAJec
EsbvTm7wTmJ/TrvzSfuIejDCBwSDDh95z2tQPLGzAMG9fLbeVXxNi0J7zsLk1+xgtKSYmZmiA4C6
VuXK4fM9VTGvcGEEeq030gQm5frGN7ZhSHFSLq3+iuBiIwwPhOAHvr48bggXB5cuWu+QPjW+orYR
Da65A9vtMAcoJkV1rvCsfrltxImlMehXIw2jlP4a2TYqVXwisszc6P0TtMS2RRQplRmvxLMOXvOK
QTipFOyqnqjU5fdCEk5r88CydVzzfzTRI9GHsktZZKLJCFRg+TW0olbDLlZEHD0jYSgrFFOLLnc2
9YwmUoKBLQoYtOrubGekKlWCMyU8Q9WiwHJXA2uSdYl/qAZXYR5kN98YXVZvjNlKHzeRRvUwvXvo
3saV6XWNeYXtjAPELyiTXcRRUCaA/BbzPmiAoealg13rRvDf3z0fMSeEcoa28SFfZTmOZ3txxVci
kkRL+g0ki7ZxL0GetVWJnrad8j41fycc3cu7CQTsKU6Ihag/OUir7OHpyGBYhwXcGHsXIQab2l9y
OvQtZhYcaObLGd1+k6cdGW0wb08e4ZLVfPAqlqzOyUL8s4FjTd5Mo1rL0VggENvZluBnBPFGwBa8
rzCp/Dq9khbdcTPI6VlHSGuOPrljhenVPbGdfCIDLiNwEdeItqe9zX4v9a16g7kXDbl/FwMpCXHx
l+hQNN5iaHBq6lZFrDPzSxKb3hBYwa49h+kou8CQefLaEIHGUweppERe0unuSQAefvkzjKpJmvsk
hZteZn5IAvPd9Y5XIDOOzN//Z+nOMQA4ufoAZFH5Yy8oiVoWn/j0eWr6GhADohNMJveDD5Y1bhfu
znVJOmkPue90tYsoICdxk9ndBI55GZoQYx1BIATdkKzwn84hbb0NmY4gXRcLu3wz3tUN1T0EUDe2
K0+lrzV0FZTCE1SWnaUb4uRfYuQlBeEI9jVMJA3V7Y1wS9unydcI9+zJTnVXZYY2EWWPf73IYVZM
YTjqI9A4/cU2iNXhVielXHSEMYNrh34KL2Lp63oZitKzPVQklpvj0Gjzva21NECxGQq71jpb0u0g
RPpuyevRzI2rI3z85g69UAs8RgiZrFx4obLFgfxq7AJWszKgqqlKf44HpB/ltj9Es1RNt7mcGclu
C8uncLmz57hR/dforim0nZ70qTGF8b4dgxXs+jjptKf28p0b3dM4xY4FqtxDeBhKzXjf4vO/XK9U
wxVqiapB++QqyvXC8LQuFv50khrtPPADvMDLXr7u85ijANpeeRI/+3uQ4OU+B0U6s10F2SqXAM1c
gfC8EBseytbvFQ1Nn6bsZ2W5+I2Yxkt8lt4hSio228IB5kJFXwFUra9UWnQoENWh7GxMfnX2DDUk
XMWMxlf65Lq+aqoFcXu6agHN5dKtMdFZSTbqlhxft1pQ0HJDKAwnzSEU7IZSucwfIpbtkaPZ9kMK
whkw599VmQ304emxE+d98CQGJ1wzJl1kOROy4iY9HAMHobOHuh6UhW0KrKUrTJfFRec+x1YHaV5/
BZkn0VdH8sAxR3uBfvw3SuJguHMS6vjb7To/e0X5DnH6H6Epo0iH4MNuN90zG347sYoYjvDFjpeg
JC/cxrreTJ7EUtcMoQ6QwtPZ2WQdTHfxyWQ5CKgez27k/jDD5BVgTebvKr7eN/Tdm3Ik7i7QYWO6
R6w0P1eJabGq+CVRznTxXIwVI6gWkddqcZz0j+lcxj1BDVdkg4FNYZF2oVQiZiYiImeGYoYhdY7r
QX2wLLNUBmUFnbV462SZcbO/OdXU7u1811358EUchc7Z+YBnhmJpD/MipTarn3tSk5fhxGfFZm/G
V2RyFW45n/aTDzcswW4q1F2L5mk1TtG5WYhYoFsagCXH2+I0DCMgVcQYY9Y2KnyUdjRQ123hF7R5
4yDg1nq1w4RrkcpGmqIhsITNMJlNuE+0vf7lPeAtmLiXxIQ6Tz77z3vuZMXMvNqQH3WHJ7JK2wjt
ummXar36OAH/PsJz4HtCiKKSNyE9L/7t9DnV8rsYjBf5VN4Lf/b4VdEWPe1THK0acs4Q4E6Jnvdu
3f0sNgGBTUwC/6EVIUd5LPy/4VE96PB7ZgHxyzCtrCkRBlGEXNJgrRtAqL7sOtyUzYVbc3fo5BeO
SFlKAT+AS7C/uixd1Kgnfh/38mR5p9YSS+ET+u7TlK4b1+usHhd3ohdnPwToCsS/vZzNE+yDH1Te
xFVfS5nAHAVfDxcD2dAjXtrV0PIembp2ssbgPcOYyH6A1+fr7wiZGfbwfEW9YhKl28D7joMZLm9c
aE4+moiWtq6vBnno+N7LPmlhw81furOTtXseVIYDSSmJHktvSwpCacSBuqbV2HLzh7OASFXGcmEm
cRpGAXoqhha1M4vgRFXTFasLm0IkWCuTgO43hGitYPXKsoJUd8d8GpV2QUW0BBMqDDrqmyl/xVUp
tsLYuRSk05mgXQox35HMUKuS3bGCtu0oZazqaI8R2AVnbP06mB/7Elfc7R6IlduQgcJlt+wnWRcf
D0vfhwhMGnbMQ4jOCPYWzTZkUdQeg2EoHgkcJ63uxFVqJ7RjL0GZxHLujlmKyCa4uDtWjWI4JBf1
6hBI3oA2KlbJ16iAPGRi+jImaj5hADjBvixT3UDRnT6U2QykkN9RxI5uGrW1eHeFqm6axVsIgAyn
7M9iLFlhyxTA5yMgTwtv5xVjTgwamsTJ/ppha16QT0x2Re62+FlgT2PQc5QpT05+KJF4N4XAZiwi
SuF3l1dgEP+b9aaHv9xHVWtet1CgKliQNnMAzX2GaHLFd8rZ/U7mjHfabpJCOUqLsB6b1IlKEwf0
IARSUPA8GZnuqmvV57QMguAE7G45GtXHnHNQvyj9CgeHt7bp01FcOaTLg2yZxuFJ2iH7pPNOHrw5
DZTkYDusO9nY09NGqXb6O5/oh8s2skSkhmP52pu9qrtA1FfveI5e1tHPZdNMXlHhRZgNDIKJe7ur
iPIMm2kn8AZHyJziy7RlxwpYsdhoRCTN9D+t11DEiC1gUfZZdRPYehdn+W0AdzVFKo3Z8XzskSO+
LcXABB9Y+gpsMiCiDc6AXoK3KeRoqQKabm7mUHT3OFtkignpnbZAFZcGeiAzF6/21HAFA2Z9T8CR
qXEJP/3kqkxRCg5nmh3fwBWu7w389mXbKGjJno7iJAiQ0vABJ0B4nAT4UCNGXCwTPxUwdRuF069k
CGNagSC+CmzCNhr91CNokqTOlMmCFjTKaBFY/Gx7QfLYC5tyU0MzAgGiMc/up6GMYR+5MIHbcVdF
uV+1jOP1eQeZVy+Q6YdgfoFcctlgiNxmyVH3thM6uJ02dS13GkMJ9N9suy++WjLG8iLRaBIXFnDJ
vF61Zh25tzE+PAtkYxMRSlMy6MB2GdpDAhrBRwq6Cb9TCpXqIplNoKDRARzvy8Hv/wOTIvV0eM+g
ALQvislYycYD0KNTd4VIteCrPOZ3jgLJjqhoB7iNzewnAWqMVH2mgkhnUKVpcx3fne1wAAD+I6Hw
GE7L/XnwubTsKdkC2J+a0cgVvRc5WnTPZX2ntm/TiPsBYfK5erRRtrPvnG14/pmDT+YibB5yuBty
6Qaa77NwZCK3YwPF5DUsXJg0vRh0w0a8YVb1sDDR7iaWyZEPzCYXxxkaJg5L199qY+ZF9dS452nd
UxJGrJzTwdtr4S4DuTOWdebnrJRrjjKIm5SdxVzdpNy4VrEj7TUlQ6LUs5zcywy+P+M6OSiAgevv
D/PK0kFiRjB6i8AgnyyMsUOnwi2fcY+rzpKFGB3vwNDa/bLf2/kClsZ7WYM3Kf0j3o9D2xrRY1hZ
JscfYQnU688QQKOrIw6WzUiBi9kJCOJqq/Sb671cLq88LwWhEhHu+sI5g4dUh5vhwebbHeLsItzY
p5H5d6NQpIDd8LAacTT3gu75F0RLPePe+D4SLQdAkCTnUFwT2YaVo2an4s2TpT7l1XxUpc8JfTvz
QdffjXKWYJE0q3CRJY4bW5+XYe4kqoZcFV46zxviLAvlh4+mtGZkViJz4gOpyCOBgRUCXo9OsXQe
qCqRAHVrW549jr7HS9TgBcWm6l6DrzoltKiN9ogQQkqyIj02tXFt47uEJhFAborKjb2wIkNzpH+j
0TzaaCusGxs9FfUnBrSdMu6aEqnX/pe234L0MqTKxgsRDHoLbVveNre1KluMXHo+Fd75Q55D21KN
yJXrQjQDt+9Ax0VKeB/cg4YY0C+OSB4EqsRxs7UsVNM9AI9/0DnycWYTrjkhxlLTEqoYEm5V+0T4
pw5dNX5UZAAYQbtQwFWQLtpwpXPKyFSinvKeiS/Bgy1FdlEbL7JJp2x6jUy1cpC+aOMJMelY3WHU
0bp5UjoZSc0XJWgi8RJ3VlxqzJJlwFApU7Aw/4HqFtLPnpK0KiBQ3oeRn2F2XmDHIvvoGOxzetf6
SFlzG9GdATThf0SfU0SWjjyZ0y4UeVocVaMDyDCtqft8ZWgJCvbRJ+KrwJGtRd6dobEZcMAAfKI9
3NAHzeOZzMYj++sGhWzXeLeoYBspSMndLOLcyt3OAf8TXyiNGSvUVo5cz0PpWd6ffYnoFB8bzkm2
kqqBEwuX/+Gg2hUW3lZODS/S5fRpyuetr9YqcU+pRO5YaPx26PKn3XkPXZ3zMk0Mu//f9uVoLAWh
i52J8LPjeX1mrjNV3x1cAG7z3lmpextbXMiI9S2Cn8NwkAfRezokbbueBa9avgqDZD6oCHd+1Mof
gPMvVlGOIMfVnEzTdC4BkuXzay/0a8dtqgZk9CrieqlW467O1JgF+RgnoPGJ5QeBI3wEj2i1vi/x
QPkK5BvVkwnZrDytdltS+mroHVb2nfb7D5aWx3Am4diOe9QogcYdgfBMqkOK0Wwyb/lNBolJZTUq
0o6IaRZ4mNiBltBbfW27NrLcLxceiT0QNa+8A2X99iACzBbBF0O/GPDbw52pGGqKGfowD3fJj+RW
7M7//Oe5C/g0NaZ+TNfA7UCAtdWptlM/mZJbeXm3h1n005ijj/Ge9ymWjHdiLeNqkfsY6AqsYvd7
t96mb8kMeRilVHrZNUZpl0HvZGiT+Xka4oQEJZHuTrY+KPihJh5FOPXKwND6J9y+HIy/aXWdvmXe
1Ijw0qr2xtX9lbNZUfYp5/9tLFbJknneCQTY/z1s5w6S6anJmCUKWKABoryrmbGDD4AAB5K5xUJk
VNehev7OYrPIPHM1aYbKbdcZ5s5hzerrrNM+QsLkE4hBTUYTfC04oJAy8Tn3joutWsAZLKN/fHld
FPzxaw46pS3mUg0aHKpWWvqg/AnLz1VHI8N+BeWOlIvB6FGCkKSmCZevFFZ1xmSS5dJtiowAkyJH
WGr/eeOMj8tZBCj1oUnzkNPa+WMXgWA1BBml/0hfL4gdhBPd+ZFui5pmKDhIu3m9oMg7vj4Wjesb
C88I03VuPQnX8L6fnE4fuJtp/TfDm/Cm8xzlIZmMvfzp7ETZJlZ0yIFchuYJCXwzVQAsLMLutsUt
ZksSih4ewmVkif4SO9zlqOt0eJ7hH0qqRu8CR28t4ngWJK/mGdiBYHuuwMUHHfdGsETZm65iSm8h
0QYzUIFy4hXtfvHNEdkMcvamtDYOsK4gQRpjbCmir6NiO7lRyacKsn42fDpMh3TcltzXxMFnd/Lv
1kr6WsuphRZvQkF393EvgVYfIm3/ezzvYqe4xyolnaIZc4wG4e6XBmWhMSMNb/+3IJfVCsObm71K
DRy8UntQL05MwQyVzOAouNVBgnaRWvPRJIVDiYBzsqOSqOWVS29Z2YanvwbTmj2CpSaC3wEt/8Qe
FOUE7A8Oa1byBxUJjUiN0N7AOQzWB6mIBTRnmIsjuzN14gjFU2WMw2TO9dHa/6oZVzXvIQB/P/Y8
+/u1wHTVEzyjjQvV4o1t/G/Tt2h+6cBz7IkTbcziDOnK0La0FI13l7ucjBTnhb2vZOVxqcv6Z72S
Upkw4Q09YqFd+BUUC8vUDAQ6hxghhTKB97hn2zKuYEoyxj0hTYHRFAig7mtSwnaLjETUbl61LpEk
2xYRc8RP1P3ZlwhUOQkspDGbW19rnie6X5cCnMGdvn42mn9Ouv9bnPDMNrG2nQA2DCKpwM4FvgYt
LxlrbCmifdYRPcr0ENYXHaruX9kqJXBIH1TI1QPywV/O8Y792EINw34OA3Ubf6aMSKNqeVs5czbB
Gi40g8drAwS3EP7RbNg1wYlxq7uWheDNORVrknKEIYKC6v6mlRcx5tQwicGehtmlr3fO4IF+I95y
osUAOCILRdv6LNUVDqdubjS6jTIfkLawPhVD+L3F5s/9Hsp5FqKao3IhAlwRU0EQaUXY2eETCTPH
Ylfb2q05XUbEEnLDBomMHmrlk+c3sP+z+l45EdRRj7V9sF5UENuyr83hSTDA8RGB4/mi1iBSoDkT
G8g57w7UmhjgKHu0K7XTulQONn8N1UJekNykqloqP6/amQptesgU7F/GDMbFsBlHF853NROXF1Zf
JxAChGgoRzpcTkinXksQxREjQLJET/rQGKxue9H7zSef3InRmE/Ck6pqRZTelKgil2JBxsff66r6
q0mW71Y98cGhTIITlaP3H3BMhf6+zzLPjsim7HRLp4t4TaP3b8N6mA1247+QdJu59NBrB4zF2ISM
0hboh8xo6+F1aXPWNGoqSeda1y6Wbt38Rr8Ffy7tFM1SX6uitylHTlKbs5UDquee+84v0mqE8oVP
Kff0UfiPz8yLPnvetzLU2ZWCIbMGAG/MIUj6SCdYlXNXlakVlmMVCOfjotQ0eeb4Yv7qHLHPyG0a
HHb3VXsKH9dTXPllZWwhjzSU6oEtzsHjHX9suSlHz8pIB0ast1rgAfkuR/f5lG7kQNsOt2g39rwc
wYgLket6qVRynqMZEPl//MWFdJNTMGaIcduqW+q/YiMnsFTqV6eVF584QvCZ7M+wcClmNwH4FiS4
UsiLOY/8Pn80Zyi+x3B64+qP7mJmNyqit7avQMiTZToqvWL9S1G7DApn6c3QLcvkeKzrVq8jekyF
2QQZPUmSnuQIu/rVXs/mLzkY+KMhPoXJMkQ2+1SPl0WgQ5ZwTE4hkJOCGxMJ9CDPVG0FtbMDKLfR
ttYG7ev9WOWqScVowAwKhniYQf7ktyaBWFTIzw579kQZgRWBlFS94CnFyO3tKqHf/Uo8tiOePhN8
cD/ab14HccJfZ20D/5PBrl3WxBmG/4dDYf81bVPUtJqgoIUL2e7vwU/1QtlbNtWbejim9b+4lZ12
oQgFhi/BUEV63Skul1fci9fMQLX5IqKVfmAyQOkEJjU6/4hv3REM56mFf8D2nVe3VXqeygk5fs/t
WJtWbG8f/dHBlr5yrsBvokK1l7NVDYSQMfNwM5NyVnegBpnocDjHBEppDBFjrih35xeYBt2t122O
JhQu2+JukF+n7UDy/eiBoqOjXH4E12nDtp4UPRhgxV6j7/hcLV9pPrzgyumNj2qa6FpvIdPU+7zb
jyZlrAf+3xiAg71o5SIP8rz54Smk6U9P43vW5WVx74Ig8CkEr/EAuHEd73lB0XmHD2UXMjsliGUl
H8rv9kcdmaNpS/us5RoZr/2Wxyj+plPo2+MX3qKPq9DNmp4yAlj0upiU7j4cTuMH582JIptQrcTz
uoao6UJs/MN8k9cdzY62KGgy3E6M4SQXF8xXsyVoGvnA352mXaTmzw3Py/sf4T3/isfcL7TQ/2j0
NGIIo9JnWsI6imPgF4gRHT+NiIU/alQoUkKNmasmpVswKEKmE0P3HYIOOhtjYCWOQnVd389f9XMk
pElYJ/ZkObhwSBJ3pqhl8lliTMGALdEK9ECDibkEwu44wAajz0WufgB9+64IsBF8JmUmnooiCSdA
EQTJp1HysPnpttZxqWBjaYDBuQQAhF1Ij5wucfqgsm7TkPRoc7wLveYHSRBPLW+Bx+wmh2GMB461
EEi0NiCLBg0NSRI7B3cQnziHGsEbDhSjH0gPxfHHYnS9G8KjxUv2bbOm8x4cHrWOHhxIlJRQmu/8
MJEH6jmlkXaAjGYcGbIwS2PJFTttNlSV74BeLZIkuhcf3GWf2MNtA3KTS4ClPC1UVI/N6bek421b
pH1fc8D6zMBAZq3Op8Rf0k668Zvi3p9im5GimCz5H8S57tZsM/EzgIyCVTLxXJzXC4BhqTKTN/K5
VIiYvInu0NimE4HWHmNOnHAtEzk7W2CD2GbEiYZVVOUZiUD1J4PA3SQis3PIZHjouFEJaq2gK2AQ
WwKfLOj985sOFvLzX07fWIU4RCjwO551xjuKjerb10zGNh91CH7oHCCotqtKCxnLO0tpT+MC6ugW
exWb5Advz4pSJv40JCW5VKozsumfj6NFj0ZEciw84QBr92EnsYNA2p2ax9kVeqH4FiyjIlhWLKbM
LmB61l2Flbpkry8aPiFAacFoaA8Dno1ujJmu/WtKS9m9Wf7LN9mPxnpV5TGRuu64VdKGLZaaNf2F
5fwd6sgcMocsI4t/Yt6iLhMLqbCkyrhimMyOjsggcGJRQzDtafTEfB9z+qYWLJarOGY7lR4ku9hd
7PNDlYJ+WesCbTBoiFoBnC2z8jGmRjfOYrOfa6GUkUZj4I5moTasr4E5VQi21OtaAKUd2sLt6Q62
RYS0ajyDlWDtvEitn+cLR8fPKB6wnQHr/f3zyzrdsWVa+i81VnlCCq2my3xx6TR27H0DHSh2RJdK
oFrC0AClmCh3YsGH+xCjzyIbZBL5l24IiE0RKpPACFYpjekVsiW6cSmBSBWmcjVr5h35oaLrmUT1
I21gOqnLwxwn0bO1IagbVyDGO+WE1Pe6tud/NXFFXXAMHHMBkwWzEN+BXZUmSkUsHyvH6/QAi8IE
c0dfX0ZeL7hCeKgLd8p/SX7hNPx6fjliNAPpAShmtU7zkSqZ2hI/cTpzru5q96Vx/rKRcsAZK35I
AE5pzwxUBTZnNJkBx4IdBRHzWxYpzDqtVfhdYR9WjuLN7HiP8/kj2hcLkNx1AFP65KHjQuLu+fWn
Iny5KdpE0I8SvvdpyFWtOhMhrFGdGujxeuOYQ0RpPFEOC+gwdbCrgm5TZsgvqBXF85Ta3ytU3a42
4JIvDeyvZo6wcwC9MP/3sRF0J7PUz7Z2JMqXMJ0zxpMZTXAt8Se4NzerQsBAZsh4VvniscfLOp3O
VWHUzbAvUieSRXoe+XVBF8XMUpwzIEZe7c8Oq63F/sSjlTnkZZh6RXA/v1BUpUSPvQf7zqWVyGvS
BGJkxbPWoIj0VsYHj1Lmr+WT3Yc0KhXndUpRndZkS1rH7aB0YL4TeN/rXUuAwW6w0xdbo9HqI2BS
5avZdVf74PvPKdSd3uo1fKAthpMBsVwLhNltmx8vD0IrmyJRDHR4szdYThlXxBH+MXLbInojrEsi
rKmcm+E8Y6tP4UMM4iTUKoTQjgCOVDf0z5/8t7yvyGn/xWaIt5DgOWeZT1yIDvnTsv8Ls/U2UMgm
dG47XXMezvvUd4MNMq0cJHzM0bzlabOAoEc4bE4FkId396uptHSbfMpagF6Un/mhhvNpzCnJp0wl
D+lCRJMZ2aQ/wblin/KjLaXEWSrbdv3//iMTx5es6cqk2xN+RJM+g9TUxJupRKqo1WoHqDMDoG7P
0PiOcSI2CFm9Qg0vrxVgpJzT2sFnXEls/hnd62v8DPjuub4htE8q/c4wcSQL3Z5i5IfVfvxgLmgg
5UhCr93Ys9uVPu/YAXwyFAb8b+tQsBvrGHH0T+8m1OAB5bNvtZGvspMQcd8cuiLREGnWnkGQp086
oanxHKReSwBivkkpbIhmgc9r8YHr7tSfFdyjZJvEvxgK9cUJHL+ZkONdrXWPmM+ks4nj2AxrM3Pt
Jv/vA9QOkGfAO1FagMwyT/DZm12MSn1WvfT4X9AmlLnB+hPjQRIdPvrIlkQNwu524qSKi3haVjUj
KptyVwRITlKJ56bBScVVtVdCYsrCR1Q6eho0Wqg1netfkd1hvj6+WK3GAmXs7h4zo/1QbjmkDq+K
uAfdlyzzBqzaRQNSGQgqVM2FC2n04Xyt0nVlaNrmvgIlldIYn4s99RCoaYpKl5gGEOe4QbRbJcJc
VL5Wp0meYEUyIql12ZGzyDjMDd1x5Wj/HWsR8d1xnehOuPIRX/2HhRaWi+PxA3EcyY3W4GPiLAoQ
lsbDZRERgsk+zIPZ9OUNHRsyCxQngv0J7IDhrdoVP+m9YG1tPYHrx4OsjrcFgLKZwnMSU0F1KImr
mZxhCiZMlgNJjKpKEgAQWzKlZhWElw72vwp+av2PEZtVSKXvEGgwe0GW57A7JBKzWMOS0pXQNeOL
LYmP0ZlZEpgsNVDGeUC/Nj0bpMTwAo26BTVJC1e+8SNXpiDkLruOB+Bf7cUaDw8x+PYPp7UQug8x
MqkwY1Qemn4Bck/cuJCXFvL31D6E57KxjMAKs2Avnn/v9VVmOk7ssU2Wyu0RrMEnGMjRZysprV0m
SKWnvnzrPU4ZhyUo2RR18Rm8f2dhhULlVsmGfaYFJc/02Dh5WNgn55pph3jweeHtY3F0c01bjt9P
KdsakpDu8fgzJhHIF5jwowj3xUUlVCe1UERQqP5mwyaNu3QydSrC1c4lZDvb+E0KD45iQiR7mIsc
/gYX+AHEkfSBXQnOkQz+qxXaZbqYTVSCw0tB7XqM2KZVbaJjy+WHva1aJkj825Moon0u5qGi6N9W
1V5oKYeklh9uTUVg+3XtzCxCmwLCIWen2C0I4ag+reENnrzO5mDFtVh9N0K20wrtv/nuS6R/Avqd
nYPWxGaugsQsxMl7HAxyeo+Yse9p3r229F8pCCNMSZpvoOFaE3eb+cP8dVn3agdORnHBuBmKD1bO
hfaXxxO2CHRtZsowe53VXLMuYDOip0avP3a7nd3CN6+qwb/ZcukSHZpfQCeuVkWmsnkLh89feKSp
CHvevWtBDBQy1OIarsShUsdgY1Zi6zndDgRnNj3yR/iDEFc9CKb51DZ9TYYl6YTn2yieBx10BR3r
Gt8J7gRHIAfAE737dmb13w70uHeWJoDIAAZL4yjHv2p3V3pokWHgF4ypsdNMVM7SvlVWgEBEw0Dw
0aldcQzAx5BsNgLx7UeGNNkVkCzZaFfp1t3WwydSWluIV4FaIVmN2N7LCVawtZtcUFnI+yyWt7ne
VpXQIyyeSUOCTHcC1EfxBsnev1PdErfh7KaIgqs+FIVSlzA18Sh/DmLJfnMOi1QIWOgRsubkoOYm
OGwNq4pNmqmb+EuIhOpikQ5cdGWhDNsFR6u+IHy7FHME+aMNnqjzu22je59gzMvElsl/5gDSKjtF
l8632Fnqt+Vmt9W+nAPa97/oZ5jR7AbzQbyXD6AYFw9xjwPOUZ+9vpUHl2pT7GCZMI6IlkMVYUvS
I6qoBaMJyQRZ/cYwU3nckH8yvfbKkHI9SmXgO8hrMSv0q5/eCIbH1pO/g6TDAcxoo3dweRXY0kh0
rjFExGT0GCtpiBBmLVHJMC98uLee5osIB/6jnn8ih5XfJh07XgGcIfMyHGP3FIbmxu4Nwf9Jy47+
uqRpjE2g2sGMC5z29kpaVD0UcoSqc7dbOJgyzHhyyOtlwyRGTLDxniliU+PgPfG23tCMQjtYyj1E
N2IatW6tVDgbsyium9YAQxWb1htcNWXtG8zLR4rGHWW0RIO60Fv3rulyyVSjzt4cg/LWzWrnjx/5
7mUAkTEe/BuebsJ/Sdl22qvop7pvxtfm1znHRdG9x8xzCV6nJS8Q17NKHcrUZE/wWqEHBpEA0uQf
A9XtRQkyxz9neoXJkHYZC5/BwRHiwWsGBjDaMpTb0+IqPIlz7AfbEwOPlyrRZdd4QeYX/mCCi0Q9
u0r7juSbw+lsGHm3cx3FnbOUDGpU0CIsmb5s8Ma4OSdVaTqDDpVrtMAy+ratdP8KHJSsVty7OE03
28RP5IxFcAupLy9MnRlkn/VMkxSq4Uft+mlix55WNggDZ7t9l5wbqYkFdt98x1B8uY9hV5b1p2J6
gCRm8jBMWA7UlZ77MsUzyRBwuB/0L6BUdXLbNiJLW6BBS+Lxe1rBfp8ihsFyPxG8ppkfKESUaQs/
Z2KpL0PyAjXxFlRNSOs98RlhkPPY7twY1e2N3nW9gDPc8UeMoYWCOme3pvs8sIjHpy+2rnmuLNAG
05PCAUQ5PKFfc7bzv8LOKupbSPOm/FFjH7jhrvr+W1eEyCspv9HmQUuQhp1DO4NI3qDplSVHsAIZ
UsMV6gUUBtRAgw8PJBAm4U/3yRhw03OBJCjPDaK4ncujAq/t89eMMXz9MdOuWCMjIreVuovEvpfp
Lk62DdpKEdJkpGqwvHLLcVWJ6QRiX9VOmrUVF63a8hCrnoH4zSq3XntjzsEcOKOsFCwQfaKlSNZU
CS4/9bZRuNgN5l4ClQe3m5tPV0FWL6Ndxpn+e0onRwfS7V5IltTaVYmUQshPJm4InkqyygDi11Dy
wwakHpp3X5SUaStEd1XuZUI4t2z3blzaFmKDE2Xh1jY8tu/TkYLL8SbPCexVYjP9aSBnLtJrOqDu
aOQBL7aepWbHKfz6/mP/hlLh3VAssLR1Eq6iHZhC8lhRLZzI4Umu/6G3gU5IcVzXmJrHf1XJuEls
Eu4lUdVnAo63Hb/y6a6xAqqCrxOMlex/s28XJgTPjyuCtkG63TGHGNwe2hU60OH9Zy+ZjOSHRmd9
xJBJjmKZoPCBZ+QuJMALkvEAzZTw5WMmRwthchso8XftLvQOhsFrsgYUwZfQ8+G6L2JVGPBzJzIH
U5N3Gf7CfwsodtWjkHcHhtM174a3IutOSxOllXCC9dIsb7StL+KLyuUrbYM3vAWkczJZNkGeuGkP
FFWKJpgti8+ulGb2hoHjo/+y5Chx4tvEq5NjeixthnNRxWqkjLzO1+3xADnF/8I2wO5ROeeL12To
gc+2qLWgu3BW9Lpi4WgKCtD9JO7IJHj8KrfqDs2X3nRKIOYwf64sqXn5QaeWBcAEQGmpneNPKLXY
3MPvUbx5QjbwiclmytIk9VpYQwIc6xPGslt3iIhHTJ8CRj0QDDwRYu6QhPAUn98GxJJJr1HT7Hcj
pumYJ9Iyv2DQJ+9MGV1BNffRx+xsIvCbtFoSyBULE2wB5d6HRg361jf507eGTVV5TYRChMqEd5zb
jZqMBgWyGAvkUlKQ1PpUASP2T69W57Hwc4WR7d+OFv+l1PhbLuGm1VviVuet7y839Ni0Q6WdUP28
JoSW7O3bDFnuP+rETZk8Pn6nhsDSAaFj2+2uYVbbwu48LT7ezCEJT6u72oGaRGOThOl1H9cAxUnj
kj5iqaBkITQ7ZcRxN/G3V47AAeQDt3YM3yrzFCO7wwjD5U/VkRzUY/85h2uqi66uGqY4O2eZYd5G
Cuh2lLjnXtPlYqdpqGUzmmobuZ292+aD9mgN0ajU05HNzyqCqgoPcbJrfUl71Iz3IuFS/ds4PYfO
uOdhykIS4Qx/hVy1HO1QJ+1MW4uhG8sdE+u6dFav9PUn0hukZB9Tp6ocq/QMrQuGBU+vBik2Hm+R
1rz888glxezLIbdWweALMOU8E8v7EYBOcWt9FI7Wgvj8Vyn3LT8Q9ydLwuJCAkTh2JKUgxZQCU2A
VMQvpcdEWg6y76dbPC8pcyiuygmOS+Eo9hiwsgmkBeyf+8uP7dciMqL1jbIf4bjwIhOihxTmAXe0
u4UBZpEunjpEevQLlB0ZkUzqNw13swsES6Oz3do7GDj0QFUWHBY212WC7v1XIiMRY1mUgc16iQFy
vKxkb4VKI1WFfvaRZdZp8P2PwJYJN+EJaFhNHVlO37ZGJQYbIVrgSULQ9kZQglGoZ+6MEeKr2sC9
bnigOkbVf8L/WqhFRaxYxKoFU4P6TcYftGrUSs1DYkHAoamL6jpz3r5DjbqrQDA9S0+QsngE8WAd
Z6DZca+OzXe58jJeSfU+gGyQzENPjxUEmd/MCEiWVvDi5XEaZBSzYpNAkPGgWyWa9B4s9/bX5vow
H5oie0cehy5yIUpSHcutvV4dF0IM5RvqomHaP8rNMlZ334L3lmkaykKJ9/8WJpLBdRFkHN1lMdf0
5qJpoLLrkJmuV58VENDQfjMWEgntvj7T+tOepkzhzrWGLA8dn02/6tq17xe4ZvEKrS5CQuix+pJ7
5eDNzTfl2iCDr4eFH4KgFEVw/xZYaTpIGh4wc5QfE0Js6RGG/mFs63UHib+lBcY4KXfjbvEzHTAF
hh3jZFiUou3WG2jQ/DJubH67QlcToSoQFz0REZK1d+ENBXEjaFs32YHyGgdu0pqHRS8LOFi8fRh3
Pv2rtCYwReNfQlX61uV/swDrwxgpAUVoT4S9091yUCLbj1RRweuIz3LewY8If2IwtXpW/NyQeX/h
+6Xuj0//TcLzhTnLGFn6TTmF09KOxibllF2jF9UNiufBy/kqfwYE0rBX9UiJfdBBC0tUp/KMA9Wy
kolQxXscHpc0yGe3HG+xnyAHZMkN60G4ufEx+Lx9YvKiLYBkrB/jdaBR54ufHe4+BqqMhwY6QOHs
RhfDLqlL5safsBcVWoyNJ9uBswYjEfKEobn8jfzzpjhjiicSr4dtrXG5Z/BEwCX6IsjlvSY+HaSh
dRAcAU+z0KPSJXaDm0+cYtq7CXiMoYnqPF5iyym5f9sKXCqOS4uMrX/H/uXH9De2sLbtjBv1GFSY
DcKzFiDsEY8Jza4t2sNw8f9IdbDdJVdlIDrb8MQ5+k14N92XrDpcINEin7qxQMvdCjjSYT2wdeCT
9l9U3ngPcT+abkSmU8i6MbngZGM8JlLD7M4qouH9oTT9cU9VpfHtf5RiibQ0vJRvUop1yul3pKSq
ct/nGrQlHb8dAoFcf5ikdszCxoqQRb/WOrPUkCo4igSBXx6qKWaePcDG9LbaaZtlW0gUeTURCVu9
23sPRfT6YBmZuRoHTA4YNEZ9abJ6S6tJFsYOj+thfXa/DuJ0tUm+pd9DNNPf7e0pEyZVXPMJwKeA
DL1cjFYzEIxV6oY88Dy9j25xvo/sbLie0CnkA5DmpOrKyOKA5XiqzIcxMBEbLkCMrRw0JcpGZWml
J9+wGz9AvvkAy0TcVD8vuRE7xPORQLbG/cOgUmrFTR/YXt/YVj3c3RcP4kp8R8W4NSECKj+/awK8
Nyhm2kAw4PJfthKNKklM9IXHAq4m3Ggwch59Ld2kj03rOWuPPczMK7rBJurvBgRPHyKMBWcHjrC3
M5MeqGN9nOG4jL1TDqqrDw7ZDGcVbVsDBi71Bz/N2b5HwWFFHrydoi9WWVfsNsY0CNZ4gMUZjn32
7WOIm7WhLVPQoq/b1V+So3UwEZ1qQhfkQFd5242UVVQ2PUL+9DF6UaUTBsAA5qMtiJWpgOHEdPnS
tEXXe+RE70t2XpE8bjg2OjSDzEvBD3U8UAPeWET7HMhOKuL9GVsv2CJFTagNFzJrILDkyFoqj0pQ
cS7MIbl+O9Ii/U2WYmLD+GKhLLDliywJpfB6wAXTIwpsJX82MSlGUWAoX1c2BG7K9uRDZQpcuzxN
wGGSZadm3Qp4gkDYBC6emZxD1m7/toSd41DkHbBKzVSLLi+9dq2xFUAVcspR+7U8B4X/vQm4Cczf
Ld/ihh01Cf2nYQaF2ykCVuNYXECVbHpE5RAA9fdVxAZiY2KE6YII/5OKogOyLNVDgKs2GtKRFWik
OQjXkagLub9Jek5x9gKnZdyUFPTP2FVuvSNDuQv39EC23MtMiWDziedwZGqDCIlJwygSlHRKyu32
Axv7C/0QsNi3qMb+vHly+ka23tqpku77IbwtvqXgaJbCihDsswY9pxXeiJjWO/pPuYWHPQ3F7641
LT93iWDW9mT98TG5POSXPCwQjcInmbZNuewtvBfBR/TlBit59nFBjjzfWPIkseD8Rjm+CcCZfdae
Rfy3nmt8D/BVzupiiXTwC2HOSmeLhfxaz8TmbRgSjfNudBRPBPaG667+4JVx8JUs8zqZ+ottK8FN
tUCXs9p++Lkn01vGncicDkXnn2qnQKM09kBNFGOiXj/RtxC4Xa88qleyMO0uGM3ikuNeJDQyFrxs
weHl028OyBENB2ib0Idu4DoTpXYg1T5aeb12XZhpkgb9BGLI1kZwc0XQjgR1vr+g0Cwpqo+65Aro
afJCEj/yMGVp9AZtRNsY5LoTR1iLydipaCtoQBpTCP3l2Kk/myZoM5Y/MMl8Xkhwx2BF3zBvXHY9
sibg1Rt+Ful0rUThIrKowHU9GnJk4RFb0gLIQ1psdM775AT+2iXQPmlnG8iQCN/XLAvI8jdcdSgp
7MLP93H4I7X84YbIFVNZIB8CuHkdw9VU/Vm5rAfUzrv/+Xo419tLSptxcwKDSWcGjnqLP+ycyP+F
A3qiyCPwKF98SzneKK9M+grh3hza8msgBWisPUCCW2JQebEKHNmvg4ihyMhhgSOAYkUIWzisqP7l
E3mUDpo6wsx5jnu+11pSyBIUDJiG3Nhw1NUk5m5XrviQR+ltHsIhML+PDMQ5QubqX/UsawKWgZQ9
t97aH+7Qb00EZ7PlMMfdsSQF+Sjl35/R5NAAFFCTYwiHPzvzlNLVB0s49eNyb4/y6fT95XKBWxkF
Lvqiao+IT8CXA9os00GSOUotMl3jp8Yz6xu2AL2fdFChG/KxaKfN9LUF+aRzUu9TY20pJiTTfXe0
ldzI2l9PE8EVr3YEbSrz9vqeZmBeHT/grqSCd3ybH8iRb3o6KMiuOQHoiAWhdHzMyGjqhhVE/dCz
BPrADhiMsNVkuMyokF4+zHOu8hUusBoKvxm7IkaOnUw0L/k1UE2qX4Az4LThgI9IuVSnAEwSVsfL
28Neeqaz8aIXU/bRax08mIyfwRkzZ69uq9NYbDFZ78MLPEFsPZVP6vjhmeHI9kEt24QtOYRS6edz
2mGUXqn1h5DVwGvPJHQORr3wF8+fY+Day7DMHILuqE63cCxdnKrHorhXUyVE8wUoY1ZRQe4hr0Yj
Gdb8Km6frOn9fd++kZfkk0MTnpaBmGpeSliXRlYT4tGWuWv4+BJspV42wtrJN3dTizA/slmkiCgi
MItlBtg7IhvQY7Xwg7mEM3mPqCi2HuH1OakpKiahNkvbnKVzETwj/W7xj+ZiOZE4bqYUVEi+RNir
ICBj0GvjRUQyeiv0ZkyjtvUckEOR6N+OPP05HMGiDYj4plFpawEZj57WOpYd4Y+WEX5rOWvb5wEp
JX9HhMzASTqqTjdof5vWNzpiD/WSkhF9eT/NBynjQDb3pdNu9HLRf1epZhS+J3tPnhBwAIYmLqpD
8DgIkST3glOxxaoOuUszA+oHVcE4FZfCHXXP7tybVuYmElgaJcPQX9UsjbOwLW59JoTDPHSa0ARo
qQ/DEcDoVyiR4fX/7KrDA7/C+0huf0jDc1FDOe2Bd3WDhOG4nJjVeCflZZHhIYgdJa5ZZO2OQNNx
g8H5ac8syWuLOJiNAloQNUswE4MvlR+1DJRDKlGTL6fk6wgLIsaNF82zyk0giMui36QBY1TAtqtb
mscErGzpibf4KJ8y7E7LKGx4l9NdUOfC3olcFLPevgoLDqHlIY3Ihx/dstXMZxaTcjN2MIIvpdbp
I37XPEHEL8iTGOjxDBmJJey1u1SX4yotnKgm66bzeqPFWkMOJ+e/987AViPeZvm4TYLSdviKyAeX
YQfTRqDrZg5E2GVKEB1pk4s67XqcYhadvYO188ebg2/juA4ugBOUnC0dVkvRGMq+C2uYDohGbrgT
ChifyqDX7ru5FjuCIj0l3oHegvDVgXRic9Wy9n8PPG2apK4h77odhQE2hXYKJ9pyYkGH7tKhiUei
ytZ7p2v4MyeXglPTxRFYYcbe7Wfzj+3JFt9/pIrTpRlvhhGVrvExN973BY05GxS6H1XLxEIWlWoV
nMNZ3n0jl1oY7f2Q6/56Zqbpba7gEHF/KdaN+H1uUBCIjpDOz3Fedirq+h7em/b4UZ9gBJLmWmHT
VwqeblZQzZjENTsPpB4ZygKx1fFFKSd9Fyx9F9aPw2+oPOjKHqomsTl4ssGQhaKB84CV7EYDw7TD
t55Z9qvcdMdeH6/wpir+PvM7C/43QhUtUBDhbeJG5j84LimHePBr6+ZFIh5z4v1pJnTtpwBIzqE1
/4jtYX6RqLSl+vephb3/TtHxFWneFv+ctSwh2YXs99g49cNENkk9+qZ2g/m72m+NNLBrDFPu3cWz
Sb/8sa4ORdVOEq6zO3J0rmQMnlqbtulm/oUXA8O9MbAGO5o26sbsPKculpxTTVUhz40eJS8hIR3W
c+MB3ydgkotDpZo5iRAw3f0qVo4Y+QTpAm4RXNLP44fgqcvGHZCcoMulOjtmAfFNBnTCZACyYb/C
nGXg84mSxfL1QZWGkXNUKxdsTDmulQR2W3ghB8Qcqs4Ag0cHP3H6/SAVoubxU4/M1SDSxMGxpGoT
22XMbGW7SXplEAB26Yi0zf9dmxBjd//VopKxexT2FDiSzOJj5DVfK0Y2toa5Y7QLFwdM9YlHs6v8
ZcEyr8K5BFqSU99YhAkt8UCaDNIh0BcZexzYw6Rg5tfS6n1+R25Ztlze61VubKFUrSvvuzgULyFt
WoPx3QTlzz1sQZXMuZK8U7O+Vw3ohXHB+SHYc3UUy4ZwxbIuJ7E1t5Lw0Snl4Va8rVDkgD8ZDkrv
+m6pIqG2Kp8iJneX83rCcuh7XQbGivwMyOSUmiOj3e0Cy252TbBkkfhbWhDhYI/mIvCSHXKVPRhY
K95HcNX7jzg6+yWqwNgtUTjFF0n9gs/F8hv8T7KhZvc6GPiDo1pNjhopF/9q1aLV5zpjf80L+K4x
UmKf/bFEHp4JNmSY5UIsrWH4F+EynWCdaT1exKRIXakTciMeQgsSVxV0DeDG0crJqf2RwOnWp26n
kfJ7hUfxNrtre4UQaLZjZ+sCVaq5wuHif5ppYrcsLZwfT6hpQ9BPPjDRStt3n+RTL8VhxgmB0NRY
3UGMaLvVgJeDiUiIcs8fBzsr9KN6aNK0h/zcHqyZfTXlQVsiOloQpEaSMUNG83mYDkqxtra0rmNb
GzwAYqjAZKJVHHwXc5tEDLnvkHRBeAQvXUkzNPy0GtSFuHeuNZ/GazFplYNOQCaWj1VNZnSrv2S/
XPRZsLZtehaY7IP/7E4DYTvh7UAaJ7KBViQjTuTf62cGpuFFrfNEjz4A2v074pozUbQSjOvSVwO4
QDQTYLv47WMO13eCGMKVmljc/GaY7bb2wcgo9+2YT4H5Wh0GhgZbd1iI9hUasFMpwBJZ63seKnpX
LHCpae7SbusCtPasRBixjxqMlR9nyt3ry3F8+UvlncDOqJghaNN1MiXr1aVeQPFgJtO02tfV7zx/
p0zwT5b7UGj/bCyS37m1LWt6dyf2zvb6lUYWxTnb1hSsGxRv5riIwekbK2K41UJDL2mqKLmPJjq7
G8PELzRz3M7wLMPuvYZSky8Q8ACbtmMP2LsUajR4IT3WrntRCOW+alYGBilvWYacyH4KEJhxsQby
hq71YocuwdCSWYQG+CLkfKxZ3vsY7j8ArEDcKtTEENZBhXYTXrazRjqMunSrBzz6tdblD86RRb4x
itKL2UVAEll5c/SGtg9ZL/HE1JW0pbBn2BS4lCJh3PH1dDsrjMtQbScpjoh4oW24A7EtuLe+/eUQ
xzBUg4QUF++WMcyTN0jgBKoKrEY7Gz1yqR0Ckss3Q3oMioXHUA4FohwvtFYzdbwMlcXX6f3dKEnv
fXfEkQZYz93Kmd5wzWvPjHnBMoQ3O1eisowv7sH2TJO3/ssRn9mu37f6R5q/Xh4X8jnW5MedlzT5
7UTrESFED0RnDw2OCB/82GEFcGRuGY4rbYiYYvsrqnE+hoOG6wq/u6+L8zH4OLoBgYVXo1iRnt+p
7SgC8nbTO80ARQhb4Og9hclCIcbaSqZkGmJKxFT+4X4j/kPpKlsmgZR60mz8fojtbye1ZdN5ICnr
mczBYxZ+CLCg3CeFnb8AohXbtJbsUI1ufGGrsjvM2nBPURMCB0hlnzAB+tni78Xc/aDI2NdWrrQy
4XWLBmSkXTh8943UjiBTgvnfeblSgCZZBj7DnncIKi5BbheokpKVqmcbc08nuUvu9bYlPSpImTC4
3lBbsIUcj8oxkKkRwbtjsUhTuAljupMtRLcT5YTuG2tSOqR2C9We5DagI1rjzZtLGWhxSI3vOh0T
EEugBPjBcdPqb76fPP9BqbjCILYE0/52AaW+LLpSQwAtNbjTLPdQnK7dJXUYExz+L+Y91G+r8unb
K1w/tvmYeeNpr+duflxhWC8UTQhaqzDN1hujHMprglzRS+IY6aP3JcmOzi7zxoia+KHnDeuBKEQl
e5jnGN0tWa4b/CUzD7aB7knwFksLk8YecFOUMy1YbuDFDs1zor3xqikf22SmOIPuFIOs3l8sJmZx
LEn3ijOr6SD46Ief0D7bqzXxL0PGBNg36UX7ez48bzypcpVdg62fw57NgORrYibvJ19Upsox8YfJ
kaeRwDwCoHCfO2+MSAPvxMoXh7RU6PaOuo8/YcRctvh+8aT3lrNxpOQXzEo9lUwo2fR8tVrRHyHu
ihg2yvStylP1AesRn1ZEszlfeSbNBx436AjxN71SjUUGgfav2CazYNSBxb/pJ4IWOtsEQIkOs+57
QAlpzQdXAEGuiWXj7xVF+BpxWT7PmlI5K5J+dHlSKws/T2ctXq/eNY63WLyWpLNy2HmKLk/HB4Lx
eEz/HOCjhNLNqv1T9x6yV6PkCEf8cUfP3wYcs5NGy999Qw4XbgtUlEYo+GbFk6KeOalXm+Wlbspb
RJB/setNgmhClGT959cPRh8GKAMk4n6zKNrEt3FM49FwyUrn9hnUvHR/U8BCQfpOnr6sQiJsBxCa
mCjwSYS1IobuqVREJixUhzZ+o90yTAIkx6ZWi2i2nJZQJ+nmJ8fHgKmKwzKece7nQq7zfIO36jZe
vO5oLnzDVIizR0R3oLANCrJT+x9ubgMRT+c6F5shKLOGY1JpUojJNyZB0KVbTf4Wn11ilv/aoiiG
RBKF/waOjiqbKC4kJvehqsR7XbK8tqMlLh+lxogRjDrYelrimMdgibYTJNkkiZ9uCwx4+Ct08/ph
k9EN+M+HBrXJ7s2PmAtegauaf6tzcDozp6PFl+DX7f0zAF0uXwvJOpQqetKeI4XiLI3ueyBQI6BM
VBNEQ/5Pw9kZR6k8hKr+4ieNdEC3QcBBB/xAgn3luDZk523B0mNBGzkjCfYkFq4L5uBNfmjOu9TN
NkyJ1pRmA9cElLMY2+sm5FBJ6vShN5vP+sQi4e39DdvPHzzLYBMTVTWeFkd1maaoSyO3mJYqrUQC
69jxYaAjxKfEV9X29rXxQalCcmHE55VxX+MMxw9LmdBH9qm9zUaEo1EiWh0DaEqJ1GGQjT1r/K+U
BHG7jHJmYzDgNKWWHwgBDiUtx7lXgsi33JytEf0YBteG0RKKPxkfz3JNvGxJC80f/BsKXXNvxXmN
pm2Toju6+k/aYwWxUTEZ9KUjSeBfmgDreIxJEzy1KEUI7Qu+gZnmMej9I9N9+qjtXunPCy/wlvtV
qoztU2n6xaa0/cW5KUlQomUhDe++V0JUawPn3vPXf5abNF7Q4saa8NU5m2KW463HtNNHeJdnHUNx
KLFKPotlUamKiuQvIng27BvBTyzM9MSESXal/Y3JbejQk6n+i0Wcuz6/bru0Z1xq3/AJx3XYt7T/
w4Ynfumk3iUuW21s+LPn4BKHwQiKk6FZYHAPbVv8j0q9Z7gssRVKprzydv5Tv9k+EDLBFR3riyYd
NBIdSM4960iRip2hKMwwjsOGLak8W/5GL09hTzWY6WI4yR05mn4iSYpxx0dXVXqkTagRqpbZWQDQ
wQQOoPl2fuB/w5kRLocTuOcK/2dvtQ7Ij0+956o5K71PI0nxYmGJl86i5jXXqAOgUR2r4N7hPPJv
rVlIIiVUdrFAkr6/FWO53LISgexzOuCj+kpcHYLpBVGeb2ZRdyqrTX36EzcrC5j/IRieRgEEU1oM
ieXs17hc33xK66xEooYZZLzgYr7AyhnW6yiotphc3GDXNqNmGQ9yVibjukHG3uDs6caIPhDGr0Yu
ySLZLNeEZzgUNfeAshW0ScveHbBP0CD/wWj6eCoXSt3dnM0nK1o5giMLcCrQy5aU9sJ2lGnLyEjw
Gl5E4BnQfERe4ZvkqtqPuk8FEOl3/vw0IlfxEKc3v1qLKKIdGwO+gphGhd+Ap1IYeZNbcztIRg2l
HhIpVHxLwTd1F8EgDN4f0O/onpLKOWisxRu0FA48BZRyMyODilrgh7OecTR6rXtGbhBZM5ptV9D5
yfIh+1g+wSUISjMHuJYZ7EdEKsCkzyzGGyvR/bRM0jV8VpSndqQ38JHTyEj4I00RqQ5JNvYV1d41
YfyVZ/93wsWiC8qqHWbyoG9Oo8CWf/UuZXXg77YQ5BPSp5ONseG+LmNfNcxRPbtEOIEiDPeQsjWI
ZG2EDhveOWr49MHWL4X93HqM6NaAFwr3+Ay0KNWVAUMkg+NH34eGCtYgC1KbU12LzxOIVnIhrmAQ
bJM0WwdPKt6N9WUBsImGaROwFkZeoSRQYVI5UjRB8OPEmq0kyFJcBq87OD+40bpDrUHYpSMazmHo
FRgWxPGYKb9xIjvuw1zxefl1KkjUs2iUERB31fHOmpnXD/jSOAvXx6a8wZKzcea/oGR36u3Hb3Kj
oo8jZHUvo2AVNmM1lT9kxAI1yTp58MFPeXsbXpbwwTv6IGQAZ/OokFJIvJ4YsETDOZRSvzlSehN0
QyscTCoh+AbqEYwysKyQXeunjw7wgBbLLVarRp9unPvEBKpkLWVqBk4MsdV4l/gihxEJRsOLPITI
DjjlBwJyskbJ8FjZ2plxEjeWBZOrCxcJ6AS52ApNw6kLsBrH6yksRrUF0azMyleNP2n0i6LiYDfB
mA2hc6QUa5Kl81sh3+a1vyZyWSfd5IKbaLED500/OLmpjE2+GkVGtYB5mx8taeKD8/FmO0QP2YkR
fln6KA9ahbwPmJ1/WJuLb04wW5Gb9zKeo7lIKVbF6X7TrGZRXPziynDrMG3Ymrmk4hVaGtkfKkZC
1MNnZdXtqxFFC7GCwFt6KeWXWullwLOB3PiWNw7cUR+lUFPgwI0ydsGZwRL4bsQTjsFVJvuTXr56
dLorhBeYTAsOxfQmHjct1jhXPF4mB3nhIaRGPsrfx3pUGslqmiKI3O6RAzV2vk44Hs7pYssGchUj
iER9zVr0H0RhU8LfPGYy1yA7RJnqWMlfa4SVAc8rFdWuG/1dFugDh7Wur6ykHc3DdiT2qzNFx6AE
GXsTk0u4TDUgkkYzVUuNT6Sy7fH8JnMmJDmF9l8+EvE+dLgNkul71Jh2qtV6CxG5qrR83aZjL3QG
mCSpkvSYGmbwUFihjHHqBT0+vs/Ht+9/gnhI9M108+pixEbE8bCaobeVS1g8nIyfKtDYV4ZMm/Al
R+fcnQQoEukuiE8pSDqFOvMFrXTD33GRZ/rB27xMTq1xeBz5W5Bjy7tiqASs4pM/5IXuunBIbXFI
faFp09n2TdRXakhauvBgC5/zkW2Kc3N94xfah+Is0ctM1k+f7/f7ZYSALgns7x5LtBcATPDV0u2o
pwjZ4g182NmuraSYmjI/gN4wi+K/FGkgsvcwIpr37RE8snia9RuxUz8C2ytFm+hlqFFruIuKD+K8
/rUxI2QuWmW9+eUz5+YbSokdO/ByhMzEBJoVdPbnIFjvF18/h539AtR5ZqBm8dl2LxIjeiJJSUxg
/5pKX28rctwgwqOraizE9rsMr5meajxSVwMzlKm1VePSZcrHPWcbDGKvWf84QGtgdAfdZAEBFBxP
z/X6alkJGQ+Sn7VArWY3rnRwoLhtoemaORyOtjuZnTJHyfIgjkKjX4vNLllCKd2qijrIxmtXIOEU
h7MUw3VdWPblf2OtP0bUqcUAJ1zZruf6JALZkKj9AbM5orsfIOK+pPBCr+zNAxoEixZdIy/WtQAE
3QZ0ilvqm7ij74nJMCcLX5FjX/Pp0q3EWhqtEJks08Ydm7ui36A3ghSfPTe4AKNbyK8X8zq1qXZZ
rvhgjQAhtKp3Q2fXuoCdqjhrWBz0HvywN7NqVbYcM1EWSvnhS6nEoS6xJPu6x6IJmF+z1x41LCF7
q5A6eg++omg8Fo8NRAGyi8cSJB02W7PL4ohUuITrmEse5ivXk9k6PC/ijDNFMBxqv3LyyC1K1pyX
hSgtNrvwrrtzrKU0rCpMoDSy3K8UfrGbl8/iAhR4SOEMEw4bq8r9vjVtTt3+7VL7V7WPs8GCHwt9
K2WWhpR9QhUTZHN3C8TWnNgP9CU5LqXRSujtnqz3cRJt1y2kN50951mwdL7GAxMAc9TsW+jGoUdw
RjyjzO/nF3unCsRaS+sJ5A/kz4IzBoQuPw3gctBy7gKohgrh1jD5iqPS1wGZKQPao7NvwLr1zryI
nQVCQFfXPyu3Rva04bChMI4XQ/ZpJ98diBXg1TMWZ/FBUJRezpWnAB5BNiRt8e8QGoMJ6WjS7QCA
q3b7z2nAOpF3jIuhg4ZlE5Lc9Lo66p83cYRy3XMcPmIeJrJkXAOt9otoh9UaakRWAQ388wKNLrTw
+ZgCO4mK0q7lfzxaWWIh9CCyFvcWbu3jdwJPC6POofmmMzg6kUycAs5yMt/QHjH0QYsjLf1q1rlA
7H6aB4Ccl3579C/CcyFqAPY89pSiEGJjHQih/bfREt6Xl3de4R4/HWLluVj980EKTi98jvHPQOo5
Y4+04PR9jgzUdOfwEeEKovHbuVWSHTyDSO+DzzBIOU7TMQ5Ex4ZNF3EzcPvoN0ULnwcDM5Hd2OEe
hQ1L6wOV53kM4TaPhp+MHEJM5Z0LtJSYEWm2L5uEVnFFQPEXjbd2V6k+g2xadAZevFtlbHr9/4h/
xsDdBpb6Wjz0YJRvtq+amovsukeZTgoT8bdGQFhXnWD3kgeGPAZkltNBQ+uGyfC2c2klwj8gY0pW
gxqBIqewAxfJKuxsdszvSzuVNCmojuEt93N7ADv07pxv0brzh2JDIUhxxAbpC6S7in1hQxD1ZCG0
qYTxz0kcAy8mzPlBfezHn0tNSHWjygF1ca5ETLLRpOo2DRVQilyqOAqjmO1LWmPbHtqCCGg1j/Wj
z6vEcR9sUOC16PwFvnstR4Bcg6M2olOxasz5OJwhTEj4C1GG/ds0Maywhrv/uitMdpJuRJ1tFO31
Fu9Zw6n81BkrlmMwgR+pxeKTCcsm3MRtAtt5kWpVwoNjB0YBWDveijk3hc3+QBa0ELQpWILBGvsx
hWoxH9VVnJqZ3OzrxaURITH1M+addydOGMv/jFLph18yVL+nGF8bXgv+Ln0qaVS+7ooGiHyfmp7+
Nu4VxrOm8OG78zRaQG74nYwicSBf6hyQKSux0f+fcepsmU3k9zkUzwpywnenOSxGmB3JuDq/SGIO
NtzUUbO+S8hvZ7nS6QvFFLC5EjNu3saSUdAT3DQSbiCaopt1s97a5OlYFP0tp1KaNW4Svt3/3WPr
+2ShnuiTyolNbpOf/aFi5tiLmXPZ7O5cW3U1VZ9PQ2wHGHErc+xpwTt010sMcyBGTfsvNY1Zbvtg
FYw5Xs+wxcISKumbiYirfRRgkRgKdx/vV30GrEARYkUrza302Fc226MURR96n4bFrolKq2N1aQea
zWHiGfPMss141FeRQYUOIZ5We6neyWko/fyt6v7SGM3TT5qytMzN5l1fgpPsvIUpUKWFP6c7p4b/
2aeLjIX/GWRYAdcx8QKNqu0zV4pwxkDLe1rW1P51fKZnQA044f/XxJdA1JFYBOcco1uKptHevMEo
FYl9M7GwpaND3ANquOaJKAzLHwJqRPbnG17awsIZGr7L1pPlQdHx+D9Ak3Yn+hI5LZ8sW7+z5FsG
j8Lu0xBl9Icx9pf5nObum4qdU2gBGakruGZT99Ye4spI313/ezoEtmjl0P/jDJjnOQpXy9EjBUNR
BP6Q8Uki5dU6oWgMlGv4SFFWnSoC9ZaFBKfneruIReRodxde28irUX7fEnc+UJ8xGnhW9vhQRFtO
3UBNpOw1b4GTT1wBbVbjIF2rM2pAemCm8yVdJd0Skj0fx73nUi2iK8Tr7ZsbCuG8tiA8lM5s66e8
LinnJ6hoy8S145QvKIbCZLh28Evj/e2DIdguzdZ49BPqDJs9t2QJRDXZOgdAlOhYx/6g3OeJVmhh
r+UCkqTAr9lXFC9NzBv9eYdQLwHN28G1CZgbZ3gq/K71ia3bYBhgDsv6V4ux9JZ+l36qvqX3Vwrf
Q/fV5MNWljOyzhU1d3EyeB51ows1Ah8PWiBuaQDdBXCJ61Ll47emxHczF9aKLe6BDUIkUwKj7Huf
anjjV5bQF4A7LtzPA/6VHEL3Hp6vfG7RUkatgbJHF8g22J6h+At4XQRL7dtx/3ZUxrtXspMeakSy
LSaS+qIbbYFJPLRagWwiPKMIby3PmQT6fXAkJRzPWBvtcOnl2pLL2VRiTd4cuxJ/mMrJ+krQEh2K
BVpH8lC7rPClkPLIOydBs07l11nX/RjX71N/Xr9x3IN5er5dpeMdoqSsOh51vL67FY3QC2b1lxA0
qRt2+3HYu7mvvG/EHNkBkdIzOXq/QXOzxj+a5RL1somMmbGeMa55EAnz2CtQB/QkajkkaOwC8Vin
MsAyP7NYdbPjB9+cSLXwMXOYF0faCbQM72VZKd08E7UTCRGDHK0wOq9SyiIJcPWajKXnr4ioDGxm
u1Q0RbFnpCAG7qxGRP2xn2Vokc3d3hsWTRAXEjHcMXTfhPyufYLVrJd7du8sQXovreRwB4pRAN/D
oObEPjJICTm1jXSUfqvOlGLPjeAx9SupJTWRkfPlzk+Ae3E3bHfItHiYqyI9nFHwKiEUvs1sD4up
scsmav1UsdRZF3h+YqYDNOBtq5CYMLmdfPrQxjRVUHl6w+4W58dx/MFW8pDtTSZpiQC+TrpFPsju
UzM0nMASkQBL2XmiTx9YMCEjs+GkdV4DVn+fK2YsVH0riwbocwdo4QJTGInF2rcLJs7pbzC86X6H
8IoYl1RaQcPqdl6Db152yJVUV5Hb7RxT4j4cuXsKx9jg6sXYSCqRSohexo8Xx1QtJLYk68mLmJXi
Vty0s0sAJpHQkhW1NaAqAous89sv33OorF51UjQiY3TrueOhUkzlHYv6TTWgdmq/WKrGw+1AAPKU
NB+O+EuDL3sxbWoqXVG+PnM5LpMseAkDbJRdMsxvh9lE8XOtzRZ/9C0YOnKjDnijTOcOdCcrPD2F
LagvS7dRl2QPuZv90nwW8MmFK2cPnxcfOZU+FSRdzr8oXf4u/6dBrAxKJl8fKRpw4v8NPHL9ecj1
aBcEbT/ysXM+Q4ornUHFZ5SjtQplvUdm032cYBwebZxfaUyPD+XrHQdY1ejMfOP4qKCrNk7qbetl
wfp+nW7AyZOglEhfEGbetUlGoa7rWBBcplhfy2m6oblR3Tbze9St3+Q/yyb1/GipBIn/rrs375+Q
PXxyPAHrg2X1mGyJncxdPSUxnp1gU0zO1mXKVjfUJv2PLEf0bIr3hfg39deDV5nsLDyMxWLSF7aS
nAtAzLrzk2AE8Fy7EPD3bNTA6pUxEzUPMLesZbQkYnq0fXT9KLVy+kWKZpDj9NiC8i+hNzmtZ6y0
BZ/fMspirrQFJDoVcJLEBrz6/ftjXFIsjY5/fo/iRYgaH8H+bBewcVUfGjJBDuXcEhKRdcTN+6+B
Ku+VQXE9MkNYfpMMr+fVYOLHYU24uiquWHzTbyQfVkciv0tRmIgpUr8EBnLSvlE5RZbJ42k2yykX
yBNpdpSJD3Iaj89aEH+L3CSqXIriBQ23fhrM0H1Pu+7ZtXTBE4wxm/Tj2EyCayg5n+1kOV0+5n39
Q6RyXnGlvwV1pWrDhREkxNWUb608DWSnBUrtaZ8NLHZKh4RUOGjeisz5HyFsygr/r+KTtYVMtO8Q
umjkGjRrq6pDp1TeA5/vLkmRAKZmFZFZ1fAEYkPSIvD7r9W1w8H8HDRB1n1tDeT+XCH00ACov3v/
Pu0KNZc3LhZs0Iyn4ck9lUDFQx7gWCU6oty9jFi3/g++JaRCvhrcv+49+1UZ8NY4V7yrNqBuik87
S0r7mF3UDYzo+F5A5he9kU2MIGlh6RXJSXvSzYCXrZw00FJWpm4WyCiaD9ks10UkQ9ooOcWexa7w
Zjioa2c+y/oqDdiKYDITBcg+YcAypN8ov5iz/fwcGrG5DJRVkC9o/sSsv7r7rtswM81diUohY89c
bjkq59SKedPjF37HXtjWatyZQWyc0etMQgYod9AJfdT67hkSO2QOHxekqPsphM8YGE//4iqjzekx
Jix9oPNW3jHqXAajwbNBKTdE4x03x8JuAx0sOujJggavGWV1XwrSwXyZ0eDDPCy23QV0BPhVLC+o
RvnYwXfuQEs6BKeVTlnTVDiBNbRQlA0GQyxAhl9Jn+Gw+98UnARkrNsxbQQbPO+vlfDEcABOC6Lq
7zOwppFAfXDRXjeuZGAdVzYUDjU1vsRKS7+47QlCI8cZTPXPHIDGCN5CTBXh115TXJtujVCluZ0m
byhWFhZO8wr5bIFQ+XT+dKwWRgqBqRBPYE6RKHUrJWFWCkVeAgH3G8oGsf+RsqTdICBfpkeXqR7j
z3s+j7+d+haMC3d9+eP3v9xLwFFLLRD0Eo6s2rwk3lrkNZEpEmqAkqbGQdLLIKPQEMKIyGZ9/3gP
AtaB4nNPcmaqAz2lhIedKlS7+AbKXTje3AgMEdoKDfYws6ZfnGx40NzA151o083sP4DjXk4QXtuM
VTDCqNga//1z6k0XY6bdS/8gkQuGV/GkImQpS+QNL3xspQjXKQf/XLRDJGk4nMxxxhThpiyFicja
6mKHdfxV3wNu1uwsxgd43Dcl2OIc/jTxqAfXvQUwRtZGS65p3NzIm6UGZcqxArL/iJE3KDw3lkcw
1ZFNYztcwoSw0v3ZoNJqt/rA30wCtO0tzJ9MPXdYFX2VYbqjhODqHjDrSWuJQendAJeZWE1PQWJ8
hBajdSHxSMRTEZPS/QfVdHVdp3w5DI1xsI8FddhCiWlpt1WGn1pab64IK3dHlJcVk7hcmlPAUI5i
t2SPs5fCTVbpOgg5jT26zbPI5Ny8kOou6NYe4gfFPGq+ORd+A4VKZNRZi+569pQ6ynFX/66V9Gjj
kIzYVQy5dj/ioFntMzzP5s1VlNc5kcmNiUNk1MLYo5i7PMI4LovU3t7WmF79Cif+uD0OBZGfnS0B
a+L5sXekWbvie4FZz3EVd/ciUkDmCDQ2JSLGkpxdAO76De5WA5EWgAiJrNabQ4Gq7kZJaszx2Rxv
HnqB+agy572zvmU3mqNSSGv/TLDqCQO3DfMlfDSboT9RV5tmDCmSHkY+27a+IOamfWBOWdVOjPCr
i3aRgnaRgrsuTl+MGcCm77lF+juGWKCczjM07IaLvRlLGSwN3KA6zHXtaho9D5EAz0enikhKQXoq
S+D9ltCzd/GV+v3RcswXybqWPUBpPHVrPjHhd8i8pQfk15sq3tJ9Mkw9Zs+QQblRgduzP76pdU8V
lL5oUUJtmnA205IGjMKDZ/bZX35NXJapUyw01KABAK+BnATjz15kJQV1wfzj3Yt08HIDsAW0z0Y+
X/RRyvs/35+auaNm38ugJp/ezj89qD6/HxBXJbd/fz1w6D6pMS//MGSkUVW8zoaXLqoxsH+pIDn3
oGLfVOgq1tY9xox7rTHpCJCTe1SlIl8adg0lcihsapZXXIZHBypRfczmoGk8xQeiak+Kx1wJmWlM
yJKXg05v4UCAjgfy1C6YMEtIsNMAsAuQUran9BidKTk9xwuXo9fI48F/kgohLUh9SGerommcLfCk
o1AtpWExDtgPmOTNEoUtPRbdtjBJVp0L4eJ7buDDJeGES4znonXIXN6dU5lFUeBWPQogMMfrndO9
1+ySQq9X2KFAUyIx5pO4nanoTkorc4ELdcQbLYSz6itlz4qIaAcI/YPHyCizYpzq6NEfCB42uixn
WopzU5GKVC7WxMDbfY/UHme2/BnqEU7sBzi0mjbwZCNr7fIJ/zY8n5Qv37KPMyZ5OBAjoqAd46PN
hAJbc5vaAxSoySfUUsHRdBvhnW9vr2F4C06VaONfaGOPVSg4OPsa+aXnMGED1T9vL+AynHlVcFbX
vYp4cijuvaeHZX6j6mInb7TvHfVZo5CKJH3jeMcb2VR2we6x+DAzYx1DzT4iamSNx5FUCJea5d6l
XlDSaHspEzN3KkppA6qZ8vM5F8NZb6wz5Ae5h+DPco0LwI7U5CS02h26DQ4Rj1W/tZh6p8Nc5tgu
vkGLOicvOjB0t5jz4OFdyMJxK+yA+2bTNAykpfrXNaX7Qi4aJozp3ZW/TwxJvmjPNAmT8SMc0nj8
EAz8ddkh3w0isRJLFaQvBU0TmFES5hC66x3kUdolTaGsdI9/sx4FP5756J+mdlPCpJpNboc12ctc
YPE/PRiAPizRgwnjGTGW2+g6KbdN2IBfQLG47rOOrxByTN0uzsO5qxTgjSL3qF7spVNtBikQHTBl
hOhKdVL0+IzEYfxUxFEzi0Xc4RqVTqYkda+l2ZKddR16YEmIlTmKWNjBreuZcwMpeQ73j/qU18Pw
C46s9VtpIM5GXis9nI2mFdk2v6/uElRy7FKFQcW8HAsh4fUWxLWKMJWFqL9q0VcpVVJLuEuiLTiY
WT82qBUAvhDTEq93+8TF3iofx1dsFJaPOhemvUfc/VbUkajIw1PHZhqqNA/JoeFB58fm9wcJ2OUj
DK99jPOdksVGsbKPn6yBHyhd6FgE4Q5WakFgdASDNPtBLqZgeHtF8K8fdLf5OjSUOjOSQCp4+Fz7
AKGYrcDCZLD+jO46xkys0H2zJ1087nUfZXMjjzmKNlW36Qev0+QTS6tpUm4L3sKSTKDyMATiUAIR
u0iSpibfc2o4XJvL/ClMZYKHlr4SVFhqb/Bkzh5nrq5pHuZe3duewXZDtbhbpG9iMxjClqv8xUG5
NK+BXmdXoO4IFaCR/x6JATf7cMD+2Cq3pTjW6Hsml+HA+DXNqmd8ENH2NA96Tzqhwv+SSCno5y0t
WyipE4sIIKkEeN+OW2Q00dkFiMHdtiKsgz1ZBvOaDCyzG20GRUgI4kOiuXArA9giN+s2mlKfbSO8
/W3UmQxA7583M9QRGsDAjBdK1HwR6liRDFYiZw8aVO05gxdxzU8aMF4czPlLJEaxgqvEaDh5duXi
AZEsd3EgvDAx5Lq7kS+YsjsJhlXd6l/d7yguzcx8N6tkBO7HTPmvXJ59Dpv5HbPB/pTLciahn5a/
0yjSzgBoiu6LZSC/vJlivv0z9enoFOV+JAqYUaS2F4CBnbFAHZFM3NtxjSfpZzP2DN5Pay55hdL1
QDVcE+Se6sID2r/e/MIL11IiCNOzYjrla4fShakMVPmCKTTWsmf9XU5s6KvxCdlagfkH9y+iQPyV
L6edTrHChPTpbRAgh24SyzqQ1jdRqNvvb0o418kmNYHIZMXOGusdLKk62BZ6pOjX3vocBFqVFumS
30vK5JrAlvGHq5t7i5B2to5mQWLOFvgASL9d+ZXQ9GhuNZ7nGZi9VJqMpSVFOTB53O2WlKZODfGF
L6SW+vKeFsbtAMBKKsnAolk2pTNyikSVxesO4Hd19KJsBOk+vV7Om4IkQXMGScUm7X7Thk9nhDsg
4BnDwE3V1k4NAd+SZPLTMCNRs84xHTINwUmruo9rdtlQWHvSu8m0Uml5VxpJNoboeunn7FB6d9bO
cwg5LxId5mRRjgoaEqWBihj30c8/5Bfw8mA/NEi64Hb3zt33UCukHhI7nwMUuJlSvFgS+IPwtsHw
Ojdx6SmAkfsq1oVpwZDTlgjaXF19+6u4qXykhwUGPjg67bB2E9THqLkDZXC9OkKhQdo0VesK3fIn
TIDayTXJfc462WQZT0DPx2sLdl6uc24LPN6n8xuVJjlZ/D7X9SOisHdwV++gr9m992mjSLwsdZB1
u+o2vtoYuOVjuL+xp3K1Z/887RZIp7bY/VMuwdEzVnnC/ZqYEpqbHVL7078j51EV8RmEHECKvJ2q
iluEVRjmMnM9qoloXdsZnQV3aU57yXpVULSSS0McGk+5ZWKeqUgr5I/C2lbNm0+rl8yir6gd3c80
D/jHJNxYzL/aRWfJUUvq2LjsyJ4Po0FYNkkVfWzm+mf8903UuILUuApxerXAwR6PXvXoZkx/zxfT
MdVgXiZLGQKtzCEio6Pbj7sRSaA8fEVJ2+QhY+xMlmqylGv+BjwxvRsopuYdETG9FORNK1epnbGp
3v53KOer5pp0/DvNh7wYDh2dqyovPMM6c/n0NR0SNPLoMUGszoycrIhoUXZfsXdO1Ngc+Vxtj58f
a86VhjBRBh57mOQRF6GFhDNxKiK8sdM9B8FdYMLSq53VYXxMme/PlBE/sw41KmUjdP1dI3xEiSGR
qyxtyge5m7AHB0j2264HrbH8l4W4fwbqHXLU9/cL1iL2Pn9PwG/F+qYPcu/9ivHgRpZH0lBvP3H5
9JQgkt+5f16xPa2+uVNuhsf9iFhJueKXxCCfw0RNNDN1uOgarf1HIlPMsuHUwMFyBsjWzzV7ARLS
c/ZKeAr8zcyrTtLsZaukTSxemCsKxV05GpjaPovx6uNmT6UlyxgVypzKvylIVqH5gDTBRhZnK/kW
adz2aAITopobG9tAzH52RUOYHJMfh86kEJ5FKgwL3Qh8ofbN/Ss6ZD+eUyzwq0W3cAm0BHwrW2WT
mqPKyqCY9UNmiRN7ln8ebE+Ml96TnWt4WPju6fyOb/v05EUsUo/vhn1xGmNJW9xMThBN05SkFZvz
ejv2I7UuY1+wv1c3BQboUNnhn5sPQ8Upk0HUXW6sxSatGqaMBDbBpaX7KCq0s8yNxnXDzI/jwjKn
MgC1z5uu17o5TIHH37ZhT1Wd2YwUhMdxuE6AI0FnaR2WNOUuJENnSlijL+4mPSSc83+PZdLYh+w1
9TMwnBjQGjfDM/TBEMnFl9JVa/rj0raPuB1NmxY6OTw/VTwFXg06W+xbdCTeAwNXcv9Cu64aIfs7
xs/oStCieY2EWie+jv3D4jWQcGp7Amib7PtjtaY25xOJeYdbtGfiLjjm4GzTzA1rr2qdJHZVC5A2
zauzXG0VWu8X8zQIN/Qyjm0Ze0Pn674kQTMFu7/GGYlqs9lGSuaYvpUJVUfUpX1XTHZvx8F2eTUA
yKjmiqwfWmJ+FuhvaovNnuhoFJV0y3KkVoSZmFskVHh2L3uvmpzBuxApuwS8UE2I5iLtWg5o0Nr8
fYv/SvzTK0m5zJRbAAzB89G5ug+OlKvy7IdQIDQWvmOx3AeegmzD7svD/ySjTMtk8afYqQ4627HC
jXq3uDA1u3JP/GmCGxRZ2mz2965dR8h8PWLO3kvvIfyTl5rwTIUg5MJwyGSkiboVWjJ0EuIijO4c
gE6D6Ad6qpj+A+ciw8+9QwzzdI0ISBfhn0E0Dgg35DuW6aBI+yZtCkfWcOgIagXIa7z1iykXDAQb
5D/M/k/RnuniG/bha9p8APpnhan3rWjWDdsYWp7Ilu9HCyFEzlS78YNOot5/9xd2vSuF/qvNZ7Yq
XfrAZyyOxpqWUMBSjNI83jkIS3dmD95sAfkkysdWUnXRz9v8frtvFOEOltWTSbQF1GyIGV4Ll9LG
415NkDpAAt4RfZfFxw3U6r13lh9Xi+i5/wq0Lh2cJjgR6k9w2TtXrifYuyGnd4EmDEttv7GwYN2g
FD4B4vSZxDTDRlRQP8TUoNVLZe3Qfj0YufVZkdn6CZF+xATVssMmKSeI9gLixyxrExCPEwjEs5UJ
CpsNJf1Su/81ZmW+XhQnKU8e1Avesys2G6FIL7UmdyU2BCZAN2Tb/5/WPU+CkO6UkxA85WXxSmpM
H5eSYmyoRCydIUrx6aAE5t/etzdyhwwRrX3iKtmO+P/7uxaHbrpYRbEUkwp88+r6eIoxXfE+7zAM
hMLxW/PSjD6qyf9cBD9U4QSwn7F8ryhT4voOdcwA1xW3IQirjeUa031f6styEzCnxdZhVjHdf1M8
3eKrBOmpTh8NqOYgv64tiA7uJyF5ZeX8BIcHV/Xhv7jQvIsw7K+umuNS1MT00o0YDzEvWljTL1zN
QADzx6VQeWW+nv0JrgB1QFi+461cXlS9SeJ86E8/dcXDBOAatf9WZdrt1ctFXbmwEEQGoi4Twhei
jZKDShnCgfM50N7RR6clzeDMCHaGbgsKeDrMPR4GMo+V2IOcOwDCv5jjyIiRVa7Gr+NcK29h7M+O
bHxZqBOkuoKTt/jp1Cf6agheoG3Mn7DXzkRqEBMUsxXrGwtmfVLbi8Urna4nheisGzdI7m+3NE/U
duk7Pp6sCmXQ14PRr/up35bX5lfTSzBrm1hvHiCpnGK3hE+HgozCqqo3IK4LBprq5X12jy3L24jv
q8nWxtRE1wFFC63Dl9oUu7imlfwZJaOigIxP6Lvc50/YTdJGDkeDnsxZbZK+cH3OE/UCAaQ+CVHw
NVmlbDoev2hUYnK+++EtyNOq36j0jBuQD7+7BFlZYEGACNmXJp3InqgVArOHuTk6y3xsmN9z+phn
XdJH9YwDjhPKk0nJ0jGYUUSf46uTkhATQujOk/gD2q+epK0+nf8QolV8hwpDzYPr45fAV60n59gL
PRDfK/MHdGhjpmGkAI+9G7FCaxlI8iNXf2cUKQVBJp48hsJBShNjBPtX+yy8UK/x3WLxOMi4nM0Y
onmc7uurLPymhsrUIxsWkaTJm3MrjmHRMoMzKnwEODg1Cpm5EqK/YqW52tBVXcJcTuyta9khmbP+
Zd3APzk4AzON6nfEBnwOCWzAe7nnT6y31hOpfdydxALSii+JwEngkTwYjkoPSmxWWpceH0X26DOx
4AOuJDweS3YtbARM/MIiramR3aJi5mauJSBzi6UKhNwJf9uxpxc0Q6HPUbLSLrRoWLJtRubnq3zR
UcWwLGI0dVKa4Mzp5VS+LKFzaBN/tz4C1queUcVplVouFQPqZZzJZeg3QHIud2qp11/VMwiQk0OC
vzVlbGdVKs3lFZ4Iwd5QvtDJpx/x2W2ssFYxxiADoIrwyDnIZcR31z+93uHoiqeI/F7XX6KhtHto
p4PVtNI955Ce6Jq/VuJk/WdsaG4l5kR0/MzKVA1nTQmtQ0ec7MRwKnHkdXKtJn1eSiTaJpOueKPZ
AEiwAdhMStqcsXwdV7GzWCDFHG0ocSwO8FwB58eGash7m4y7ypTodNfdFi6bkDLvNkmrTo6zfDXs
HFEzEgBl0NETLwsTGmkryY6cWbvpm63hyXzrFEjKRPDR8DSSNV70jpgxEqe8BjQJdOwL/s3MGmTJ
+MZ1qWU905qjRbtKH+4nF/3iO/bl2JVriCZcoXX4v8JYq/TvOearvi8x4Xa0c5Ro0wtJIOYJM92D
08D1yfKyjevvF7anU/F8w1yE0AScSDK19xhKOoV+qnojOVEg46P5gkrFiNoS8MpUWMNIgy6zwP6z
QMMOA7HRtawZeo0Q4GadwE4irYI6Ft8ojaJNMP/qSbBSxKz+b3/VlrBnzfxaBmMCQUGkthwcowoZ
KcN+SJ7O35ugEFbsVZ3/v+7dQayueMU/4sCRbhEAqOpLtVQ94j8pQFk5Mx1ZMK29DhbMNNZq4dp9
IvOB6aU4Rzplb1vZiJTmld1Fb21qWs5XDMNIziKV0bH0zb2PVAxEHFrwWdS1S/7RoaoM4nyjhWyY
fTzKUqAj6WXLC8Dmkira7WrE5sFq9Mnbn8uqr88VvXpDBIIVmX5F89cWSm9Plkz4jgk6a1PyGr9x
fEunNgQHwfGbqikfm358DrBZYO4Rf5gs6vyG+gJkbKRGjXN0aWB8EMJC8TsrE2U0nCcQ03rd0uNZ
LjTzZgUt+T+uLlxw8tebxb3AuudHnpaAZVm4aQU7Cf71sstEYNLtBN88usIGmZJcOuH7HudiRh+F
txAXE5dtT3ngkuvs9jblAyZxVcZsD6YEi2BGU4rthajXQO3IiWAmKSCWzjBQlBMutOxhEq588Y5/
ZRf3wv1Qh88MhtSLe9DogKjX5h5IZej1wZ/tMVJF6RjHt2N/fmJpjlPmpgu6HP7jYwf0PAsaAkqa
GiEQ5BztTZfT0AGOqgW0FGgDvWsTKMv7HKl8r26MirjimR4ukIpwNwIHXqKvkLcrUnpFlloxpjwl
yQu9IeMQsELIPa99CmeYQh3X+SvIhcWCAqlPKMavuuKodu3VCnEiGytEohMGShGpelxhorfueiUq
LUEFmzIZ/LLMWFSW022uj1FuphvLJjJ7wEG2h7K896viZnHf3WL4qCeXyiforW3HSOxEp2JxAUiI
Dnj2Mt7Olf/GU/N2f7VntJFeVOplfS7OZ2W51urj61p7dbFr+nB1/vYjzwo9CO80YVAnFfsMR+yE
VcpJOEfLZBjzCCjgaVaQVi3P5dwyTkRplfpGeI9gfNdp8p3gNUO1g9JFwoSbpezyN6EMKRp1DSpI
kPPSJvCrsegiSVT65RdZrnwvV+NpXkNdy2/9a/U+1HylTB7x6b1zV45x2LzxZEARGBHvxu2EpVuh
hVD03DbpS8qliynPFInsEfXw+H4nHkcUu4vGXHfukyT0nMcaEAkV4G8saHthjnKuKn/Ips9xsh60
gA6HqNN3ztFCEk/E1pLaJb2cdkTWQZH2sS0vJhZh3CrB5mzwLf7YMJryzX0rmtdQySX3bo2tPaEM
DyBgkr2F++up4cYYui7dE8hftGLeNMDsiCvuQDVFuT4NYU2e2ueluuM2QFK+hyABoeuVoDK+ss3N
3wPWjWOUpdjtZCBXCaqa+BH2xVnyTsyARJz0D2oOsfFxr7mBzqFEW+LnJSzXBrIKp9akwdZMLykH
ZLKU7mFING7gRBVG2t9aILP8d396j3TUVIOArGDx0aHqoB2N28JCDr7eZPv0irU64s7VVp5t25oX
UGeU66FsBuUiNXVC35lp2q3D94DBlvUwAharYhHf+l+Cohq0A5G0pvVrID7srwPqs6xDBWLJubuX
HAMbFcn0K81bYPQRMYqhVuLB/lC+r8haEUBXbZO+BszFsir1XqSIGzAVS6RYNfL/0xUFrUtUlCXk
w3KqgfVRjWtfgL/LTIwEnGYr3BxxUklpnM2NIeRmvIlZl5IJN7HlP2eW6GRP41inuAMVm2nHZvWG
WqcXuwzSCT6mvIIrcl+ZXHGfs90k7ItYZVg0vufLDGErt4QnYCzpWM4d6fMQzEZRpP1LwA90Meyv
YJ9hX189AlYul4DvNDZExf3UffL8chogmRfqP0yW/KzeXsSivpOMUyK/SNmaRVE6uZuSuhF4LGv+
cbdBzktwF07fr4HYX78YLmyioGbRJ5uAiG4K/ej9uXNJ3JjoReanuOE5x+MHWPZwmjHDHE2rghG4
MNFgO+b9OQ+L2Es+FzCttYZbcKAWwJ27l4wOGHNDuZhbQOS+AaY25w6h0HVJH2xJxMoAekThE/CM
DN+YG9fC3MQSww0KwGF9fIC4G36zPMy2m0/rUAdSkSmCzio6bhNvveh+Eh9pEq4/2Zpsp3HoZiqn
8uumJzXfzqUn03YhAPnswyvsI8SqWvhJ28w1a5jqXvHwgJ+8CI09R4gaT7lxj1279w/3km4UZoDv
w5W8ZmVE4EX7IJt+WrdVt9w8rGluBmApvsuSYskkPajG3oQvWBGoLsL9ToO2edAN0iLECkoxy987
qMD26o8enEKsKOY4oULapTRLS+VuneUR7FbWkc++n3P+14+it4xRVSPcp7qYkd/LJ1k4aM/xCjNy
52LWskOhgy6XiSLjbY9rVY/Geibc0CeRwGOMfXS0n7vS6zy4KbSOGFsfd1h0ujy7RYhUjFfU+yJC
XGZwsRGL4EntmohCh3TqE8F5GyYau3PCF1hNf2YhT004uDD9rZBbHeqBCPtSnCQ6RnEhVN6C4W/8
s+W3ck0bdpiTq2k9Dme1w/kPqK7xOu06ymORD6o3U3jNoxFj/aJkeOHKMiPK8hL6xhTscB89z5X/
jQB+EsI3j35SPptcZhc0BTthsAG1Q20eNBOpcELpXyutsVS6Joeucjl/daqXANWlT0OH/tpPfsvq
C8XVcNlDCdqnwYdbXllt44agRk4R4t81sUggHYdBUP70aafwivdrEM71VeKnK3A+0gUNNGU/Cnle
L4ErDRjeJG0KezQZjzkqGa/i5qGdkUdu5y6qIqa9mmfgHnnl1Kh2o23C1F4lCosGdt37HCu1/yd6
fpg8JrDdFUDcqGnpDignOjJtWEDea7yI3BuWpjjwwMceZDiYBjaPBQ1SPuPoLLtSGtxA5HxIQUal
m+ZUyVk1D00HdD3cu4RHHlBuybyy7hb8wrps8KPkMzGaL+DeRfU0SdNl3mctCxvKIi/5KqcuGoY1
9l9vJKJYNXCJv1v47Kcth1QgjsheT7T6F1wxyJu/h8A7gYCCuSNoy558YoMwkQv8WpqYrTzHTkAp
skodviPAeiENJZqk9N75C2ybfJar9r3VSD8zx9rbhLdfN+dzlGEHOMizgf8SVsiS2iIrRo0LAlMO
8Qn/cdbs9ut5SkfhilqZ4o0uP1Kwtg1yDLSWd1UQe/XdXGqgezfLyXazkgXHW6tx2anI4r2p0fO/
hr/wttrFpiThQIpXCBqa+47Hcy3qa7mAHwNi/C9bOtT7dNzifsqYL4lNRDcWs9H1N75MFYolRq2j
3U9eBTCC4nJBWN/CVRz/zMrtzYt7vjXbE07blJV8bArDBTb0jXJM5uuBvZE3TfX4NOmr4lZe79uj
tXASWHxH28ENFXy2hHpZfllrjddUgol7TeQb6gPlqclKIQkbuKSHdTWK/g4GdvB19NWgk+70mjRw
qea2gvVVymSmBoU+P8yxOOsA/FPmbocrfqOHOSk4W/+s5HrjyEQ844pDIZZyd1ekgO0J+PyRwYa/
Rf6vQvIzqMVPBmD+Vu6+Ix4TjRpDIwM2u3P9f5bBQM8IFP8E12qan77wnGrMD2zr9SAARQCsiJkC
KmuKgGt2Y9SEYLlfAx84vXPepdF+/VRnCNA88EfKbA9Mo7ybFxOkFM+OWsBnDJ0X/7+4xI2IscbQ
CFuGFRSvJwp3G1xzDfkL4d8HXk8+xV1obEnpzVXpop2MvI1eWsvtwqWZ2vP+eLPQhcH4vgfmwM9Y
Q99NB7nUo+ehnSyfkTH6NKVY3jXHSJLkmH6CJiHyzeNLOGShoY2oHRhhM7LyKTZzebWekhmV1Dra
Dhp9b+iYZBYkvpGiKvN/NmpHOk5bQrGJUQNNCL742SobqwCRTcLA262EHTEUvCpmAL7ln+HxvefH
FBD/bgIESH0SQS4Di3WK0UVeYsRIcDER/wQMW4P+lnTJLt7tFmdqf2xWsDmpL++4oI++ap6CJVhB
gboBjWK1SSyUHQnvG1M7GRmLH6OTShsbp6OORmZCilix8Nwq4gs2KymM7G3VP07LBesE30qz3Qh4
OWzo9jzxSVtgJ09xDTBsBo8IzmxWPyhhJnW27WvuUsr/DrJw63q2cqa0YkbHSDKLWbI06KyMW6nR
ZznCmcEnai0FP5/Zjsz+JNRaGIQDZbqn07MngDpoloI5dBWJ+/r6LoSZNIY3B1e6kQ57Y97lB63e
Uxm2T8mkJu1j4b+yJ44F8uqBFRPgP3tYdlBYiCRNbI3q1e1xaiF3Ob4eQ7N8m701EhXtVTDlagVD
UxAQ32XReMQhtruOjUh8Zl6tr9jh4aojyK5mCqC6C4V51QDvG4X3WfFHPtOs6NzEjkNgOWiLvLh3
tlfFTzEGtGg37UEgfbRftoidmoCgUj1X1NR3rBdQleU5M04wX+E6i8qaGYOcKTxFQq1QgkPdFKbu
vkY1fkYE4ZOfHCKpjxiRb0u1BiGrTnn9mw2FbKjI3EAwYMG7J3ZmzjcCYzTLqZaWasd/jFw0YYyz
b7LNKhZi7SX65MsBjk5yWzJnWpWubA2QH1R76w6YvtmqlJAsy4nQbyRipLyQeyqfrh5vuEsXVOn9
nU6oSBDNIiKeuQCGJjy5g3iBfAVQeufk5QBZemgBIJg3LBO1ZJyL9d+VR0Ume3x4jMAeYitfzuDX
ybA1yX2Gf3W55I0a9EY2yWtahuxnRB7HTO7eM36eIkb19UQRIz7KiyZxB3ikBXiBfogF5rqnvr6G
KUJffeDt130oxUfy8oxUGbYVOSR8/+mkqZBJvEG1H3H3SFsT5cwrzwoVZkUi8PIiDlyZ8hWmwGlL
u82c06Svj4luSc3fQBPU1WkbDMzMNQnxRfZwT8S7FLxt3XZHBgWJC8n39bHlzClSMF77S9AW+2d3
RyxlDpkPDfaAteCjZmSlMzA/9ImIJfgbZZKi6xkERzaPSuZL6Tyq6CEziH30y7qwvTKiHh4CPM9i
of3u/aNoT+swAhe09/cLyH6hmBM1jirbNv1xF0afmvOHTkkz6+Ze2Kbrvc8G0H1rEzARJW2cK51E
YNSbZL4Z2MoPh30EMwOvOdTTAVGI+2BD1m451ke6t0M/Bt0elqfoEGh1YFfSGDS1fc78kvIh0DB6
S2ixpL/Zk6wNA7+91uygdGNe5auP5wDbSEGF4x2KOa5domV8tl1TJKgZrfmPmtxF5ExjVa04ujIP
lBqRQduYbg+1Cfu4cI1Iaxm8GppCU+JRqcKLjIh1zcTGYl2ofyCN/CoJgTxUb0/axINayrmrwRAD
ua4NDoHrF5MVP21ST+VSzsRZMcv35Vx+0NS79kSb7t+UQ2tumwDrI4mY9HnK/loHPhBKYSNdlDBk
1hHR79ar5SlkhT4WeQrbPBoLdMaF8DJlfAEWY1uEm6S3iLxhY2AWWWEm7ZGqMF8AFPCR+76flYXV
DUL8bO6rSsXy+L+3WvnVSKGBqQVqOquvvmGoTm/K7BYLc/nbcglcck5tmZnqe4I7kWLB09Xq+YPq
tcj0ZqnES1I4KKQNRp2nGjxecaGBKoFIz8pel0ja/7Q5uICJ4gKsJ4+RwHNWIVOu7YStL6dGii1W
10zbBaqGXtApk8jSzk5tdum6YWgHxm899rHmWR1DtqRb21NOCMy1m0LBLEKMBo/1I8NFjjh5aNYe
A2ASLgaydq+cSPjmkV4o9LpvrRRpySHVZFAeSYwq/Zg1CUSHaOvAOXPvJkut/izI0laECCoV+N+1
t1dgQOieSwwLg49CG6IsSssQubed/CP9IdSPZ5g1N6PWf/mj6HU88m+JeWpL+BvmCL+DqVFRyAi9
w5xxmjxF+rfMyO3VzW+8NDyeQIWgrXrUYL8f3gCP++dl+jej21w9/vPDhPSnZdWHMQYE5zB3oo+R
g8ShTZ4L+4HVVYZy/Dd0DFTUAKCujdq5ggljdump/f6vg6BR5JtQ8ZWX3p6LQB42Fjwjk7knFNvK
X9Svmm7vq3L/8asaP6kvQf2w9ohtQ/1eoKbomEcZxixpVPxgzflxmwr+gcmaj3Za7Aor2KZTg+wc
288sbkoSj+HGw2a+uzIthsomewd0FUCbZMb0Z+vodO0DX8XQYuPYKwhmGpWCS5TpSwGf6UGnzAEZ
OSIfhbGDNiuVATGq/BJ8LIA+xbpf/oQzgOdSvF7kdK41ZpudiMOjSm7uhYCX1D8xN0dzZfAIDZIv
sHbKePzgR9MqdDBXCPPQ0JgZoWLROf/hvHuXXoAFOhuRM2q93/vxSW1AOpro++tGBaoyQDd8dE4D
OXk6+cEJZVvuJM7grNpPOGP/LDp1kEkTdNKvOmZANbEC8oL7jYlqMaLz7Ru97yVKkuCuDWIpvMWS
GlZ/ijaRjjqHu5mVbCOjYuAqny7aprzutqu7PU6a/JPaUtNKtOK7DqmS0IxN2kyJNYW3Olf3RDfC
SYT+vi/648n80EWpos11ni+MLu2beBdCZegESqfQhjm73RQoOXDIVfGfnHTXax2AI6P6u9wDimQu
RkE9MqLdjZ1FB9qbCBEKQyt+Mv6miMgylvZFqMKIMOIYgUg/5jokPRz/kubU0ysiOLdga2ByRbx5
7fC4DxVj92rlMy94u/QYYs2B4PEru0chkAD5oN64SIbmvBKO+qIwnkAM95MpaN2OTfL60yd7JXPB
XdCkvMif7xleJ5fyw6dun69gCFkS51XLZgIZLdOt3paSXk7O+11k+tD15riiAqli7ShV19PclN/9
0pbZjeu82OQ8GU1qluZZShDDfZIIUYbCmpcvfhLQWEp2YU0/hkFmPWXwfTcnt1yAKdo10w5pVw2B
lFo/RKkart1TvEjbz+rdHgGssapYTRmvAO54V0BQyJDKJ7kTrMigxNazFJL6M+EtEQFCdn0nye8L
bSMCvVONdxJf8PE68dskw49Alva6/r1Euos40ERam9SffPkJhtLyikzvSqNuiZuZA2Kk+Od5K5ZG
9FOh38m+CdSR9QdLHIZL/sd+KelPQvpYPr1aQzp9tdUG+c1Js7hMsGLRkvrKunOZkJVkibfqedo5
UxfjJt9E01iEi6qdItmddkS0e9/0GHsiTawKP4fs4LhnnHFKOqYP/lBEfyk9/wFe9GKbKzmFEPnL
eJKzvxkp1+cI4EPAE0vfEvK6oD+NAVFP2sEHiDiQpLf2sUwjvxkXRL/zbqWxQyCCLkN2YuLmwNZK
O5Ybz1vA3omnMbWYhVF+uhVXkMWTYnogI7voJ2+sgeUAFsIgcA63aJbean3pKtOF63ufGl5siTRQ
8YkX4c4nxLNDCRtDEJ/s9svWVo3OPDBUbC/qwz4gvBrDaJhMY+WsdLhe1Zn7VN5weASjSiUjdmV5
PCBv19g1muXreGCT3ZJfwGF0OCBvLNmZae72vkpdlK6gR3OF8nwb/Zr80iwhglC4sA3X5KYxdfYR
6S50uhC3SkH1V1l/egRIX+sBxMH5UobnEiodEHoWrTIgeOh8BQ/0gGDSYE6Exhz+x8E63ssN9+Da
QbIvZjuTCcUI9+NmNi9DljhYrBEJTOzjdXb/yXCaQtOfWqlI0Ap+AYFVtpH5/4ijP3n2IUf4+wXk
8vsa5BR1aIEAYoxBUmIQkWaf7vw5Ku50VcAmSPU7ZLg2FK1isrUkWJon+qDXL7+/Oh3oMovgPs+3
C46YrbLTDuQa7QcVssRwWJ7MTxaXaphxRN2Lhyk+oxp+z6iDdcdWO+BziN4o1lE19ddBY3pVIGF0
fxrOSsY8XOhVFdn4VszduzkSePfvkvKVr9ESM7Zqtye4bhLLC6zLg4bImL8NRE6jYeAYI/cqmidR
wDEy2XHWq8o15IkjvE4LEKb6OCWb9tvFALToy6L95AI6eHIVXjT3M53PMU6e/QA6ezIrTh2qVokz
3c3iF51dlgFbRIyimvr195m2IyusRQv23Lz/dXF5ndlZZdl8xtZsPQZ6M81kQILEvt8RqliebMT4
cjSXqceHIzRs/OItLtmGw74t/L4zyb+v5kf3rr1EmGKEYdDw56Sfx//OKl0anI2+LOOtm1nsSH0C
FQQymQc8bsX0UEe8x3Bg72gmtAPrzJB9+uBPpauIOWGrKIs+AiGfRgy/pKkDW6JmCwKdzuW/+VYz
DxPAp4c8swzKakiC3OXGQ+p6OyDEx18T4Rs5wZ+FlrP60EZ9MNg5dCZS3bVnOFJf0NxSTFmTUnrY
sieXCI+nAKjwDV4KCb2OWXUIdfF9MKbGFWTMG0zAWCLzdoxJY3y+HyJv605nNoLJ9SCjyUamUaRR
LNz/ylc/toGgyo67U6wv2So6lbNil8Fj58KDQUxErA2Y6mMbyeQSj0/yN9YBsy4jQBHyO/mcP663
yjEmHS6iKllD9spJmoU33Qw7eLs0kXgCk2geBSeDn1VRcRxBn8AblB7UzuqpX+8V01wrDFiXU/sK
hyzL03uapJKnGUe8QDsuT1RJgOzAUnWnKQd15U8yLI0esibSH0i9WFz+ev3cFmqAEOuZCZ+nNYLP
ah4stFkxgU8iIZuXBZqENmydVO1YYEeISvGCtDFYXC0OgdZS7CZFPkp2I3dnH+RWH/udPMi4S1EU
9j64VCFOMN4lPzOfZNOX2UGmDiffUrWxxMlcLRqDn+EKMHmJfoFNoGfzh57QGWA3nDhNTy5irBzg
LcvGGVY6Kh7mJ0JsfZpIkXS3ZfUygnOj0Tb1jM9PYUzT7tx/UGNHL0SXaw7C6vaHyfRY6Dmzq7e2
8zKGtpD/ZBPH4/pxk+9gxYxu0V869JOtCIlCZF1+fHYcHx1qFqCJgHeycz4pIN9CZXMFwE4Bd/ny
g2cH5Fev5EYwsyQ8cvcKsnW1gmEQb9hRets8uWeuYDmRuFWAdhQLLl5TVjNLJmSVoiFTh/BQH7Fh
IjQ9fbea1zX7HW8rDd3VLKdKjLu4ozGOAqS8a97m97cbdt7ngRWrsS+v48ffx7LYcqdYsRj4CIBF
FXaoUBRtbhpe/X6buyTx/YoVHepx5bFrwtNFMs3tjnUwDs1di42OhRfazUhULSUotrDcKN+u14Om
VeYTTt5U6bwyvsnKI4dgHhiITzoHZTCPQHGMpDWdOrD9I9woZRJxgsr2+i5jOfMbDF04JQ/FiZ5U
4qNAjNZd7X9GKiWDzVuJakA3LgiozvY8F+UfmpjEIwAPuTmR+3Pm5t3y4pR9Ji+XeaTAcwOtHj2r
yKz8olQFlKs1pU0SVMdNGJGglHpapZ6bhyBb6Lu+gn+vtsBThGWs4bMAoSrVlR4qlWjYBAC7PUUW
D3gLj6L4GGzGlOz0i93t4md1cHJyzjqZVlfD3nEDCy1W9pOX1TUKLDfYn+7lWhW67geleAxcR1Cp
aoeTmn4+D+bDpTZSoRA6kNooURG+NdouY97feyYuPNdJcb9LnAxhvU7YMM0KU5hqkMANcuq1z21v
VKWc5tgpjLgjBOY89KDxImE+QIxdlZnP1FMACzCKCciSeqIv1eZTto5gccoOVfNIYEam1WTQ07ew
KgrLGPEFQTNLlR9mAeKWF20p0LYuHWhhmMi784+lk1Z38nUM2NREtSZjTVeX0tXdLYhiPisN4VSy
jxkbIFNYcqYBa8cDI4UnoYNXo6BrPB7c4cjsQjNSWv8QYNqUkuGMjZ/ybaGYGT7i6AwyEz20GD9h
Na3geWI7B544IIBWUKNUzg6GTRNnmdQtEaKk+9DEiguoBC3MqPHYBHfWCOBa/HJ3sNmJojNeDdoD
Oaebmg6eWuwf2/HFY6V0roAzdVboEmaNFI8M4d91LK0jMh2LGUqqET0WkSxS49e0UL0SRa+iGbsX
WvCYe9a9s4GwrrD8VsXBfaNWhakmJleLgNJTMK7yVUC0q6MJT6hnmK3MqLSmYq7LLHCFXKiDMOHM
32wOa84K61r34P2iGnYlien+7CvVdkPmne0qBf6YRlW+xU4h7MmhYYwX4Xrz5IZE2S/EnvtA9FIZ
dx2+knLQmh2cj312xOU89TEqr1j4blJQUi0Wj4paIKfdbxSawuMnKxG/bnfMgwKR0Lsafw2R1yT7
kVnxJB9HRAYKE6sAZoxSbNqB75Rmj7Jtr1POwesU5iWP5akEnHNWm8objYFM0tK60ta/pyvrwqwx
bBKjX71qW0tvP6TRIAD8tMdqgYmuOD/2EQN2wInp4fZNE6PNzv7rpWvg4uyeEiajdROzNgt/rpjs
jIn4kxh2lSZyOF8Tx2EHA8FBhGcar39nrpSYoctNxPw1246CLZEhW7FOhjnu59col1zzUM0PaITF
KSEZCIDbgt9btB7SsgQPN+wIolL0NQjbiCVFpJhe0kME/e5UWDBz1R6aIYEEwMbrNaVbtX6896Jx
YRYtIzao/Mplu8mp7fQyrYslMo8fbEZSv8XroF7R2O9D+OnD9/xMaOXd2CCRABZ26du7+cIk1E1R
35yDL/SgL2qstX+s4Mmi2P52OMawGFE60G/1074F04oDYET8VeORCKT4U5ut2f0idfL6pbDIl9mG
2PYvUk/6DPyzWLZPUPdEWuaChVUgIr5fVFOEpu8ss7eMBYGL0LBeE2gOlxq5tWmKqPcLQ5xM8rtG
6S5vqutjIOWvE7tPK9CL7Kfyk3ZolRxyFjDK10uGGM1yutwQH73qWKr8Elw45V6PoFrTnVvNURmE
nSPA1+zcbzPpjSHE1NfdbPFUymAGgMljtGWVMoXPw/OoSM6h07rHiQD/W4zHJxQRnXw5GTKrkhqy
BzWrqfk0S6heosZ2Ey9nzBuDrVJayyY6w7/b1/82xLNgW7tKisgVm6B8Dg8cIt9BYXpM7/N7IxXf
W9ASPZNusGOSOX0v1OsXcekRJy/OGqJ39i/2QrAZEQ8Sf9TroLJMZS85yPPMVFOBFjdGMPP1DDsF
ZJHMfw2rnZhA5lHptlDNiXpn6LcJ9I0cGyC5zHmiqnGlP5Yl2lskvkmZCzU8+TZE8Z5j1tr5qdlB
qMG83oKXfUayb7EH58sWHyTNLvKKDu175O/ictc7Oxaad8YZO/IVX8Vj0f0KV3Ji91QhmupwwQw9
oHbrV5vT2xEvqLdGzrw81x1qZqJWWs8MM/ELPs+49SYd5vggMeEZsXZ3SAduRfvnSb9gvVLhIJjz
sNqO2ftzNpoJsHccjG6BVpeUovuKiWzOR2u/kYLqCsJ8nb5OU3zmZUftylP1L7cmf0N+73J/13NM
B0/XsigMq6nEPocM4Y7DY7mp5dfuXU44bPlrXCN/+eGiIPcOfgZV1yTg9rd8bn3G76iHx2dltSKC
cB+bFeYhYSRC+AQ+Ua6cLOuCF//4RfP4VS65cega713kNMXbstz/ewGgCCRfdF2z8LqNVNyBx+EI
F4geb3qs/ZA5hOuu5fTv3frBZPGBdqXsG+sgygV3L2oGiQroXSNuwZ4WBiHKUqR1O7ImDvvW1/QB
Wi9qvUl9scC+2HJ95qbsYiCRHn60CPUBPpTH3Oy0f2UoVreDJvqd40mPy1cxETvwcGonB5Oc/Tda
PwbqtQs27GYa9O2quc8XFEe7m9wXMlnTHYWFt7Gs8Rb8L/do4WsrQWaSypWmxEIXcGAstzZF85We
jF0oq5+AonbM732OJSTO2E14WBoa897Q1DABT8yJJb3wmumMZz7zi0JNZjl63AXjecrVtuXytakI
QVpIORTF58wNMUiJZ6WN9LklN69fhdOCI3AmAJpaDo93wfsXq2j4g4Mp7LIdp/MQpqUfH4a5MTPC
hfua/GSb9g/sBxfmnvhbKqjMNbauVa5bs+KJ3BrKi5CDxS4Y36l0S5EIQIB3e4UgQjyeZ7lYmfsJ
DmKJSM3ofu6vUeEv9axyKw29JaVSBKi0oJco3Ay/aQM3dOFTc0T1P155grqP5bbU6j8ubTcU137T
Q50renYC8vN4FzI9UMVEIXcBFnjIqoSvgd6euWHYUoef0epSPrXtEqfDooNQ1xj/wzkG6DZBZ7Br
pigEl3evzyfY0pFTMXvvco7ujIM6m/tLqMlNIvrl7lbkSz8pFFT2ssJmy5F+4HtASyyX9P5Dl2kV
/AM9ltQSpx4A9sLCoP4OuEU+1Ym2WWZaDIDu4GFvM2sKi2mBO/7Kc1w9JJFNu4KaAu0PPrMdSk/n
DTM7YgptXR5qvG5V5P9rWmFGpHdBFLreJml5R4696iRvH1PgLJYvoJ2pwlMIuIAIwfESqiRinSuA
jWuzTl1b6zvcHhs16Pj+PZPrEWXq8QV5wT5n7dTxJ1iCseZmyLDcDvGgEhGgYjOGsPqvBFDRIYXk
jxIpR0MefH78wXrIwEHtw3GWpzVRLIFDby+lo6M4BBXyPvNV+uRIde07VA0SVkT2mE3n9YD6MjUo
kZg6s50r/JODan+vRfvqFxuTwqJOYShysWgAOCzXzTO0t3FZwOaTGqg+aPYbBUz+OJT7ULFDj6lH
16fDDYTMGg8GH7H899v+w2DpCH2hgk02qGnqYZ7pYBZdso5tPz/Z4ic8X63sDBdLYH+c1e5STww6
zJNUPQRgVU/nSid5IwwiHw7GXpJCgjI/Ss6aVr7dTnOvUPWCZbLNBaxjRl+TUnODnCcwmd3XHFUO
Pe1H4Ah/wEUOa5GKR4/mavVvDh2g8t9QXtLY6AkUls7n/AIo8a/dRnBcyI6MUQS0zwbNcdQlPsq0
5nAtc0Iq494v8BvZm4r1LLFbeuAslDhF3HZ+IrfM74AjTQE/XOgqda6sqfDiYnfhdcP1QuCitTJ4
P9ZxEPIBZ5Tc1IkY2yooaoeJPGCxf4bWGPi54G7W5Yd9o3oTPULqbg1bjZfFEAyPpLQvdMBpVKzl
2JkHB9ywENxDS3WEUt0DRtZX6fwYIp2Q8MpiSvv9kKCD42ME7njoLdsxmXA4qPwz9saJjEy8tg7Q
OmXeUzHHlXSsaFmjLbxz12QQs2omEruB2CU5/QHTcFs6c3A2uY+j7gvSLWtAQMIHXQL1aMhE1LXV
OO4N/Pft5nrBomESwkKK0b0eo1MHzih8tHUOZyqGJNqz+4t8pridm7VRmSACvDoTGzzZM/CQSj6i
GKRns1PQ05x+zwjYJ3EKmaswaIVR86eS9a3NOWnkSJdkgkkOEiuJS18w7axdSwgDLfIVvpm7FHdz
ueGcIZOi7OmDDn+F4tP9gI0uABVkVagZoQ094Gs4f63bRCawN2CQQCGN8wiM+6yHD/SWAgLFLC6W
7J6g4poEF/5vIK1EGs3o9nGjLDtE1gvs0CZb9/P2qQcIN71E4nEea2e/bNjWjAF+MB+SQmWbyrgZ
um1MWjVcKsKoC0vrn3YPVqCo/HcHqTsYR17aC5ms6nZsxKlSDjiLCr9mHVPqn/Bh/W2dJKimbsCv
QjcqBB2dPmHpMZwhGQHEWCEBJn2oZ2Y3I+nOtdNfTbRWy0GxnmcypkByFJrMlq//m91pXI6Tltsv
xDXPgsLGLGTN/8FZVFVICZNOyspeLJrMjvYL3o6B61EkwoZhsNVIrxS+CIwtz9tOBOpSxLrO+lzI
kQSNghno/xE/xD8uf+F4zhDh9qGo1b9UsdK0KGRpXjbX2/pm5hlcVIM+J5qmJPEFn+xoaDwpNUyq
oFd02NAtN6zYGWxvD0+Q5yiPVcbWpYqT2A1D3gVJy1ylB7jRYy7H+v+AF2cF6i5J4CH1fv2lcJfi
KBTtLrTSNoW9HEq5Gykpf9hmcXvx82Bb7Tfe8FfPY0ygJj+izPCYNEiqmcMD3I8aPdtlbeYehtxd
mi3ZcSeeiJNhb5mliENT2hX8ocm3vTdr5jGFVj41V92YhsVlz7YAeFHUhEL7+sAXsA728gY5IB9a
q6DcHz5deOznWbWl/19BakI85/vufK3f/BHC2F/kuYzEJTK9R4rAvQNUPW3V6ag7UES9y0fToCzG
uini7bRmE5IwVbHH7EZiEiJULH8Jo6MEtGVyd75n9Ns2+4GiUXSg9qVp+NPV441hwdiw00ombSL/
gY6PPQOT2rbmlEBD/3+/OIqJNAP5/NRIHRacKfUU9QL9k3WKd10ZXvus4V4j0+NWkvx2d0Pxt+vz
H11KifLCYoEBq5cG+N/14DzAnhb+g1KRv9VNEIgZw68ajZWM3CC3j996wrz6+vGByZCV7GwOPWSk
YaDHZlx50v9oaWn2N+BNgI1inFFY1SYMMr7JXxXeUrzdJFx4FTKnJgcBql1UBdLn3JjPtpustFR5
AYvlKvoUBsIVQ9EV091byKplfH0ecq8f4IzsSk3gdwxebAgKnt/mRWZsImw1o/9UjOH76ilxYehG
M087WzO9K/qQjRPgwI8ki3rAlsLMDPje0f54Q/VLzedb0ggS+Z0DsBXH1ZUQdvFs3VgPvm7TDK9Z
tEjUii6GBCXduV7R9SyoxGaA/WVILZVVij8jZlkFL2l7+hFnaI1ysXIU7382pKYTN7gxMrOo/RDf
udtCJvonsIsVFemfqR0s8OKwPxY6deQH0o5/kh/+Sm1UzXbnsY2dbo+9RL7qu9vS5wrlSWi2rr9L
SC/SrZg/VsAccu5qbiwgll6cAwpw2++z7yu7Qg3yiSI1w0jSdHXj0TgWiU4Zoz7Qh7yzUMm81FAz
UBb6U61AimO5kTjlYNCZJtsQ+5FsTSqA8Pc4AlphvG+40KCczoX0UUzxVrJUX1JvH//Y4OwPiWAv
PBcbxRhheoHVYvajbrld5srMxA8obOeXCulPFhU3a2iDuBLlrYyw+04G1T1OcaL7n2FAIIR+/Q4D
+2u5ci5j3XPFjEEynNxs72wxVgxbX6EXadX/pGazQ/AE6xLHcEiizMd3OWeW9A5wSvIFrVl3nPaM
k97rag/J8ZuHAJNrk77VeFzQbCINyOzX+YogQ1ho+B2JXBJjfigPEyrDcuzOFTmacYj13gFbrywm
3s81jGp57LB6cJHMZJHOvN00tAyblyl73RkTGrg0mojF2HaxRuQTPGX6ZPbsHsIOqBy8NLru1Zkn
/nLr6nugwI7to7pzyPUN1SQzsY5UKS6Q9jlNe7mQclG6ZKak+hGpd4+V6yspjkj+1kiCZc1Q0613
t0z36oq8G4Sidsco3TNt9kb8zfkmfbclEm3WLa/ikvoF5n/SMyPdHlULfqd9aniuNnKFknMxQ4Tk
Gvm3i20gIzD5keRem/kTqKmMfcZxsbYokMafPgvdB2yMTQowQay71EXjDqLDWMACxJJnnEvDK+EJ
Abh/KYrFNi2ge3WRGgvHtyGRyjc+peac6Xm3ii/aa4DRfpVtCREJuRRdGChgGOFfp5P+23YKl0DV
bOvn9UxyI4YSqPmEB5ZhvIuXHUozYEZqNIHva0XbxMjKQarNmE1MVMIWe8tUn6DIjEtlieyr1bCh
9tx+I87X8G35XojJI/ImQbXkwKiLQ9sym9FQtq7md/tTh2meYOdBWuQmWfhHB2tAgFUk3U5RhAag
IwUa/N6yoN30xgsrbNYKsF6wQPcWUr4t+e6JuAzi6CoFZ/YWZNVUB9lI1D7HJI08CM4wfsM1KA6l
9gmhDTIoutPcKQYAPgx7boAu9a8hE8fJKx2JXbXMSOoLswlvQD9U9t5JwIWvP9Wav1AGsrLGQLR0
b6WOd0nrmiyaeug0GjSJIG5vfsy3l44lhpFWT0NC+L6Zk74pbeYYcC3NE32PtXcQ0HTNhLKZ8JWq
TBdn82fghqxyTEQyyYsZAZvtiImexiESQ/hv1xy+EM55uBSzZMdiXxXYXpZ+HDJMv+sh+lDr70X/
XMNe3Y35VvZNEW170BJ4Sj853Q1QMD/NBnK9UBv2zo1ymONUl0K51LuXMMEc00hmZA50sbG9EtqJ
2NVaNnbe7W1sFDgMch7ExiPWyAJVvb5lpd5g93p+dZIbkYE0idwwwnJ8y9+WgL3Jt2RDQVHSFc90
YyGMLddz0wIxsRVeRjwcRGzXiPKMp3630ByC8aFews2ldb9JETQf2YAcN11dEFTZgJpFddTE8FmP
S9AEZSdMik2Xx0PkhM0QS2e/k2DvXXVfGPhNIVrKx4waA/5bBptcr/O+rG+vWlvE0CXhOEgqevJJ
IZsW2rE+hZLyqDDb46z+DKCfd0R6rdz9pXn7tO2SVgNJVgjB6szxGjSR796AEIML7uwlX1xNEXD+
uoswRzNG9LsiURq+Kbgl1HiU/Wpib/3Ngiuc4LJws1GIYDOw+35lVJ/6SuXMEHcsRv4100btVRGg
h03K56kCWHbnSiPR98VyuPZuxiu18vX5w6l+sPxp3IhxqdASBqZhcydpW0FC5t5AlY0aNkjrG4SP
EocoiTFsM+vd+FF0FNFXCAd2GM87jq6Pc02n5TdnC7EM6mcsbql/ngCddUNPigvJgynCGFIxC6Vq
qPXyru9xuJ1j9IISbt9u3ygIE4dEKHs6hXLaUyQBlO9IO5zkFOK44gOkPq38xgvJkKBrO8707X2M
2qSD1sqOKB+mI9iSFkY6u/guBocLce9yRptftOEO5yeFhJt4oXirYISHXBPsJ/XpSR5H8T13ihBw
QNiGan6ytsqF5P0TeqPMGon2uDEnhmsYeRRLWErlzQ3/CuzZ0528Z7/ejGRlym6pLdsuQEZSDCum
tbQ1p+LCuLwCvgfe6u0bvQXVbz0+KK4NNVYtpxGYZ2zGeM7AmFgTbjZa9kA7T+ZGNZ8gdDZsp/de
TozUCrehj7zjcclpTTc9rXaw7iJ5JTgEwDe/wDEPSp3D/zo+3uLGlr4hiEo20k/Cg8czJDksvRff
iU4+4zK2qU18CONSEU/23i65QRapBBLONzWgvWLrj7auZQ5AR0yf5bZztw72a63hqXqB3a7NEXyt
Iil1/LBBF0jObK6lxbBKyl+vNIRKerkJ4R7q3S6brgES06UkBj1Gdp3ODfB1uyY3If5gLxRe1MSq
kcepHGvcaS8w+D6/A8zEBCE5pvWM8PsY92PwbwMPsfO/UebBaMGCoe/85JjVk2AfxTvKxwP/GlzS
L3HjJ5hqk9RYcpCf4Uov0IrOfGHHbOyZSlDO5/ZhYc/EKdnmjvC+jdHQ0LUrzjVVoJPXejgalDSo
OvfvFVG9wRyMD4NtfPs1cNmBUnwMhDLpE0d6LBdTJefn1kv37vuOj2XKCwk5EiBS7vDvriu3QgGs
k37NK8DzzrQ/hQO2TUh2BdebGScEHmUU//cHIoGwMdIBW3E2j5pyYVTObTt8L6jawBCieH1CuzzL
qfjtdgV8OVgaiLpRmQkZkpFpAK8xZa7EBgPvi518M4jnc3k/5PGpqt7uCTYQwOpb2VvZQmieHxzD
M1HlFy4jjYYOy6vPXXWT/O0VRBGbIJBxs4lu5FEnekxG31mwaomOS76wICsADXJhj7pfEJZUSwcj
tnx7UFbJxU4ctBPpug7iqEAE17H15XNkO01F4ebQvVVqc7SFdazu9GD3HWaVTmMNMHCEZcGsx0On
DwKmyZGNUQto4ZTjDWlYTZTymmYqOMAPkccyygVZwUXcvIUIEjzHm4zQk9bz/sVdWpGuYsXtCa6t
ePYejXFdfr9C9gFINP2Kt2qQA/UEaZ8IocT1RlGyGsq0cCGCdFqjuA0IGtkMHp9EeQguYRugsUGS
I+OIsXVKK1z15jGApZNVYI1GEhs2BGmetetC9c0LPWzICAmEb+05pX/siW80x9Zu6WDmaEoM7HLL
GbJ/31eThCimW4ObbFHjcSMxoXop8Q0aHgkAG6HJ5D5LbzYndVBC1uTEkYhgP68b4yZv7nPyTYa1
lhgJmvccKFg4MNHiB+wfAMjGQr0JRRGgXnByFnx/UTRS0YeeHlgfRYDGzJdXhdW3gJjZn4od2tPF
M5C1oRuhX8nVhnABY7/cRbXkeBnkX/XqPb9QMcX2Xivt7WwDhRy0ql4t1J3jWLQAPiktLQpPZa2s
FT3AEdJ4UN7ZB4u6kvlJEG6nToueFWjTPBZKvz0uoKLokYejCXpyHCLRAR10Ao5wqO6swAgrXVSk
ZsQL0JYXPuhl0DxS5tX1IL/AFX1FfzaEtgIqh1Gna9JgcbfF93R0nbJpqNsTEYnQXgxBMoxMfaxX
22xuDdjvNiiV6KJ4qyswZFrRLFLiv3tXJ0SH9juanMGnEC8TIZBnxCP44e8w23hzCrVRnj6VL+c4
L+sQlhjecBBk9aLeSNQ7pRZ0HWvevxcO6frvlYFioVOiVbzlx8vfLkoZhR8hXxa1BucUz+59QO9P
unQynna1ZR1GDwAq0wObFlGcdUphZ1TDp+fXG6Q/yMDjJR7XPZZPlzcSUCP/tMV6xm3jSvXSP21L
YnikbAhTiQ6Cw/ed3Uenzcww+/Gsgul2RYuJVSq76ErudnJGgfGqkOo8VZUBm6KuSE3DXtsZJEUt
Uk6SGQao1eG77dcCxgouw1LYKJGDUUhPw+WpiXlua3RS6TnA2oOBcjVpTEPa8N4ExjCzp7SEibdW
MhNKLfKVWlWF2qAECsLQx0jyoOOfgP4syooPJvP5TvO802JMywj1IWVzi4tRSWMoJtI3hx+h38cp
Y4XSlEWFypJ2P2PWMQZXO7gaQVA439EQL0PPmenxbZwNdguCChVJoT0Lp+JE/Y+MS+UXL6mtyNgt
z9YPoMd0CebfOUDB+5zfYNydjA84ZJMoc3GXOy3lsyUnND+KN3c4Ro2vmYcIhoXlOc5M7Imc0A6J
F2J8Mv7U7/7R/RZl8nOtmdq9pcuo+cbXjMMvoBYX9lXmW8MlCRhoHwCfssNDta9GRIMacNSXuFjm
Uo5FXg/efTkSPWVwldrkXKmLseMNcQ95oCQ2R+dXHgPhBaMWuy0P08M2u2GUpihaWkrkNXGXNxYm
oDXoxxwvwYorN6a59SZCXp8UtpnM9eHqRo2RtezcrO2EFPBXWJRyUNCHsqnsw/1bIYLSWKumwtmi
oO8JMtyV2IajhyUujoDu/+e8iBAzrG8I88cK9PE7MnQI4xi4MjkT6uOyxVtAqNosbT12zLmTkvxa
oeDPGKbaiqwH8hw0BWeY9KcarmOLGs0BGDkHTog1MJtDEkcUlj12GqqOQC0YSPRT+DaKVUU5TQxR
w801mhz37ojeaq3VbOHDW3TQE4DFsmgS/ZIIDHrH+RIUSkXeK7UgP9xeMDB3UEQQGvPVWx62Qg3A
wI0VycJ6Wt4e9t1/8NG65YsenjGkgHPCroLYXyyqq9mN8ewqs7EhShODkYSorldJvFl0LufEV00k
AGJ+yLOXkU9fIr5S3DMCwJbFoWGnz6MksSxFpmIxTXe8B47tFz/WjR+Lzwgb/0IRclmBWO0JkEiC
WQIgLgO+DAzNHrh2eykD1pptmrgJ0jAgnuD6tRv2m25IyCIR/EVGQ96xqJaRqZT9fQubSgtjtDjL
ogYSRXSKO+5FECsoVL+WSVy9IGlE/8iXES9onwZJ/jWzf+7pRJUCAV/WBPxzBPXD5gPCx647ygoI
0geeEDhn679PEx9+Gvn3PtkVJBFaRDLe4OHNQxeNte414zPjhBEvPRRA38gPpSavPkPpgVmjefB0
U+iBDlBGXCa/o5CuhSJd/MAClH7r+lRfnEAwixcjQ0TrfkSi74MWIgk8ae3oCR7T1FcXfKOcVsOE
eelAcqdrLBBwhvRf+WUWE2HCVl+IJCEVWiB/X/Q3iw91hKQVyUXKUYfNPrvUeSr+6zw7+i9KwlO9
VGTIMRAcch95k5AtM0juy6lqRk7EqDayP4kcA21DdjWe7dsuCVqMZ9Mnll3iPBOGcsHPLDoHfr8Z
/riHk0EN9KLFaRQFWdhQ0Xj9c0opMxOStu/yUilgdRi6WekP/u8QvFVMfssxaZU9n0kLfBrZf9Sa
QRYYYabR0extWTtSJ0QBqBKI4klbbLAxMvUyD3BoOdTU4AucgjclDCDnCX0yP+yqsNe+31hUyHmQ
3EtbGumZoUES5fCeIuX7+GaoPGuTgKTTFm/5JodMa7f0FL7XOixh6RUmr9YUR1oWYyVAnOp5WS1h
Xe/P2TwWbJmEA2jqBUVgPruMXFe99BvLVtIk2n8dMgmwyvizGLYMCoL+JC91Hfsdfzwd8svTZPZi
0mvicMTNEe2IffERr2HnLYJQrXYvQJWhQ4w2efF4a/h7syarwTMAxdltiLlC0BNMFHrV4znyZgWT
jqwnrTnPnLiXNt8RRGLZBeJy+GaiysIsPxc5SwFa73UX60ZviOGRvOzy/xjUvoSCKO3eJBb4aFh9
wteXctyVmPbDtL60zBtJwBVb92DVt8i+CtH0KAThVzxUR82RG8rUVqqH20AqrMAzoFN1SQzPvEnt
TbaPO9zEgIHnUF6BQWgMt269aDaEEsU20L7vj5VG4RCl1lwJeegYnHZPMRVlLgQNG1pzXFkUAqFk
l5LI1NB7Vi2oxwHKY53Pa8iLLZMOl2IBmeODRqeb70eFk/3yp8fRrnSqV05EBH6i+U7P7F14GHID
cAHxRuTUYx3M5r6mAAqals6Kj8nt5o1LflmTHQCqzYJht5nrza06H0BSxMIW5Dx3f3lsTBmQK1Vy
d6HZtfI+dGxPNMMm3pkxjvyP9ASh8aD32MMspRefqpcI4hlYe7jQubR/lPb54WOD0+7k6pat2k9O
prSdbmeHGjcOfVT5io90NnaMCO7qc4CF+tf5MYd0nraRMv6tejoBYNDy/lzhpoMAKbG6lR+kjADf
odZQK15svV+FBKuK7owB0oGDjjf/77jAEjhSldeGWQyyPPiSMnujXgE/mpPiq4H15OSYEhp/FZ+h
zqiKQDXM1qLnUg4osdrnEG/1uQbad5u6v9SnHeLATWBy9EsexipuiNnaOvk8K8LjDLFgiOBSsZvk
CCI0JlkTZCwHdyM6q+GGScK/V5ubS4R/e428mziyqfzbKrBqp7qdW2v1kPMGo1Xm7wQNEwKWaSqL
cFkW41/yGRAZctpYA0QM1KulG0IZub6feaFrwrppWl/Y1qV17FxXdlwiOtzOeDY/ehYUm6D2bDYA
uPM0lm6V3HTZ64taC0H31UINIoJbLWJCEGCxZRp8VmtozKVPxoU2DazdiZJVF6V90plmyvbriw0Y
UO2SUuHaLevOMzraXxtY+txGJM3BsI4B8KbwEe9V+6GEG2xMkY+MqCwHNBy37o7xzs48vjKJ3f8I
HjC6xFzcnpBBUEeII+d6ctaALxJTIOY93ak/6r/j97i9Gf5QmeXZAexX3z2Gs5fJ9TIPCjc1o1o6
slgXr1njv4VtxmO/Q5EMe9rNetI4pfpiqVjj75+tPDWj6O2lh0PZ2KFl3263dTi+Em45v12DS8J+
3xhYmK+XtPTutpofE0oaz9IFwhbyDQUgwnMOHVZyOsRUnSdFNUB0Y2hZxQwHmhKLYWosb8PdSw0s
oT7NeJcAskm5JQJOPwLjYrvjQbxx66m+VPYmP8o+7C9WsXKwxNdWhsj+Tagxg3DAWEvUSEjf09NP
iEzWj+7uSs0QyVohe11Zi4cPXJHOhJmGonMoOhEZK1ACO5rOgUfIkibMbex5QUZyXHkpxk9YMONe
C2yGpJvs7+osXON1VwyOKDxB7SiewDMMr9nb7YpS0LNPe2ZHT/jQWShv1irdLxLgVhSTIFOZPacu
wp2gj62UkX9GUhzsuzsOIWpCPk95W8P6qDX7czwdGR4pdI4iW5w1CjohXRxIhZSp9j4rRmHPYYRe
8t5jVZN2zjTUVEN4jU+GNo+SFMF2gjnwi7xk2k1jkzIg7EvcZqzAuVDuohsmoU14PihqzL0vfV59
GlmrALUJaioUhicn4rH8qWUhlct6Md+m4Djtg8+ZlWUY9F34lRd75KRdJb8TB4gI+cljotOAlnn0
cQBHRpePfatejxpt1GwfYi8eoaSHGii9wqfHAw6z1il2M+PSYsaO48GbOPIaqgBuzB7aYTxtS9zq
FVBQwIEceBLPp456K7QIZJJzlFiTx1+r63HNoi6/yLGufLNtNQ/iBU8z2/FDiKYyQ4pZdjNR2b5y
jX2qloaqRnaPu2COrFIbWd/z4ZwF1QLXYBztxaBLUk7ecSiLe7nOZhXAy4aGGbNngh2bGCGqnbpm
DRDyyv4+x/YUTSG5zCb9KexPWZfoVFwwRVOvQNb+TDiX0bAuLSx5sdut9QudduYUHL5G6cOHKJci
rMhAFSghOlXT52TK5w+bjFxoyrwJ7izJi/UF5ngnRgXHJ1kD6aMI7g1ngTPingYogSYALF4E32dy
bDmcwyONeI51sXrmv9jG1yXxsqUjKcZEYe5cXDPXosSpz+6S2LzySWOJm7zQyAgQyDSebY5hhxif
3I6uJ8EiQKDiyLXZs1oK90ZWh/dACDJMj5wvVZ65k+gYSCYqUGJ2JTYVXvuAIh5KMalKm4KMop90
UUaCsYv9xMlIAvdvCKV9Q/4kvedy6pqYCj2KOnRb4LD2haB7XeLXak3PivIFC8GRxAdM62COtuar
yKYNpw5Z+0AiJ6xW805doGi3hcq8g5Dv9pmJyvqgSmjC6dEc7zMAINyk7OcQLU+cmHpkCZR6FSmR
VTyRIthMEmdUdRI3IXzov3dMw29zRHjXFzekBIhHO0xa8TM5jbDVljXTBm3tCp53jvbb+TVjEY4G
CMDDY9+525PulqkJOi3omRkVM24LLg0f+gaOoOvoa8PJI++Q7+TdR0L4CXHLzWMUhdIsbaBeiL/F
f9K8lhkaBli3Cw+6r0YZMtmUra4u/UFraExoN5xJFsUA+PJd3H9GxMCLIZZaD4Iooktb8nfudemP
Lfl1gpdg6Uu66D5Xfp3mbA3hskBQ6eXHGvzszyfL1Ms6QwwRjM9Pf79PbdHKcW97gR95zJ+PWt4V
RpM++gABrq3g+4et5v4QgPqhG26Qs3vYz2/YNSwa2G4GP6BQ294IueOZoY5Wmv3MoBSc+LFlEk46
t2NvwnTi4DXyJ4g7fA33zUnkmcurtfbtYpmkKPaQwJGPW5s6LEtp8YImdncfBwXTdsEuLyOBEsRj
KTrwB6qLaNsq21YRrl/ttbvDEAnXDwg9j+Fwv4gxj6Ed36QJ803LsfMeRpd5l9ebX4J3lo2QMMYG
lJ4+nRwYWqyc6hoP8XPVB3TI6F8ZUqAR5nB1t9ymVyl3RUzAWxiD/0UBF6GQLvoJo1zzsjX5ADXP
yAGJjD5vwdOeA2Qmz370DanbHvaZSYv9hTxNoPFlc6GoUSADUbGWB/cl6c+LyqwoaHyaf/gC5pkL
dSCPdYi7NegtQ5CnjVxXSIRPIMY/tUSrf83oLxKF1gsIqmHbH3PWOnVFQ2O+dxcUCoZnEvZL2MD7
p9XGMJ4nVSGxvCrxxnAToy6qoeCtnwXFn1OEZKxQFHzCpH9C3ga7AYFrShlVd86Ee0jesx6/3P/Y
0/Nh8ixWqTepCWGYRrQlUVzM2EkJL736M22LdYwj3r7cFnX69C5y0iTTPr/AGgvphsdAcGkRfSvr
HmUe8AXPqY1SPhqGUOfsV1o9GdQE8EAdYb7luI2gl1G0JY6IpQ0YKIogL7eA/nQ2LPQ57g5MxTeZ
U9DgZsqpZi8bGpsz09GgLx3wbVfY2U9/Zbzl/JjjdgUG/zrXfJ0jRtoIkwlHDUU5h0Vdf11nftuB
e6/qVh2G82vV5r5bXcgbHp60xgMlX/WKa0zFu37sIzmadZtoAttPNDM3SiGAl3us8FsCQLq9scll
Kra3a7zOmxECEPhyQNY8we/B0fMaZg4nNyF8J0+gP/KZ2/JceVAF0Otkz2HTyV9M0rtQRl2TLTux
w/4eE1Ue11lFGeThfhaG7+UzGvnYm3Ut5eBb7JCzU1wnJlYQh3TJweqLtks0jnpXWRjAKfoucpZC
vh0rbYbIHHZ6YWbmcf4Wq6dUCkb0J34St8c9BQVL8GKVQ/EZnVFRnpjOHxyH0nLER4E4CJ9ajium
F9+f65lx6Lw5t9eVwaStRPUC2zOdZO+RhvXAXBOhu1QDq2KFZVckeyjoAkhUtaJ1a9iQTzvnYFjB
yeY+5EgmqjgW9ghzL9ryXX8qQ5GWv4aVdWkYY6i/1WKFvJG89790+lZcjnkWsMl2dxswKunxQ0CD
bXWVl17JrZTrLWb6qJgmI2nmBfCS5kd1BFGHAVfpO4OXBkaT/35k1B6i/3GbwN9u8l/jjoWMM5XB
lMmugBbfSuaOidmp39K/aGwXWCHHredywhoLtt/JJ2oyaKFMWZyJZB+03jGfuoIo+fteDYCZ444d
m9Zqx6ftqIyw7auEsvm8ZIWANruk5S23Wo8nlvq5qzF3V+ARP31jbYLfrTJ+vVAP/94KvXHgzqOA
pb6Tn3BIOY0ruNjlncQ12UpfubKzZDiTCs28J3ecXlardiqgeaf8JOENbdie0GUZFQuBmw+abATV
Xh8It2nlNUnAzcOxxiSKaGMWUbXI5H/Oyxf3MSBaHosbEmH0pcczBMX0stc7iQnmbl0TPAqzOUn0
LJ8NIxUTcv5lYoTXiewjDecrbO0xcbT39/7l7dHwuPEb+K78Uv7bRe1lWhDNf2wsRhErUl1Ypgcc
rSjOCO++OsjabjjUElhXNsYZiv3NDNZveVNhDC0g+VZrX2lw60739azbvUE6qQiYqdRLHAR4cOEr
8TAcQ+LXP1eUKST2sPpEOLAZaFlftHl42P0HThd91EmTZZ1Ljr5th4xTwYyaRUjnrG4uSZXZ62Kb
fxzMTgQk4GupxsCHJaiB4I4Dby6PTmbpIpiBzFdlkiGE4ueeEnfSB/tIqrXVjlDxzdVfAfVMMVJ+
CmRHfMFBAywM95NSPJMHdQM7s7DThnoM/41Jv7mZ1e2AYc02y8F7vllWxea6zBDDfNFmzQjeIYsb
MqB7AE2CfjeNqAuGKmvLJO0Cha5tVJKbdEtsNciFc/aK7rUuUynMosbGsXrZN/I0XSiogxgW5OHd
fYd6VLJ2AEhBlRb7KP5JMgGlXZhHhic2yCK6DfMPK1MDxX8aCKs2cdD/Ralzdx6rVndsaLjngcGS
kX0tZV9BlkYix21rsu5Ls8Vwpevq1bNKnCa+eZTAMTR+4BGErCLAeQC5i8Anu41x1v4G19XVQrnU
QYlXiYPb3btaqE7UNavbzlDiD3INHRkPJ3H0k3RBL3f8PN78ajxteZlEYnHoTmSTJgKPQKpmINgI
J1leAeTVp2+nffDHxWYgd4WVHnHk8zmAg2fWG6RJwRyre3K4b7J8U76fXbOM2aiL17RL+R0BheHE
8unphsyASLSaEHi7K4/FAa+Mv7dyx63XTs1JfCE3sj4jgQDZmffhBUtZKx8B9/tzyiv9CbHCRduA
bvCTXjBMbO6pM+Zl1wVkgqC7pufubcDwQtf5HwsN2M5WGar+t8Llt01SlSJzJSY8W91mptMzVG5k
qxEIP16yQ7uE3eltYtii4qELfcKn1Ro/U4MClXBfZTW7jO0+nA0mSI9gyena4mkkxjxWT5vTt697
FH1cyW3HDdwvXoKdoqQ9oqfElGHhkq5bk10c1gKM7apbviCvM/VLqip0PtAvGrXjNxgj98rxOt+Y
2gp/wJCq5S7qesO9hojfR30SE1yNA3WOrBqA5I74+mBT7EmMOtJ2iDvoJIOZYbNwmo4ttZcJmjlj
Mc78uY6DPSGLcvAbXhF3RS5dOnXYyPiucTQYhUhve1/A4RaWYUJhkxQnS6flQvnc4X/MNmEO0YSt
rOT846+MtXig1jFMWa05QiY8SGAZHuKTPHhEYWLroWmXTxn7W6PkP3ioDFjV54UIKT1pK1ikpGLH
0RlkPZjw0umjEnoLamHmEBikE31twXHHXqWrKi/wwa05kP228Ro/7RbzN9aWGcaIO4bO5VbcMNf4
W2QlLf2iBMG5L2Rnk0aZaZJj6cFy/16YuXaMnekIdGdoK5W3lLd1VAj+aTGHynGH1SwiNN1ahLMt
7Ce3qktcC10JuAHkJH7AKjAQWAzf2bkVMGoRHRnakrLris+uqbHzOi2c/64WwZJxeEhoMUu1VPxO
csdN1JzloA5TAIfhCeuevMLXxSPGKHD4vMydTlKjgtH0vhg5f1bz7VffvoBOB1USw6wrss3oeoI+
1tLnODamXTlq2WhUyD+/UXZ9+Vg8eTNH2twnDfDSyyihAv3r3k9Yo2gPvndm3F8bvH62QeN/KeMF
lbFI+9F6yIS6F/KiLXg4rPhSHFU7/NoK0MgTQsNVoV5G8yZzptT5hmuqewZbJzh0s7HIweiynvU1
B3VDjWTEZz5fRRiDFBC+adOr9HCUIAXok23KvPQ7S7PqE9qndwW+4f76S4SynqCzqVf7vcjkgfe5
X8ab1VSnu8Tj4duQLa+chtb+V3mEe87icMGPzCU/KBbLDuLgRgOnXpXBrowpp60iAlfrLqcajJy7
GtXE0p/bW+LJuJ5OsdoLbOMN8mo8rRXqUSJMyxNvWNhCTa0WNA5n4dhHQ30B9IBEzDMerg2snIvP
DOfy9nn2uw+/fQiuH1fRVB+E6AOdFn4y0bL86UEVXvdhtIkulvMCeuG7CFuL0BLpXRn6GU8uVGjC
pZGNBm09F+VcOThj/fGUayeinkqcwK4lVHUpkjLTdQIk9EeOrkajHslfJhDfVMtNOTgsfAZp1jZc
07OkE3miv3CZ+PafLDkPpBzlPswUppdvCzMU+FeXD+UEmEOw4Jn8LyafzDKEuC2GUdBQ71VLQ2SA
cKIIc3qBIEaQzuDzLPBDmo1qhpU414UkcoWOb+2e/ETtOYzVH/MmV+aJ8C1MVdEtA0Ek+dFbYeSP
icvoi/6+8HSK60TaPWRYpXc6YW6IVYraDcg7BjZxmMzPHCYPeZbUqlrUjiatpB6e39mLcHRHqmlG
8iXelaSeK+Yhqx/24VLb/azb+4EE+ntBy+WiyUNY7htE2nG82DQXNuaOxa7OfvlWMHTmiG5vnYDv
jPWOXK7jKF4SIU6A+8ij9ocqYeakcSpX2+XqecZmCoIw1D3NZWY2syupuzxxWalRogoCPO9/FqiW
v6xeees2rDQbyEMKosq691fmCxuSYzeIcESkAvQxRmAoLWiU0qr6JZ6VqaW+LiVS3XxAJnLBaiVq
KVcGmgQ4+y1WkJjW+PRTVgduftLkYFPsx5W5p299dAZIY+vfciuaUWpRkTvnyAoDHW8R54kJiTIN
AVfGUW7wNwDYB/ey+I7bH7c/HjhwEo56XT0pkoPz0bSoX9SPO22l4sQKqbw4fBSch7jYF8ZnzBJB
Z5E7zrhggKMR7Gne0if3y5fpRxDHt+8AN4i+z+gAJFC6lW3q7g5YeqHwqgJrddtFFrtBqO9TyOwp
MQEWSivrOZ142+4EEnNLUYQvpsAlZLO9W7TIB4phdXFhrgsBnTTNzhakLspCOlkAMDEN1GPvwNjI
fuFnR6pyekSqjdOMhqW2ZK3cCVGiZ0/fAv6mggqhsJ1jTk/Md3gYsV9Nh81O2AgzZBAfMJYjKPL/
STPIoErtZ1hB/jMb6rfNt188bVHR/Gy5FTwM32/jYii+a96xKogq8+fGhU6mEawYVoMw8QLygm0S
MSF1icmKTbTpBghzUna1OFUZGOedD+fzB/Y0FVN2TeFZ20iw9Zov7uu9qas9isMNqcnoTLeStUgr
2ZB4VuLt1f5cvEFjCb7pEe5cllNLmodD8a4XTTpemrV9khx27sLJ861XTc198pJdh6ShTe/VmvC1
CvfCU6rWoixQPvjjoJ9i5fZG1DZN8iGcaxNzUc/TW3UL0oYicXfiMoI8zeRHXmxOqPjgvU7zhrG/
F+R5QB4lMXkNaxYCKk4iOZSK5j6+8W7PZCytflDgi1UhnXRRJPUzpLD04RyQWw8ZtTBDf8NJO8x6
ZcAbfdQ0cIuDG/EJ1oFD36vg6SzPd945amddt8wJfwZdYTa5Cr4HqxyP84LrI62y2cXvhAbJdjNh
Rj8YSNFoO/O5YzLkfQkII9u9/9lgrDjDiogJwNdopIfDCvyhY8zubWxX3MGQ90L0O1XM1oz7JwSq
SerJN1QaBSNXY7RmN61DkJhRNFH6GtS1ZC+UqZgO6U0kRxYlhzJYURsGmQrjG0tkkoCLbN1AR9py
N5lk0gG9VcG9hNIoXOk4J3C27BRc/aVNNfb1A3SzOk6voWCT8uLgLlop5FhFzx8eqsHxu79SmAx5
fDYKSKQe85zBwZp9GNzRbfyyZus4LuRu0P+4OvVvYVy/TK7G+rQ6+WK7/WzCCqUetFm4tZR/nB8D
dU0i/pLYu8e11w4lNArqpgUvca2Fc4n8jFzTkxcDqQ56Feywnx1Jg+bwkgZlQRPcsjuu9KqWS/+C
+NZjZo7n43LqqBRlue63DsSkzAE4eQMSXZht0qScxBZ0UZjWfHowfZjNpbB4Ka9LzKoEH6AGM94f
fyN9ZqmRVRShFxhuIcK2b4uNmjijHrsXD10BgO9BMnYgGft9w8g5DWm2RZtOO2wRpOv8Wh5knzgj
NhQzJgdL5V+v8aEFNZmYdfzTBdgAxN52bi8ompIGUy3Pvch3l/mu0Txz5ADEopO0PVThrhgSUdR9
gVLJCXe9gTslos0hWsCD+HHBkr/Hd6tO6B7L9VUh3pD9aT89o33g8s/FZYOnC8kDaFIfHR/UTYq5
KmNVzAHWcWT++7ckDWuaMeYx9KFP6MlNuebAAk/ITqfO0ktyEQfxw45IFaXSPI7TEe4r3BBfh1rx
A+DIpujsgc+Wji0YAr4HTtNmGES8wcmW4FGtDsSI7AlbuA/HOp6LkKVSVD3A6FtTe0LmDj7HAZi6
wKwvky/48XBWhBfo0+E0lAX0bywEK1oZhw7bqrv/IQ7zLXwHJNcQ5EP2ZTWNPjmmQcPfWgdtP3P1
8l9meaA+et3imdQ2S6HGX02l0vvdmlNrsF9m9i/nWk+yWnAu7nuvODY60BxS75Oe/fkoWcHfXbv6
Q6REy5j5/q2HIyvQ9sipbb8vh56Q29FcGmBzKSUihPAj9NF2I5g9c2WewBZUCv4oxHDJblkwKY9F
ZtldzBlXL4x648bGPoRqSRkPFvVde7s38kyD+APLXZVwdRNQJrYDaSviGR90LZLU6qbwT1brgGsl
/pdXrJSaCWI26Gfo1Y3BJmO6hfrIo+z4bQ5NuUWV29svly/ORNDJ56bi5g6dXTD93hHXllk0Jcnx
oziKV5A3AbOuDtkZQX1Q6QJTGIhZFbtxOM9lUz0iz0c2cPfJUYmfq6daW+8y/hQMMW6coEBMUCmp
cKqDu/nem0WLJ4J7T78B+sYQy8Tx89lPRvE/iUbr/Lhl8tpzUrMXyVTKwlnnxyJx+tRjILlU2xjJ
ApZYvwMbfcFBDIPQ+37ppMTTPPCq1Oel4qk1gRF/IGslwsGTyI+6Uf7IJ8BC/zCXf+w4+oMlMzFD
F6Iypv76rUUkBFVdLOvavGS0qwt6i5hfltZy4zddeQppVgpB4CsaHYh7hlE83g1GWHgpSGURFvRK
toj3HmHKG7U3O1pWvV/4Tr9DV107CaUf3HKlQwWYy9LkXTX/u57i3cupxxmRmeyma1VM1s7I1J7q
9cLuLI6zh1kqebEyp41BNsRyXt1btcbZwrir7+hJtg3K76T6dGRl9wIbtPivCXw1n1V4qsrL7nMo
oPBENYl2S4ei25b71+dYHghFob48y3TdlzJmyhy7lj8QeP4G9iPEvb7RG3HZ05u9+mtCd6isk6Wb
RgCjb4YsW8XdgNTGVqg0q2asgsidWKs3P14fr1ZTz83hbLtCsWHxyf5NSgAzco2NQ13Ow3/+pekL
AZRWczLzJ+T9j5tpFEpAkUSO04J38fcQ4flX1E/NreEQI1gQa3/bbUgBxLoqrZlVK466Hshfj2Bo
bKnYfvAe26s2BuNIh011cGcSo6QJMJTqLgR094NAy+G0W5m7I1TjPvq3M2uO6WIgliEi2Kz+8tU5
EvKdvYQIzN0rA3FGnE6YIqjxx0ky4a9c1+NSJhFMZYgM8IuMhtOna1215cmYMbHQOPeCzTr4PHXG
T1hVgFOyAGjdQi7jSg4mAQyvtAqvfTJ16cwN8LpK+2sy9U7XucmYNWPNTuAtptxJRQQU8Y2x7lyn
DA9Kf90TUVRwRGbPIEzQNbZCCMaUOdD1Hm5LgJm97ntXXYq+75LcxDs/xpzhsYE8T41ZjuCyllQJ
mGlsmF8ukGOCSMDyL5BZGtJuXD3Zqu4SyIHPLljcXYE+r81h3hSpRfeGJ1FHdECZLuE077bfQLt7
W83UKgv7AZEmQjPTpsVeRhCwzQIdi1T31lnGI25eOP44KWFJQnJ12hC8gDt1n6HjfcPfnvsPbooH
mtnT3OJs4i8ur1VmWNavF2hP0MniImVrxPxvT+z24IWEY5B+x59P4ooEKD4ExDHZhWAjJdWyU3c7
UrwF6/EdKpuTA2oIdMRVXoWJTnzeIJS4HuxjkveTgczRLwIet7bSG7ty6pGAZufaagnOrtJ14c+w
6Md4ru5pbRC57L5EDon/MO089+8dn0s/DkPotJzK/C6MS/LPmHZGJ0GH1vJgrim2K6pVad9R1It2
JY6cAfg2/rtRu8G2a4wSKflKgFnz9FMC+bPI+VbrhHXgfF2NYiRLBzzSj/kNBHEp+nhR1ex59bwA
iEqo8jl5/6VfN7c4LXFYivM/O0lul2m83P50k6lisQiQVy/pbAIEEyOGGb/mQUM/xO3uS4T5Bdd6
mTrm17Fys8MNVtlwAJodUYID1cEodBGEcFsvMsxfyB8V8vTsLzSMkIZ340aRdlnHsBhb3E+tGsG7
uTYt14vCppA2YWVdpUpOGAN6IepK3SdsghOkJwxU0XSyZx+tmwYgAdd9E43FOF64ciWQxEzgjpLg
3z+e+SsHGlXGY/2B80pmqFxji5uMcxHkbjwur1YqXym/FRmmsBsz/ANqGhm+2FXAjun6plXsI/3i
Iu8MHKkAT7buFkJICAybh01R9IQ1zEBqwQd84oooDYuwiAMjIqzF2Zr7ozBiSoMfny6D10B9kffz
1LbZTZ4CJew0oO+MY57MWD4hYZlWY0OCa5Px//6VXXPq9A1Px7yI1J06mXYk6kS+j3hQqhQN5x3f
8ihowau9XS/CI9QgSkkVkcQrEVo4AJewwKIY2KGNfIZYVFPx+vQZYeDALXr8xaZZKw6k2MbneF1j
t4XmGiMDRt+6EPnIavx7rR0T1WXrCCl1mB1h/2uNcq40/xC9zvjOiITxkgeWzRcvt3W1MzIcVnID
tTDWHKTW/UYOokdsfQTWxufOEkpZgSRTSFDnfAN2yV3uhcVd/42depE/wOd45rLdrswE5rnuaUv4
RVu/LFNJ8zTsDcUGC5OgM3u8gG90zwdacPgHSIghDnQMZYEHX8xl2k5D9hMYRmPWT9s8F8o5DUoi
hpkURlr/Y9+0jt81xqacP6HbTvOYTrRRxLFmmEOz9d175NkKPCF5O/uZVTEiB0ShUkeYkEs/IrBH
qqMze8gOO0/GzzbOmkb+mLWA+wPLkgl9Pl3COw89/ecXfeW+CvO44aCLToxyYr6VBK7M2IynU+mU
8IL0lkxBPfhIdIC4mc162OnHVt2fyHoBW0q3B2AmEdN7vdHrCY/JN2LkU2qTSVvkJfwE7MriW+qW
ddU4I1rSo6JfDXdNRu03Zn73wVV5BzteG7gODm7PdEkbvSslzE2+WYz7u5TNVJGsAcduOex0ObHm
DdfCVjRYS9YMULt1vratgdOjhH4M2SYJLybgjXz5sSaEX9o6U8lffa8X4uguJXVib08YkcAgegEb
GSTRfHFAdYOVA8rlG7RepwqmLaoiqiSSqm8HrS8DSgmA8bHJo2cmRSpj0DzZgeoLJRB+OeAusBPA
ph84AUuu1VXHnTR32SmcJfgwIw2zlS4yFw/0HqoJnftquSuwdNHTZSz0DVife9fDN572DEV502cu
ukvYZ1rza6uUmpP8PmQ7BZE/Mc3HItM7x1F8hHODY5oyXZ59IGAqY50x9HUZmmfllcqGLFrR70vi
+OxNklYB5FCLAtas86cZmfXvQkJazPJY08LHJmH60HzfdiyihG42EZE7cPKZrsUCY+UBJlZxijve
4WUTXHJi8bhDuHNZAaRTQR2HV7qFtp1KjzZl2XuwnS5NmeL1ireAztJl+RxRY5h4X0+F1Hjlz3Ve
KcWmFCg39G58Nrll62P8IRnytabOv2zHooyuNK6gXhlordMY2qcET/BjA7kL/QJFdauHEpqFPkhO
ukxpzOHkDPDHvPv1R+UfA7ZwRW1TwwHWp6tyQnHfZVmfUivjUnwjMNXs5f+vn6V7GYUbQLcdVdy3
NdwBPsm9zAPIMLvXvuhDoQT/pol2EWpOyqcXzSfs3ZSl31A9we/5ooecHsjeWBqsEhWYPrVfYPRc
dgWz4tktXa+BnTRiOjjSnOJsIy1SRKc74NgYX75ohEFdyV2VgcI0Wzq2kZ56hkgQaK+GwvHFh7Er
8fx6Ok/+TqHtOrjNRKQI3pDphpintMbQ2ngmh2T5yxo3ZIQNjWY0lsVrFQBpRX/Albo8ZOYWzBTQ
D0f93ZFh3Df5cYqEOe4fAamK0OzLAgH0IT0JYumJTK3BQpoZt6fbDL372qqXPcme6juQgXctvDlm
bPsy6dKPIHTkvsZmeKZsEpJykRpEVGD5jq3U9rbRzNsFBTJSV5kUmudnmrgDJBt8HKlwt0wo0Pk6
e5P4MgpbH5QWoD7gKXuEPNFPImSS9vbat7f3e5vabtZgZhdpBTNGVp/xjjI1QJFwVhc+oQt5NNZ7
0+O2HweeVZQ/Yj9VmrigiXyJ7QVHUJs68Kn8OizNOO7Exm+Wqhthxoo4K8S/xdEO8pYHrU1DG3Ci
Wa4+2cuPcIYulikFD5zzVFeWFEzrXFDJZw4GdKto/tCYPWNOSx3rqAhdi9jV+TV7g+jNLBMMETcm
fXlsDaGBcRGNg0iMhxYkEfxzSNzSfqZUYz6OR2aPmgB15i2SwZEiwhen6XncdfAKx+sudg19cU0Y
gcNEc5CQ3pO5yqFcv2Tr4Q025MXWSpVvsvrVAMo9IKHHgfsrWYXq0KjfoPxyr4mfiogRqG5N60mt
Iqbw+5vYbtkGlXWr7hGonq1sP2MyM75mVFBvq75Jbh4ev7uiL9kYWpjDzOhQDLZmwSqfv5xbgx6P
pFjlCMWlhbZBTOAkcS7nUyTsJQ/+y+DxPh5qCxbe19cIoKCLfDqN2KrrA/N2pMe9eNut7BKjRCHi
n53asC8Q8jvL6x1RFRmBZohICcLwyHGkeNxn6wd4RCbnaeYXVUoTJblXP+170tKEmpUi6s347M4M
Rt2eKh7NNvUZcneHnITBVmEMgiJpy4Bo9jzP6RkDEnQO4RDKQe4ECaapJasmeUGtm6W5p1V6yAcM
GhCJJg0AKxQ6LJWymPbXr8Rz20RPam1hRg9Ci8sswRXjSd+x/C9Aa8TUVn669Umq2AbM0W4Xr5sV
a2NMZgPybIScDMohTl3AMmzKh8ET3+PKXgQ1SR5QSugwQxgpehNkii/uW+tmWpc76Pgsvppgxdl2
JfdiaTEtYivzCv1jALDFIT5N/YphWUPbn+LJaRWwwI04hA45gozMMmuM2qYQ1hpQYfNzosrOS6/0
pIVsXxpEh2BqWUzXOjCdvwCE2Cd+gyavmqgHBj0NmeV6qhDsFNdjibm431K2004PMlOHOHFPv4l8
ifvDG5/XFzaL6wlHw2Z2XXLcxb8eZsxLvVnfZ1zvIAQ5uuC1Frr9ngKw+wyBeVMQxIc4quMpPAxP
4lgoEBtAhOjotUsY3/wQIOeQUUaU2kuaDd0unTH39ruD1AYMQr/PcitwjBnwW47qu6qcCd1nEkhd
cs6+e1i2VUw80JXJkgQ7bOukRwoItRRyNR/k7DkqwGdcnCIWoQvz4lBfRjHjPHjjiW2MxL3kXfZ/
ZYOlV+/2w5I91bnSVckRDznnBijIXjj8KOhrCtTnWw9W6H8lkbt3EGRlqo0L12KEHGsCPXOp6hB6
twWqyiVkZ/qLXbYJxmvj8J0SiFeGte5ryJnX4MqvU0b5CIgOHHosEp0qjOrVHV0I5z4/h97+bkYX
j7bsaJP4fneZjf+U78K1rIBXoJSczgmtkS+/USQxGl+H0goMAvh8mBmJTtIZLq02/NS/ufS48hDW
LFJaEIeZ0b31S83lrOd8/eu/OM6tlqklgQxbirVFGObGxcLYfnQTiyCu9/4zzUSSJr2NbmecewvZ
iAQpaOjn4sKsHxg3B9VdMIaBg9+5cCmqq0wa54eaJxfQJypSdyyszhgX2cfuB5OxTQuBlCdrENAe
8Ssz3CcO/mjW0UGWB2uGnGIzc+i+bYWB5DwXN6RI3fzaC1sgp4vdfLir/Pa4Kp/ibqrEri8ET5Iy
602EGfSSXbeZmHo0ozM+d0SOqLsKhTCT5Oi9teHz+UXqZ6Yz7qac0B1YehHlKZHE/0qIG5UAPEny
diXv47PiipUocyVjCgP4myrZ+naTvJ/jXr5/XF1k5H80OPqoKW66n+KK2wsc50aYepTY7bA9+TFp
eU495gvK07KTEhpLijRQlLy7ulWGfS4e5Vf9A5nv7FPQTkgZN7QxPaUgpvJmSPSJbe2gt9dp3Vii
+S1Isn2tQ14msHrevIfm/1qqeNqNhKAL+ga4W1e9nVdPd+JB3Rmh2H1pWULGGApMf2VxbeWJzxQc
TdOb7J/YS8j7q2Ki6yfxzfWDvUZukTk07genVAHWBVxnXvJJHnU1nKn/3TxGXkCLyDoBq4AhbfPK
o0nglWNLwYcvV+SRaUCJ9iJuf+HXJvRpx5w5Y8eTt0Y5DlftbxONX4bzswiRk+JcLraaiXgamNa2
Z17fEHo60wwfrC80Wd2bnkdMcr9lwsvOs1PYv0rxbvZuj86AdVQPJys774ZJre4sqNfYkKgB/bMX
NGiSVC1GO9OMCTGK03fisyXKfAZ6CPCIyElrzcU/GDtXy6pLKXtSspvmLpH2JZudApZVKOXZ+A6F
5KLXcsA9/H8V9UEmtSz3YhQA2RWkQEDLQ8XgaS8Yj7ZJn8a8uZ+SwH7YqYyuVtIlpsrhdMPOWS71
t9ARLOqo9SMupinOvsaOeV6Y1tDOklsEcZhuNQBSJtZTwhwxEMc+LSBIx0QET3ZQm+d8n1FR1STC
q0TT4QVZFtq+5eS8KH/yLXwLMkbxiATso5zbBj8Dtngt5lH0YdYgWtnlAS9wPhJ42LRibcqiaRs9
lW6pFSkQ6KZFVRZLsi8DhCMYCmRdQDuV8oRU6yn5ElXw5cnSRpV969wq0afE+UR38w8nzRw6gJCs
istsEnw/src2/b98OPDiuyitufbtXGrq/inVjmRkmwjVBkR2HJy091wbsp53M8jsOZuHcuh8dWMQ
6TrPc7NXsPqgxB/nSSd93yl4i7Yr0SKTealX5h1TeyINXvAE8npMoBfcqwB0rByqxQICI4ogCqWv
x+EuDylipduk64c2Qf5MtyFMEDAbOJ57BpHKFH8t1zSaVvFPc7RIPxl5APiIp9CXMupPNwNUKUUT
/tPpWXx3uw+6I790z7oCsCb03ibZFoMdGqwOQF171QY7srrUcmCCi/ILRYuEa7jF+gRYZkWYnHgg
JMPpmHyKh4jxMjGq+/HqsIgnphTKKA5VMsslDCVpQNk6A2C64Csy845b9jsUZ9fPGvWfXdGjZkrX
AX8aL0x2mNR+m5riHlrdJcBIQxSd+o3kg3i4V8a3T9hJm4r+CXk5jjBZiDEhK0SFvBKrTEDEceMc
xsFkJ6FL1iifQnRsJ5NXAqdEjIsEykmCGsFnlYBKzVCMLB4VthkWFetLgJx1aFmkciJXv9l7yPZl
nvlGzs2oXS1pLnQAOrXjnyEQGEip1T/wI37aA8Lg4TEYpfA+D8eUv3/MOqIO9EYWh9rX65RhDDXw
NN9BdF+5TLszMZR9y4BHU2hGgILkoiBGdzyXze776l/Yon+iiFAI7l+kXbtOn4PWN7mUSobgsxJE
dCAaki22fpsg948+sdTC3k715Zv1phVo8dO48dZQuoLDAH/X/6ucQ3KNBhPG0Qj5CncPTcumEB2U
+Nu8Vd3gqID9o4dbjFCyd1BLfH8vRIco0xRO9x8FwNcyXt+p8FFjltdqxT63ZvJ5Aegn38rb4USd
Xb6eOjWkj0vDfOurM1o+O22nfae7gFLI0SQL2H7SCA6/Az+/82OeKqAoRrWonB1F/bDZdbFpJOdI
cx12NByeP+8zX34I5H+V4EVAXLMf2uL0Q5/GLJaP1b1bgpjIdsffXFGcfZpd5Jz/V3ptIiY34oNn
Uvy5ggtqLPLkyc24mF3Gsl7cszq3SeOKzjY6A1YK3yOup40PXoER1ozAdzHif3m5e0m2Tz6dfXNL
JkQ4Be2t11UABsV11oK9zIk7aj2TFVzuKygBF/1jgy5CxUSDWWeMzrR9ML3Zo+lSuKyxVYBFz/VQ
fruI/EqUT5oNroKDQCwAu1KDnbcR2MpaVeHmS3dtH4wkhczOumBkIBHs0NSYH0OPlkES9qTc9PuS
fYbVvJ7iY/0pXSIhsrzSpF6y/25kdywhdXXLZdGAAEoVFwpZfKvRnQ1oHY2RcrGthN7LorwNF0f4
W9W7bg2qotbFbUpNitP8mjgzn5ae8Kgwp7vJzZu/N705jkyDhEaviK9MM4M/W3fk5GabNq5gBAvb
7m8CLn+sZB1Xv84AH+J637O2VQRQr4k8vAC75uvTkcOwDKW7wDgChKiI1E1MiJlBQy5r+gWPOcYe
rOwBg7EqPZINJ226b7AoCiwfJHmdoNGtk2bYsSamMpXgOCieoDD25hYxhCqiPYmF5AKMJ+vO21De
Tzcc1UA3PnLpgSXqyPZLo7WzLXminD8T1RzcmsFC14GDTPw91r8bOl3GVGwY8WWd4leAbFaPgnTJ
o7Q5XBBiKbPzWVa8dLU7VoKVLVYGTUSJLyRSHf2xQpJ8zcepBs2Ysc0BQ1ivzximYn5rhyXjCrn+
eMe2hPqdiAdr0kUMIo3I2ExtDolIOyBq+euGI7Fuiho99caoKBQbKpI7lb0PWAhpENd2GBbJCUHa
y9ayKQjE6UkHz+3tyyDlSdqG2KnJIqX1XkUw9Kxn13RoGSnqlnAQEqj3WVAHnt7gt/yZAWMfCHYy
7CrYu+XAiEsAwhw1cux+pdSrwgKuuoe53usX3w7+KNKv25LNfn8Eqr3yBmoQnOh9byOX+kdX58E0
K7YSarmbNTDeWKBz5z4jMkZ3bpDeWL4VzD926M17LtgJp9bWHJSyTV3yABBT1i2HQmYU+AJAjq5n
MgMMouskdwN4rf/DIY4L2Byo4rDGTgD1qW/zooVgUz3p6Rwx50gXfDuvTn3/a9Elg1/QgFaFytog
JD+DTnbGDXcS/7rYTEsv/VelUAjJ0aowOHkzU7zscbiQrsB3DSY6AJo+/wbKm3IZfm6jQ9teBRz4
ZPAAXzPiPPF2sSkFe0JBgyKDKj/SNMjZdmZogbO89PtJEHjJ3KpsUGc7riNNTiDpMOkFUaIA252a
RjoDI1f6XHNhnq8F9RvzLxrqm/21V24F6VBanPR0tsLcqwpteQphPBrKyv1zBMuc7Gc9xQhE/1gQ
rT+qX6y2+deeuanrg54hHHzIAMNp+L2eALkYM9N9Ks9LzbLKKhIIIKqo99+yHJX6Cv9LHtp9W6Lx
TL7VuGmagX66cip/8nfefe34iOQ1AnPuuRGWThDAL5ilqIRvmwZsGtl08GbfGa0VHPYCcWiyh/1m
PE/zErHgxbhql6TdXOebt2Pr+mwK0hPu1T70r5XQnCcBVBbXdIxcaqiMCFujzl7kotspukG7aC2b
1dz/+TxsT/15d90gfsY1WRdJjSbU1YdAAJQEZboHN0Xs3QSS3PcKkCY8DK1J/GuLCehwlVZIxtfF
W6W3Hwj3yGzOt/im3CWiS35UcRiOg5XW+tSFTuWbi0lgNZa13sw0nbwBDKJVPdOcmwt4wy7Lv+KW
+wzlWd9PsKb5heAVRMHBgsAABUhbimPA+go/QitExiCaCSPVl6Cu0FUtMrIkVTT/8kqw/d7zgzM9
yft2EG3wdJNmIKlfVz4p07qfwyyaMFWE4XzoTU9rnfq0inABFWcAzV8h19g1ze4LbYPT49vobW1M
KghZdIl6TI5HH2mR+zLzaPShYlCZipLpBmx7nFCF683QBrG3tL1djuuNPa+p0zmFMPHVyUbBUv7J
NZ215s7KmgyEZxO5oatfjEPtuChiKWHMb4NpiaQZTehKqLP+YIiAvZgH3PWGlFZSfPVMDo0PDs0h
E5JGFJ64mSs/H8Dji51zMnDLy1C3tSX90zaK+bAFfBD0DFYHqRfxjaPRiiYvPHhht/Zg1JWSAbxJ
DTn3pvlnLt+XfSeskOSZYm5Q6dj6mzdIgdGTtPUMo3N0IRkTNkcPgm4cF/OglZOu0JLDTGyZA+lT
V764PT2rN9MKJMUCnQ/Aj8XBQydV89+gWYCfPw2A0YICTShY5MnpjYZ6tAbQ+tQmVUf+21/6PA3z
XLS+Y3Pyr+y5CFkl4I29tNtMqnm49nckxKYGXgCSmbIacAtn7okup11Yja1ZF25MXFqlC+03l3G8
0rPGUTNc7OXgKMOQ5MZgORCDU7UGhVVZjimOInjOWfQimA1Ci4i9Wjr2Uu8vZjonS6yl6eNA0NNu
wovfFM9AL3X74H07IqNR9IsIW8ppOwZoRd26iR/yd1nZSAyVEJ1jRn4Ww/8A+ff8hOhmggtzp2i9
MIPDjfa63C1GnQNeAZW3q2pEHYYvTfHQTjXay64BoC4De8KTXkSKq3Tfa1uOf5JOR0q+R8feSqDp
OteFz9TPag22FtJux9OQgi01sBJzBdVa1aIB4CR2E1m2q9Yrq1QAlBU/jZS4sPV27dJx9KY0/fmU
mak7OmYLzXwEbtgrG/jzPmC9zfNJS3oVCXkMQidnB+bFNXUzjx3e5a6G68i2IqWenyruVPUv523J
x00Rtzt0h2iSiXIWbbyFeeqDYcAcgvnXL2mb+DLza3N0eda90iqqh5FJx1b2TyJaNvIrUpA2YcUK
GgPBRLt92+OL5RtmADKjsf0M8Fu62rjSba9tyxH1nwt0F8kVgLGxNQ68DRQNqQ+zCL6falek600N
0h/ZLUbj4rWO7dqvXQ+p7qseAX/bkDHyFNwWOrxDPDpgfNcQ8R6EpvtwtyuSk9Ijn0TjreeqBxYk
RKyPwFZCXeTKZLk5gTELJrBYbN8gzCfvodsLk3dGT0M38RBzqvWBSxiTdK8aYzFYU/9tzZJLAWtg
otFxAuFfWb9dmyNOs7L8MsIDZy2xVJtUi9Wcjz3go6ZJO688bKtJHKTqifNw1D2LgHYSXQdP+wso
acTBE3B8qIxKp3rRmkR0/8i6KXL4UBU8EaC6k5ZQHv2yVvblzZg1dqg+QdCIaBGm0pOgjXod8SID
7lbj382fwO3md+JP9nK0VI8bALeijK0+LszjdpUcPuzWhY5TManDfPDju8navNf0eB2Og6/UzUi0
uCfztpQXLkFsHL2zXR2XW0X31f6Rq5YDijkN8R8M79qT2nO2V+0uwyHVCTyh38kvS2V4uXRlkATQ
ugIyZNQ0wxE9JRZrRATKTKEk6AYTcTDVvgY4gCOvZ8gWbItbzaVAt962+pUaW4XTI1Ksjo2lxD6O
iHKVr00xv5AadJGo3IChehc5Zj3Hr3/YypbCzr1Xl7f3NKynxe7gnop6nDKCb2SHzEgEqnogOAA4
iopgAt/B6DjZ7jr4sKRoMyiALJTkiRHftySZxtX4SH8ux4uCjQuSm+q9Q8u0TVq23PoKVE+Xp+Qc
Kn02A3xO4dO7xXeslHObwDAxcvum3cwYPxeJS84IZmz+l0AwtAmtg7nto7FAxIviFOFRB1X3PAy9
aWBdpLG3rPg5N3VabqL4V7mDLGLKPwzeAfc05M2z7W8T8JCQfv2DMGSlLmpse4TgOsLHJGkfxgO+
157etcXOxQ3fStChYEJOLhAkYF+Y1VYwJ0WKE7jLoidPsTPyu3nux3Y+sSJD7qaLTeLf9NBXX2xV
ZwSCikJ2TW3FuHqmqGmmtbmNApD0RBJC3ftAp9BpCVZFyPHDb57jP74xrmljixvGnSPkT/9Dmblt
fWXxGvODbZrCN9mJ4VcR06tRIjyJdrs7kQHMOCAQFptx2C84AIuDbTP1gt3ZACiUgq0vr+O4INJ5
uj+FD/3Uf5MmGhHDxlmRyBQqrYEbxExH6GkVxidMt5/+4FgI9maAZWPg3tH1yIF5QhwWZDzG+PdZ
pKivGvxZraN3t9izxhAfUXrAZXV16ymXlLH/r5iMwuxnlV0tAuJ5xWm86m77QeK4E3G+y4vuXi/2
3l0i0jfgHASoUbWN/JA72Iu1UkpOP6uffEa6A6Rp2towtOdkrVcThAIdJrUx1Zc+e7q2CJ6hLEBO
HUQOZ6RUvvrM9lIKOjNqQjBXrxsFJkCQIO0egPWnl3a7Zpxxb15ER/qDFLJZ0Jm7aXkvhWP7FauT
cnnJY1PvV8cg462SYnZz0qB1R341EPgy0q2o2ftavVME7vSLYWsZRgdcl5nt5Be6A5XowCS05a5B
jzbs8Cv0Noj1fOTUv0DMfzaXg72TCRNP2Lni/O+wmDSvZJJJNj10xvu35IUE3bBNPPqcbPShMbV5
yTYEl2ZFgUWdcf2zdsgrt/N5buErSFPgRFnkxUJhu3A1NkmljXX3fG3gwTRoBEthHjNmlk9Jrexw
q6m3uq3Ht0Wj2POMwI3IMCPPrm0ZsTJZKEnZfCVS5GnmZsWBpxkNMosdxDUJ4I1ei2iCmGzyd1NF
8i8UcBM57wgGZrUBdgPdtZwYKX0bV54cw2lhIxOwnY9LG0AgkfWNNviYsnuZI261xxeyDcrxzpuM
dj/4XepLzi1BkZasnaj14Xi8WwWtlCZSdAJOy2RF5B3DaoafmU0ouFGTcGRJ33RDHcv57o//bLJW
FiO/NS9ndeeZEiIu94Iq8raw/Ucycd5dHhxbMj8oMDf3eQ5yoxlGKKf4pMWc9dfKs6srqOTuObxE
WlFzxwniWNvE3vN/lSFB2ylUHmF11A8QR4hJJRox8zND5lRO9uO0Pu2XhXPo6XELxF7Qcplm8bVi
OPiXDf7HYsjSLPoZwWnezFw5sSX0dMYRQ5dg2fd/4mcvKYFg/dxZfIYlEMeob2F8h/JWL2zlIA8v
A7OZ9igr8m4an/HHqjtdUmFqGDR13e5eKJqq8E/yXuQMnSWZ0UEg2E/w2CAqOjLK2ndRou6h2V2w
rkuRhyWXs944XM0uHzVb1KZDycudnuVlj2MMpja1yqPGw1jm9+draBBRCvBCYgYkmnIuuvwldS31
GMOtpdk3o+QB+tLQZDc9BqF0CSKcb5NhsVUfnprPxkuvwqqGlxb5H+5y44JworrvokEuE8zza+mG
w8jIIaHeUi3Xy40g0VKOOYe46XNavnrTiIihgdx/AwutUJrKQSUll+m+ucpFBbobwLVwrS4Up8Cl
yXewjobUdN1wZgP1W5eTAPPYAy4TJTi+zMM7+AhME0tBQr5anxpijzgWesJWSajiXYZ9G6oSHM4d
P9Ky2ndRDbeYGcseZvSzVxx9aU7oDOJ9X/tMfeBf/yK6nhRaU4uqyCB3znOauPq1tQslvewZUTni
fI1bUOD6l21uPL9w6MmLWktjgI4vCxAOnXBfAH0iCuN0PgRI+61A1hl14VZN9aqs2uPL+OkVfWfw
4KWY1jDbZgdMiAoVbRVRf+JjkfjjxFEQTZV0KG+L4yf/6XMBoesWVCcoRXTijv4h6mSXWNqTKiLG
bqa6VT5teNgOrvb1I4Bkp9oYJVGx09BLkJPNl45k7GAkO5jFKIBN4zIzKZGh5BZLVnY4iDosRCsE
eit0Jf6eeCBxOhqQ8c2nsa3fln0rP25lTTeIF+2E6xUVsFXnYg+iqwKaH5n9uQvYayRMUHvonyD+
HGhQZqZB3JFuMCKz/68Qer/Punmx0xfL1OQl1EzS5waIED/AoZPdOi4Q93SFsa+qZfFkcFSzjWst
Yh+aySuVOKJTiPyX8Yl7RVadwiuoDTzsmsFzv/Rde49V/0lQt2D1U5UtR975xv0DIEir6hxmky3E
rJwUbxJNoYMpZqeWrIEy8Ih5az9tvCudYQ8v2NSQGqFOa6Dp56S/DtmGShIKFIl1pRM+cHLLhEEI
1+47iTrIJ2YAEFNj9yombaNJG3na+N4dL1CYy4Wfj7bcvaiwkQHkCyb8ZR0M5YMZE7KLoSb9tv9K
KWfuSVZwMTWvOo+rNN4P790hwamwLzFu1PAtZYSwoCdGxzTBYRTJ6AvaRFE8Cmbrj5u4mo/o6e8G
jCtrmFMl+uu88YiryW2L3mdVKFhardqQuxF9DqBSjiSZ01BYCgFaLk1xIe7PhCOTN0LuVt7NT0Jj
JkotImW/+T3AkJY+ShNENYnpb03ZIxvw9GSJyFw+Bb+3FNbju1kO72Edeo6LkTJOqchyaiQMaLf9
BU5LxnteYkhu4kDFLeDWsLZVh22nTSUfjl8PqhwxgbgFPkjXsAPYua+MTa5a0JrF4sf/EphAbabU
aOo2kqJngmDATNdHXoAqqIlpotUKKxIf0zlLzGnp+Tr3jwkkTYEZoRrOg1lW9YYMVdHSvWcMbwdM
FsbzR7G+01V8kbijFrkniSAZKELKwvxh8yh6fYfhWgo71aOSFio0AIV1Sb6kSw9pgBMCi12m99HX
FSPpYKRToVgvDPIzp/IXHJShZv5kJcUrJH8Ll2r634FfBSDrD9EogNUcJkJYZuq2Pu4Gsg+JXiJP
Hm8oz5AzIWSKjQvI5ZZqWKkWAib7+8etpuOfv217Loyk3MYXXjreJL77CHhAaARijACeyMTMwwux
Xh+vmceJOCabwi3WWUVEwyk5FRwTXpJ9Pkq75BW0vYA6xuGcgAyX9EPGRl8HLr76t0FU4FUWkImg
Ee0qh9g8bu5tEcCydfUs8Zqc27VGV4pndLOuELhQqvmGt6m8Z5Hv0+VB1PaJXuUehlkNzYCfXTo9
Puw3fF/B7oZq6Xc2ObE8O0X1a31PqWHY6LdpjnfRIeVyc9gLXEIWHXLPr7orEW76TNYubahrtrVY
x2+759KGX0zbKMVpdk63Ol/Nzrt5uo59ECpgq1O7Hfbb8a0Rp6zPZp7e6tfVDfyYmx/S3kMKh+6V
b8SZvWgJEIozQLDUR5sTqFrLp8v0QHobm+UFfJ9isgt6PjUpAVlAzkDGT4iTmaBiLtCRYSKWH8Sp
TIuCWPv7TgvzS0aCJhD93cTihrtELXiSb4pI4oq1F3sYzUtb46TRdxMIpQXQQfzCOFP7cpBc2fFL
lgb5FSTfRJaf8SE1sI23Hs+F/CiCfSy5jqWV4vTprza63h+POyccdSX6mMKsAIKKzAP/8y64ja9F
YeGQ4ErMcCRE3X2aUUGojR8hYW2C+NaogGmZ1zzS8aQBIcjItK6I3AM6rqazXL54zsHzy7Dr2DOt
Egbhsyb+RjlbE3RJsG5p/kP6m0Gos1BRoThCiBgbUwykge/SOnftEygACq+jvpXBUFKVMRYZVsjc
cVrZqh1vJbjW78GesGV1cEcst8A7EiZyDPaZjg4r8Q8DaMMLescz+V4X5AjroyBoiJVOkld5YNYt
t6LWzMYUVvYKmW1I7rlxlKhKc8S9bHs9821eKWtbnbz1lQsbCLN75WtXoSbXFfqkHrUmKVxee/iu
xRMhCT2Xu0+oFMIZUI2rYNb/0HbAXhJFMQBRvHRxIIXCcGv23MIOdFJveZ7I4EzmS46RweUO50gH
oQWp3JIzURF8ZsyGtGyb2brDJLW6jJJsk9lhFID7oniLXb7NLKiVHyAp/+5Dsw+luONBchpU00Ms
ZEIq+7gkXkytnmdY57hwRjRTiwhflDk0fUT2C1yxVIj+tNMhe2k8KMu5BFsdIRBhrQSv6/65hcDy
kD6LbqxqD1nDFuo/9DG0D9DTSW9j9C1f1CXMLbsT4yJg7i+POa7LpAf090ef1Vrwl5ogqVmFRCcH
j/CMzMJdTnFqE4ixLG1EF9MnJ7LKubOqoRtSXb8IqvK6qMems20tS+YufVSwCGY0NpA38p6/xTnE
ignG9n1DkJmyaWVCr+FVQZfBMNQ5LfsrcGOtCel5L0GI+GcyYr8kolRqGLQ5xGodN0GioLaJyHAS
G6lWoMLwIdv7DVyeJtmPQJtFHhr9T0JjY4H0NrkTTIeDgOwNuueeZj+SXScUI16Y4hUGWcWFIx/F
h+hBGYMaLrtf6mHN6sZePmpsbqfUW9z77Mh19OB63FBJrCQAGijQHxbZW/yv0p34TBiEsaB3pO7C
NsSBfgNajsMkzcr2TztPYi0VOpvu6ICh4tWcAKozr/ADOwIM6SuiKnom6JZmU3LWoOXJHyz1v4Et
UNWbo8rbH7VUuvemPb45rrNoy/suyxgtPycSeklY2Bdk7aT4A6reaFIoLG3UbsawVB2F9G5SHKIE
77uqcjkHlK/4kcRSlWyNGa5kXuRuWIkgQTiZQT8RumQnuJ9BM+lEHaPs2BksF8Cw0HgOLifV6ncm
9+2s+qOv7vWL5hY2pspfpdP3q+2MFcIk0ydjaoMQ5fiAosykJ4xmFCV4xOGBJ5lT5/vl3eI7lHDz
97yZ2+chOs5aYEWcHPZ/DUOQWav2Okef/pJB8GvwnRbVwxaizmAP6S6qXF8WhFsYQsL58BGu41sU
8V+0xZcO+T/UKW9XqXvkoO+0siztTb+XAxeUKWr5/JGlcFu6DoI8akdxRcHTXv5cZxDhPEqO2INv
6r+2FZmOPLwnxr8Punt+KHeSMvyC6a19zOPVIhvapBD2UgA2KNL33zee6cofPN9/6KpBhdDHoY2o
lbbgl556nNSbFYM4iG/HPSpUru+DX+0B/gLGhLHJ5V29ScZOtSCh8mS625Dl0v5piZ0u5uQ+zQMj
793Qd581NVVAlMaDJ9fVt5Vy4c1srPGAHtn6wKRgKg470LpWs/GzIujzqCn/pinFwzlftQwdXD+Y
w7+SoeGQ7qpUMB1/p756hoAgyTSRYwS34kbJ6Zv67w6rnttEoCQ4A3Q3J6LPISqz+NotWEiUhzGQ
QgPYxNT9B4Z2k83TMT8MDSMyUw8brdKr9Ai1YHb1KzdB2DT0x3cnNps71srx1wQ79h1lP9vQIPar
VRcS2+dLQHWfKIrwRaYxmQwIskkS5hDSiPloVnq7GaCkvTn2DNtPj8+ZRRjw3IO6J3oDYUQ5RDLR
HWOJ617UxDHMnzZQEv0NNR84HchSmVCte3NzQBtJbTn9AZC8tM7kv7PPhnHg5AGWfChnKKx7/ZGu
TGuPMiO75PLUtlesMVdQQYJ4omYf52CwBlMVlmHQRneh8Lt+a7Brcrfcrvbq/RXKMnWZ9d17HS7P
5LUu2ghI5tAbpzbzqvXRlrWSIbFdyfWDyLdnigbXWIuN5oyJlTYJapuWUt7WQ6CdvLE3BcObQZUH
HJuZ8j29iWyS1vjp5Hvs/CTtg4xKQxIjjSzkhAl9CkFz6jiAQzphBL2k8+jlcbehPRMByTsnf081
2s/SNhF6sGALaEF8MI3n/oWMkgF4IqSBupPwAthC0vqpC+PLZ2rhsV2i52lkLtMsN7ipFgD5dfMj
VbkM9O4fetgrA96gBt1cHIiEEANdLkPItQFz/JinG7m+MR4iMKVngMn32cPePkpltc7Cof65dGDf
9uCjAwtqzbcVv/0VpDoBptUzhBLDsoTMdsI6R52FMIx5oHIp6vLzyoWiIV3T9mvIykzVviS8t9RL
AnaCoKfmfbzgRDinnfw7oQ8Gs8cNEXFlSAuh0igavwAEikIRJa4YnVovE0M+LOhNeGe2DWH5SM59
B4CglJfoujgd9cFfqKEwjOGY6mgzCSIFB28p2BKEgBCE547PJb2sPzYyb0C9YikT3+/KXggCRHAu
LGFGWofn2ZkJ4YIo22tncTluYGtpM1ckRuyvfsbZcC43nGj8GaxY8gEvHVDt7tbnJa9x15nkBxUB
znyMTJ/WgSrFVnV/15NN4JIxh5eA3N8hcssZwLbzgHW7g1g2q8c63gZ86kGOgl741gmu9RWuMwgU
dmaHmSPnqOX07e828t/8ujsqy/chjz5tldyhhZgi3br8J1BZvzlo/KqtEO6eSb+r1zarhLNK4kLI
sFUVbsJLzU0B90pffjYYlmh5Vciudbb7y6WsGavRcc2hqxW11yh3rsAFdMRyehLOq9NrBzswsmYK
vijhdDcmlqOg6ucNoOsZXSV1BXAxLjwLcRq/vx7BwU7qSWP6SBbY0mChVJ1ipJ9suR+K+CJDdtUF
Mh+KpJiFE3NIoB4AUOEmfFdKbopraduuuA2FQbdr6ItxR+JxZi7JWU5lb6JV80FfKPh9dq/9W5Gi
yZZNqyo84t8rfzMitL81PwuSvwMdIykZoNFP9m7QOdKmVah0FAS0LFzKdZ1c+CoPeSdsNMDt0Ody
ebW09pHyjKuNiJb7CtEsb9GVf3BNNiQXEN3i903NLfM5RKg/flItSFMxLQ7FoMXUCFI9o/x3zcEG
YO0LTrtA1hkpV6r00eCmK/27dIeCoTC8lpaCso26TSPhyNSDTKx7VgBpcnDaiEmzkzOFI/iuv0di
bxMN8XcJiSF9xO7CByxWoOc4ZLnPdQ8WzMy3yOOWkQwlDsUxe2setf9ilXw/yFO4w0dGSe4VcTjQ
3k7dLVXvNM/jtLLrzR67CUBscP1dN29DpAtUtg1g0nywVKqTILG709sQZJHdNKT0Y2Aw+x3u4nhV
j8bN/K9EP5+3N32YpNLs6jdPbDHGfdqUOpildjkUTp1I6s9YNdF6tDAtLYI63TK9EL0ou2oxCJ5Q
ypSOJMSkchAWfbtpJBKWckc1otTaVEALF5baawWLQAabBQLR63dR61eHhncs1Jc9SSrfTEYD1pvz
/uoxG7GJRQmulf/R1ImydD1oTq+ne/Y7rhvgmKEgjWNcLu+QVMTlrlvhWyQFV17QDQ/ZHKj2HcAo
eT5QOvNYdwXb3bUCTfuS+MChWDPXM9/b3AuT5B2/8mu64I6GtmKVOJEWbKDXI/1jFfau7l4rcTnr
dOJ8IIsKdPLZV8jYFjGxrkpFx05h5pwSuBWAsJTaC0OWUJwjDPfpFhHidPgI0VbY+qUzcrP6MdsQ
rZmf2hHrQejRk7xwCeOfHlSf17r8Ygjq55oyTEOZMGZssE7CShxR4v2QgfdvH4+SPw6owoB9jSK1
yLqjQqRA9cdkU2EJJDC4YFAswQOyhPec2JsQYoT0lvHhr6/mrz1raVEia1BahOMwiaSZa8HsXWgM
sOgcjrq4XTVZomQgJ7j0yr5xTARd7/73DWKXLywpx3WuUXXVr3J2DkMEz24CNg6xVQE1JSQ9Pc/w
ehyBQs4pQFPqIj7Q12HI6LJTZ9h2MakdizJxeyJoV7PIDSKSsRJLbjQL6TJXGqREM5DDFNVCAyC3
0W/FrtllzZKEbQ/gKm2pTPmRgjv2HTCUosWnA+4Dranun+BGWdIbqSe5c1CQk5MohHT1+iQQ3Nbh
3Ra+Xr1E1TGgShl5o2kYD01J4qCDGNkI9kQ6/D/BXf3z6JvQaQEELlH8B6i+VEdFhLgskM5MnaGO
73+RFz98FTN5TDurXCZDjfFav5pk8lf6Pz8gWHmvdAIf2GDHCxJ8BChCVJ4rksLQ8Mu6AlLM9vVm
9Vz0IqoUyRMA/TV79vJynNFBQ3B+uEoS/NXvcM02dzEdkDQ9CHTDuxTF63TRrpTegQzs5Gbm9v9T
jv5jy8UlLzv8Z0GA0/7C5iUCpojjZNlIFc2GedIYghjduvE28rWE9U67H5vu3GFQYPwi3dxAh0/o
tDSkrdqBAaj1kDUr9kOQkT2Sh6FLxJyNWE9/75DKUnoOzOGQ/BZRRrMeopuUOJneNb/9HpJ1doeQ
eJKfiB3i/mxCk8rRIjDlwalBBHekBX8Kdug9S15gdUrwVotanyFKZY7f33lPmvH3yaZ3Ukknwplh
ufSM2Ke7nlKd83ikjPmBvh5wTX0Rps7WCBVkHhLmLZSkJgIdDB4xUSJDk9tI/tsUkEIfq0h59Bcc
y9VNJgHHNFvdPpz4WqCFZ4/L9azf6esvPPFWZskpiHYltlfLqBLyUpw/IlZ6c1OFeOgpY5eyv0zB
Gz8+iZoRcB6T9PytGK1mRj6rvpOci50X9nvyHqhdWwgHavOCFT/2FltSQbghYtTSRP2fRMXhiuLF
fwuVHkab3BJl3z2msMygX3AtIrwBjWJqk4Do3utPTZJX5EivXhxo/vSdPJuk1zinLAXfGi+0E081
CMTJNEX6S6MMKbB9ItbgAHtSoHI0QMoRC3bOLNNJEdfruriQ5RQJBLy3tsvbpKyfdws+32eW7hpV
05DqbzTz+tHL5F8kocbOaCYZ96pQPLyv+wUmggI7gDgSGtKuItiv/aG58HtiliVeAV/QqfaZqoZ1
vqXPYWZHPTkqTXQ/CvDfG0fylGcroOdVDugXlAFc27krpY+JzLGqhWg6Wg170Nso+V/0LkstVMKy
dEEa4WWqm93EQAVOZ9vBSYuQtpXsWeSfLeEMh/hzxyXAuCDqKt1OYr43ghfss5PxyLZ2ZTk04Rb5
DmotK8O3cM2yJCqwL7ImwAvVBs8qkBUHTAIWliootWocX3BzaCNsqd9J/ZEFkk0gNAUWJIvOGL8K
1SeSskotgSNRaYkBMNvJdmx9R/RVmXDp4ODXk8AZb54vLVCtwzPTBpPUFuc3xKIHS4nmQilLLRrV
5mnKHlvNYpzezH8Ug5+NXTanwhS/2GY1V0lavC+cuPDqm16dFhra6QGnyHmpqB1ka6y3/oJYE9W/
854sJ/LwTpq6pA1jEnTdihmXSl76kbuXmZ12zcayFiq4/ax8DuDU8eMsUFvePl9bpDUQ9GY6clFC
sQKZ5NLYL5BKr2jHvgFZDeowl8dMWpKmqoKnR8qhcC+kxu51ltxb71LiF9xBMLu/e+rUnMU+SK8l
c3J2KgsWwDhtLVQdvPiZ5Sk3lbowDdi9EOzLzL4FJT0+kA/wgsHZzCxTNouZe0ugoc32dgb4N0AN
J8ZQO43CUWi4zWCpKUt1FYBLzKd6NOFL5Z2wRewBz6tHQwcaG/dLIOkF9GvwXsE/aMzIhDz6KAni
geKvzXT0f9u+cId0/cqWSbVR+/gdTF+a2zDg4poRw3VM+2fea2yDt6T8nZ7u9exgMXmJ/1gejPuV
kcP2Ig431YnUt+CXU32B3myli256qFlfYdpN/gDjxeQFT65bL41N1iIL5VGPZLMPCbo/DDplRaJd
yyS8DU8Ut+zpbl2Va+1TeLQWaSaQBdTT7bgvBPPsMRvGzplOmOSKSH44DX4QeBWOtef2De+HpRaU
8BYBrN2VmAiCrfpZ3pCMzJonMvNvTw9P+fOrNtCmeDvs5yykc915dKPAedUZBYYelu2NR5cNQHEP
Oa5HTgm0I7C+6dUqUb4vNDVndBvlMk/O1p5X1mF1Ahkaq9gxLj3HC1tdFq3VFvj8IGSGXEXwkUWq
a2YBkgOs2Td70KwOEBk0boHtygTOs7laRRtP2fpeydmt5rvL2RGEH+YG64JAwN+MhTnj8YK6Xjf6
KaOHXhry/gjEydxixrVfB+cWJpJb7Tw4BwVT7keTh+mOsKREKCpewQaTaecz9Z3d3WosQ8zS1yPx
Iy0sphECmwsB+eZCbIf7f/rpuhMhGJ5UYz0Ss2QMS13SnKJ/GOJYzfNHOSq7GE+UYJUAccwUr2+g
EQk1aCc82PAEI72dLcWRp4/FnYnX2E/UVqQn5sZ5j8JKAZ66VNIEskdo55EhJA4MDbmjTLqwEbSQ
zhc8y0NlW16esm57qWyQyfGQPhIUuDNsL+8iBcooHvK1A+XmZyyXr2+rh4p4+VVo7pRVJLyGhxoC
dUgVg0u6p3EIbu6aPcmy0eho2CgbHLVqnNJOt/xnp1SusdUdASTgCarE1icj5iqBQEKh/1zKZFI8
D3dlaDLstw0iZJeHMPecnpCZ+2FMUF5pOgKLXd2zaWs9NEwD6Nwm4eM80CuVzGrrdm/1nioquk6s
G+HzoGCmr48mAtR3d+grRk3IISM7aUVo5HTB4golbMtHOA984g7m5vCvty9qcNbXobItAd10Q5UE
wpAlVgJHnqRwxhrkpP9IBRr0jBVt/Sr3K63Kb4AeUxyREe729k7+Yb0rOs6f9jko6e2q4uvNLLn9
8+8Hq1wOdlzz6P/n4YJ1gDZEVxVZii7vwjb7wkh7eShFi01atIy/H1+wajX1we5Iv2XPzT3cL9tg
DGPpB5VLMRU0NTNjsDlaxLsnkGRZHko3IyeFAjXEol1BmuCOk+jgxJC0U5h4cRbGNk3KG7AAPHPG
Lo7JlbAFgd93j6PPjKOYOU/p1wpB+EhILp9GUk13Y0y/hpl2uepbQvOY/Nl94IdzPDCneV/BecjX
DlBVsguIzcq9NTPphLrLV4nypbKpLMCIsXMYKRepuTSZofIP+pKaEr0QgC0hdHf7z/kFWrSji/G5
fsEOqlZhx7HnmVL0IF0+VNLc85G7aJpVRp8h6AJgZHmwtE4J+vrSLQHY7ljG1OMKYeRpfwxMGYFQ
0PnhjcXKVbf46mxBhcYgFc1a1CIQFHUuQmd4oZRGfq9QLqOd6aVqcHKAqs6mOhOYPdIKYh8bv53a
YNG57m13ecuzh1EGvM+Npvgh9o8TUMHFspKYgwcquSIRGuYCXKRdoyenZumqf1BPrMuDsaMEFAxs
wO+47/jyrixYo9TUUFND9BYostNPthdDixAHJv55dHk9CpyIEO951XmM8H1tjt8KK0hHKYRrlQWE
vVIkRG5RyCl/5NsXt3W0LBfF6eNJSaPgGd5rHnfIz0dQLEci+FF+lN1mDgj8zdF/zAocu00+RohS
ka+ZZjL3MqUn092KRL401vIbGtjAmlw5X3kBMcC0DjDFNjH4Swge+sK9Pw1msvX5OJTy5QdVXbo6
krAaWwB97AzOxKZiqVD8CJEpWN8qlfdvfjeoZraTJyQ8Op9fwE4fgW0Y/wiHRnwtBis+TuAUqGB0
wHkD/JFiYEWGLggcGcjrKr6qmOp9V+Ekgw0mZyqM9SoTSl9DhGDGTtH31v0sIu6m7KZSRBlQALfN
Us6JxMXTt3h8o0uE9z6+dtjPBD+RtBPmwYGNalOkyu22zDuX/s9uuyF3RmBcxLl2Rbg1AhFEvbc1
tJkPYLaCgReEFjKd6NzumsH8Rkuzg0QV+Tkge3Ft+n2Js+zOEVnR8R5Tac9/Ogkvh1Rv/KN4ojhw
5ZsSJxoFp/33mL9dON0Vzclgm+BURWfRraZWkbyKriH/xDEorcVKo9N2qqbnFGQATdC/WKmPUN+H
zubE/I57PKk0f6Y/gZ9roo2POGX9XsF8OPgQVOBV7jvN0+IjH0ZIB0xqBeK3/lGCP2LmRZYBDNaI
q/KdknW2SMz4ERZocp7pBxSNT++KHfFp7E5R7nXkUeMgpsQGpJdBC6EMYbrnneGbwkFRFqM0yoY/
iM+CTXOs6K1xXfd8hNc+yktJrMs0v9uvYYYEbi3C4k12eIRDAJu2Hp7hY0TwTPH1FLntLKoZCO4K
RBGxZqlVAjogE8QSH+TNbW8nDVylcbifIL7RE7uoq6/hDYuihML0KJUynebja4AmljVPuQYa2a1x
7WQt0uCWIOV1n2XHj1yi29iAyNW+gbCjr7tkOL3FtetpOzCDJ1wyB6B6MmIF50wNcQnfZppHz0J4
rwkaP0fHQtpRIl9ztGsTTnzpZiBTp2ionXnMLddjwqSb+R8UVK8hqK6wY+FicTKB8Ta0U2S4+wPf
WU9baEK+FDovhUsJZf63I/XiJauwH1vxnGXnHFEisvq3pmECPaK+eGtpx+TM23g77Eovi+Sindtc
ejRznpWZwdxenXRGlCH4x8v4VOuzGK3SIV+rIa+6/3VPhaCvEDqrHD+1slyIG3almguTb+tow2B4
55tJ0ReYOWQkIJ+NChZUtTU+oNhw47F00PfymZ02HXG1AcDBxasaCHashhz0Totjkf9O2GqwHRvE
CMHzqRvz/daokjibhgaMqpYVh1fG25WVNpfccHB9pPfUebb2wqexxIHqiZmcT6/xCKTToGcVQHHM
FuhnSyK50uNi72NDyqcAzq7o+mcoMU+pq8gREGztohrcvi3RZSif4uo7NDVSjwQG41dmEXGWUD4d
CrZwJ7YV2iB23Xbv6f3gweGG8rIYwCIfTqy6hbOpYOKp3VX6W5l7xTGtsIdAKC9ukQV6aRimOdtO
VOGWEYEMFU/aV/ZRQi39bZ4XBKinWM9lrhN0uEBbBblElA6Lacsj5JCEX38iLdZsjQ1I+uh+Oeqj
NGtBYaKnAUxQppOsrAQKfX0WEgRr5eaYThos+qoLnVefmOx+McGTJBXk5HKMhWuoBdFZtMXrgpnn
U+1M8dkzWdYGKGkReMZa250nCkg3uUVNOsoedrld3qb/hwfVx7ntwa68ZLKY4BAa9JxrxrbXHHaX
PDE2D/CeAAp3BGQoyeVF8Tdfrygb114fnEST/uF/ZEoDriMIOkbMRI1DCtzZjLo6gM5lnYV36pzg
c7BLVpFt1hsK173Knv6ccezL6o6ZkOOGU/AmtzYO2b+OW1JjjhjaGinv7kcHq7pyUMHaYa0t+Lz6
qio1M50QyiQ73RrZz5gfo0Tw9WyIXhPy6AggaiP6aYKockzW8QHGu+Kscpnm2Mc7bbLnYz4V0Hz9
IH4ifvoCdGHvnnjNCt3jhLl8iQlZuxiX7bisEoB3Bt0aZJyHx0UE5xuiNDBhzlcL6IMMWYZ8/CIs
XgB5V3+oDpumQP0mLrrfIxJ/xH/9VHMQqgrDvYN2e/WTyBkMkzfGC/gvP1jb46Nugnelfue9uGJk
ITEHoBUuICaxZg1v7w6ylYjhprr0XYgrgbNO+V3rhVF3vpE82YR0STuSVU/wESfyCCIK8z0dpJmM
0GGzNg8pmkWGvRJMLzEGeVCrOZgpBG2bsnqsiL3sI4fL3VxA7n02M/I7CwOgimmxFDF5LZDtZWZA
MUuf8SLqC87ELRYfW6czSPqWAwDjPtrwpMyTgo/3VXgLSZpMWH9miIuZ0RPfSz/PkF5Oc39JGPJT
aGhG/ePE7HTtYlE+ZGu0UcuakJbb3EZLdFQz7PXxzO+d4fRO1ymYJolK29KspGEpwBmTo94NG0c0
JGSdS7pHhjYrshafG9VNsv//zgrjuc0cqlqUr3gxhWUf3T+BmOKv2dyLeJLw80bzWWb0is8AS3BU
Ka/1WTG/B0mC/nnkpTEecxITru0Ry5JQe6H/gVOeo8c1VKPkJfEhGda4JQ0x+uxDdZETsU3iT22M
kRXA/ITq952wINS9YF17aIZlrvjojGyVx8/apFF/oAHcLOtKT+32PaonyS4oX8wfQrCwevf0Fg/W
vl0EBKTc7bANr3vh9rRCibRxJ9n35/l66af3uBHJ16FiepSG88y9FxHed+aX0V0PU3x+adKiePRG
8unEa5yLfrGtJ08qiObkKf93m2JkOai1aSXWVOEmqB4cWunPssu6dxQUdcLHNubKajlz7XQxiv8a
L11ZWCgFO6SWJnzU14J+z9Oczmpj+UyhO1ELrzDbU3/GPIwkGFOpuyvnPYHaNooyTEp0KCYOZl/m
evvV72niLfNhjAHbm9JOM3I+P7eSe+zn/qJln/Z3++DhN/eeCopJVkU3ryok033Z8LjLOq9cLhHs
rRGk+LGTLfsyVshWpaE9uZATTYAiwfRUKgQKGWLe3G0j7PvvXxYGDTsswIO2OppbyyIbukNuuXaZ
yZjM6FW1lKeFnSApJQeK26OZE7kevzk0e2RQ84ojd2TxER6AwabvQJbSrZ1Eq9K/9fSwwYTx2Dzz
BlXCiRWo3b/bwuTay12WzE25u+9f04akZDxsxl5eDAxkGmj0lEVsx3u4xGoED/vge4xg+/akr9fo
x5w/m8NwdKsAKBa96DlH/Ce8zVbp4yiAk5FvnYG8tU78ND4sbUJQaO6dG+iXCYhKKMt4+6Sihqk6
heYGGQ7GWq3Jx8H09g7NHQ2WwxtIsIgIAyHwW99ggCZ7GRmQ2NXRjlBG2zMpVD1LDid0y01Y707L
nKh33So9Y5SnS4zxS4gegIsb2bsHgTx/mF9JG2+8bM190PMRre+q9CFD/w7/kVXtkPvzJeFUbqdL
3c5sFi1jWzpzMnN9gtcWUN55E+l5qYKK8Dfn0AZiuIb4ZRc930aginY62iVeg9IOMY3pZ+D++LzF
EtKvhhqeCRPCTh7P0EE94PHZDhQ6k5jkv3pi6NezWL4SV1ziJDgwU1pCapNWmhVboDKNqHAsQs/x
XdeofgKgzd98on/H7VdH2+yPT3yNYq4SNjT0sqEM2z9h+jSKyHclW9cfHMljg/YjIb2/JtokE1XA
LqjHMKdohTQ8Vg9qO8Nhz4kdOZsSF6HKT4A2rrN7V4rzzs61tgK0U+AD+aqQL49DA5qGj0ymW03F
9DZlw2aUHsbZPD3YvFSf8l/PJD6/D19QfxSUQPHhhlceMh02YeHb5wnrmNI/e+uuCCvCOv+Ig+Ei
448gDvGgmzdUGTyrZflrG6OHhqOmujboN0aDjD6rH0opMzYUyeUMzl6V9t4Q+pi8+ZpZ2bosP2Wz
YkTk6jXv5fwk2GdNSyKlm5v+9+un/PwGHZDitoT6o0EX7GrRthfBJAW1KNn1le5jfYt0ocLo0zWk
BIWSt4TyoPkbO/8Ewi5huoktsvo0sL2c5EO4/EdVFJMX2xUbNmlxIyP2s0tTPUfOXxVPvfTVD6rB
M5R2KFmhpI0PavrlVMkk9bDHY4VxYfoCFLwRg869QhohqmbybGlnqg50JDTAO5nzmH+4Q3v6T/2A
EtoAhqGumsbIMAU27DH2rHzDPqOzeaKXO+JoNxRy8buM7Pu2ID7HWwxgVQ1iscja6gPNifBEwd3B
hbVpu49tddplw0Nd3z0qP9O2rsaj4FAw+xSpZUdJWm/pwkr7yx/rD0LMFl2nZ3zU/5Tg0xXkr2al
eWIQmISdVsKHTEDql+vR/RYbT/T44UE3c7fhk273XJ7wHuFfbRGhwxF/6jMqelG2m+TK3jdrDo9D
ABXiYPVfR0XUyq675++V4QMtXnpM+BM2OCIfWU2iBmXoBF57ddWmcegIXdFmTOOVQ7BdVX2jRwlb
hHM4VuwdseKVg+tJUCDcw79/B7lnYQV7UsVXnND3cYXMeqc6LZTwhEbTcrMgCgYEw+s9XuBUS9BE
uD+Fe94kKeZbkdKc4S+JifL2m4yiRT5i3QTiDpIl3wDj3sYbrUEfxDs8Cug3jX4IWxNEh5O5isTq
IguRqSxwvDjaVykJ07SulNe6p4gliYtxfuJS4+mCrRAHXju3IxoTB9CLMOGPQeRCbZfoVJW9oPwT
k4OpE/B9k28Hx45jAHhR5fyWWwz1g7oO/KwSJLTGQfYuc4LVgWNp4ZdRowodkBsgyYR7Z+qoC3Y0
md9c/QT/3XoPrPgXCNv4eZGCZPpp0FweqD+sjvHLckWMZq5ofJasXlBCgq5l00E0kMve7wKOXuW9
f0pEUhRClIkuZ1EJjW9m9PapFSlavdkMMjJJlO3JUD4swhQRYLUTHXdwIk9XQ3HsJm8KvOVKa8QX
gQUFEcuVW1XgxDedlYcBncqY3CGN8mnFNmVl3GlMapFc+ZXbzyGwxPT7AmgauGY+/WEImsfi3ojD
Jikofr8EJ40ebODKmV+I8vhRpQiRPvkUyGJ0TXE+QA/s4QgvQV+OHpZRUqvOmM9uJfIWLJmoR1L4
TX3OCn57WnJdzI6HLQ75bPCFI5Uc/O2MoalTp6spAgiN2D2OxsNyaxfgcY2LvbumrLluPK0fVTY9
PFf9N8U12y+daAz+2ff7loCzMuOQe36ei5zDkOHCBkSJ2B1oRgWw/zmBdJq4GxM+KASfkE1hKpm5
a9NYZuLVwiC+sbEitjUTcmY67bi0M4cemU9GdYtD0E3c3pJGDwNtIMUpvl6loCCL677zV+7KFm5G
yMo20+yLT89tHDHPJ8Mv5t+2HOhSIxGimdh90a8PZqYUbNC1j7omuZARPWZh9MHVqGoWbH6X8mC+
KWPfvmMt2+CSky8mLbVCCs9jOpDrM6BLFiwD9l5uLKKR3qLk2K3++dtop8a8KI/2WiZsYnfLeJPK
iH+SWJoxmHx/FIdec0ts+RVI7fAwSxIlpd28o1HFqQPVqZFG+gTHU/t0/KkSY2JOdrGO5FW6kEaL
qbiEELA/hgAPVxMHXxSDJgm/HGw1gbQk3IW9/nY858Zrl696niuTnexA1gjkwm+EOGAcTa/J4VHr
MoTCf4rw9mV2jYW7W0T287ijWhJzF7iCMVYTJu2OkiS2hpAiiS+IIFXH+RrHr/XiG1O5EcsyO676
CSXPoEIlKzo2G1xd+BkbpVQr9QKtAs665wwFh3AQjfElNHfFj1RW4rV1VzbuD0wa0J7VFVgTBdpZ
8vme9eZMDl0I+59JctEq5knlEqWmTPt3nzOSNySjz8DhgFU5U/aNMCsgBhBGWSMG1XP2UvD3g/Br
ZdI6DflKOCXt0JoEpIAQosL+OWE0bNbszyxSwz5aX28a6XNpTxvbe8R++k1BzEDMUCYYcba/iGUm
xXwgF8J+CzISJYEokS3BH2xCg4npaUE0hBwMPJkKUwJuMF+wNFhzJ9p8TEbIaELJEdzgzcAGdVIw
UaX36c+NRxEaoNU0eRy5gw/4VPTD8Q+RLh+maMB/zXJ6+v2GdtGMm5AIzcucBL/thxN4E21jAf+I
0teKIHIU5xmYDwjhl6v/M56VLYddjJwCQ2ltl/jbeJTIuAW5PUTEN7bjWPb/BcuFdCs8Ut/GF1LJ
sWrh/+Frk+xXOzBgW1Xekox72thllxkQgam3M7jXm293AWHXW1d+4Zz2LeUz7qmt9JzKYbbCNu9A
bW5stllDHtGLEcH9KSEyw/9UR7EUKua7rP7xcRPHbZiEeRxEZG56aZwzJu2yXm1R2jZmidwlG5Cw
8d0yhZG9YsbAz0N7Azfov3VF10agSl9c4kKKCFMgjcG4nlKsLIwxS79MzpO0iTcIc9ApkmaJobGO
1qaxucSR38UGkRTDlNiOFGh2wmjq375FAEkIPFDPiUdsQXMcGhG+M5a5rmCJmrRynCOduvGA2QVD
qnmcYncm5/et7w6sVNBAG/K/D0LZDN7zm5Tw4zQZSHr4zeQo4MWO3RkaP/iRpcgGbDKalaV6edoG
JC4GGcgmCe/gkAXz+yE1PtAQuaoaoHp8dl8uDFOlU8hOgbk+bQ4nYoALQgKWS7Qnzo0Bb+ZPDee5
rZbSOITrvpzpnvd3Z2Rvq/k5SPBVviO214nrMAbRZif6sT4rd+M8Cn94OuFJbtch1dZBu6nOIchd
FgMrjx+Y3NkKVxmafC+AU3EHpu+M2c+InPP3sMheLF/TJsipQ8fZG6p21xPJGKsErSsvKHCA4Qpc
HuHzj3celJ8pLofhnUV88hdyZ+pJecMi/+Q/ZtHQZn8+7QGtrovvIxitBpVX4YaOTMeXvVCuo6tn
yF3OW58JZw4v4jG8jtcxGtrREH0Cbaw5yHAJteDzfp1DhpUBZRmLU7jd40o4W6kvR26Il8WuVC3q
F3i1RmCwI7+gTBYge8iLwH4dWI/UeTmSOkGyQT6EECL86eA1/oJpsy+vrQKWkkAu4tKRJ5n1QQMV
myKKLjFh8DyhYEDza3W3g89cPZVbK/DiGp97aGawcgUBG5pDwgZT3T7gtS2saqg/2okUq95bHLnW
udrmkABQAkJr11pAF9YNlCGxPAUamkUTR6kXMoFhSK07J3PwMOP123hhOekYNlg5raKgtelWaiXO
ipOHXgswBmU0D6KuXaDNFx/jGiOkk2CdkniJiVO/X8N7sY7Qaj2XAYo4rSNYnRh0bkf6iESADCUD
DUwCkgTllTcfBK8bNJemgu7kN1L8VtpVsbWG93cPnIoqf8zRt0bTVThyZ3R3tPGv8oBCEaytJ3K1
N+Qsxz7sD6nLF01pLPY//cwmJuHxJAZVwoRGHFqRzHHRjbG8LwQvOlk0/UNdZF8RaO2SsHpFghZG
feMAmfnQv9M87MBeg+Dh3aVmO8L+hIKxOt1afUNBdlyocMWHHpcxnKFGTjE+yf0VMJigUOOkLdBb
7sL6bOJ7Yfa1gsNGvLHKMzsAgQl96gs79I3o0x45J7nDBvbEd98RXM4SKcDEtmXc+7u7hSVyIQKY
/U7DdJn4SnfPjOFOJXQm/bw85lSnTHv7TG+xiQp0zmXfh80cxZToj6VH3K8+5NfMgxumnhEV8KzO
fbN3VIOysIcqbxP1wljLzDsW9QCL/DVQViCVUtt6ORHMdlHLKQMTGd00rrr5TGQtYly3wZQqNd4H
ZfZla9TynIFSEQ/B5i/4tLncwtOe0ukMhG/zlW0jhtz2VOWnVCCCa8MT6V9IKHav/NhVKX/d8Nxs
h1DBIsUSytFpEHhdet5QzY0Ax/+1drIHfAU3E0SkV4lkl5c7FjVSnIMjU+bAVd66cD3pCCATHap6
GpBJrPg/5YAXjfvdKFGCgLpPc9MeblOmsILVaXW1iQTs4E6vPT7Gr1GCfNxTlAD6vJ4r92RyXUUw
nJ2wPyg07+8dqx4HwpdMNo0HB3t5cE8bjGoqEmH7Zl7MjZm4b8WpxX3JprQ5mLSngR7wnWJbNG6Z
qFD+7kxq24/q2NtEpa3faHb4XfMaWm+f7POiKA80XlBd5btInVY7nabZex2ABuriZgZ0IxLX48Af
/wAVP/JVmZWs64K2PFecqAuFq+GVHBZL/LwgiQaTsgcKpFZ3OwtOFT4Ub1CmjxYuPVkzZeoErQKX
JQ3dF73MdkNp8nwK9KpeUw+2ija/aVR3zQ/5ncFL0OP6EhN1CcjNCj6LGjWMzwBUjy+M01CUXcq1
5XC8byd73fUS7WxmApcJOnCfp78V7QOKnJwHWKoHcQvcJDXVr57yIiHjDmQg8tgQubvn027Lqm74
IVRPhixdXshPCQ/Wtks4klKqArxIdPK4SWbjBYJnWMe81tqsDMs3rU38MqErUry0bWxh4WO23GPq
tYmJ66my68g9yh/aLCXOOOZnGlXCHGuhu/LiHZIh9bOk4bVcF8DyvZrdF6f4vshBOBrOZ7CPkyWZ
5+kz14UE9zHs5amJOLHA3RzPqYVIMDb5aTuDln4MEQ55GnbilnoS5lXhUT7xY1n9Cnj5K1gRikbO
oz5r2BZp7DjyGhqzNlpv87awdWYEPTT/8670vZHKlpah1hF+U3HHOgoBJYPFlhpwKoNOnapvzSQd
gfwqKvPLozJQSJ1V+imvlRWOG3BoMhqfHk9u7960gfkgrH3V4d2YB3+y61roSOJrf+XL4t92SEOc
qiQAlwNWtia4mnVsBl3X8YXcjgIRGr0ZiLM8kGrqtC2gaqultThjoj4RoxDKGefx2yQquCy2c1cy
K9ft4AQShcvHC66jf82sGaX/sQWIcXdLfpMRq2Hc9TdPDj+2h6Fssx+W2s7kyaH4kEUjQXe+FRGN
cousXaRRris+UweYel3h8yQ0fQcD3RuJ5MY21xOcDsFRhaZlvNljWv5B8xZBd+6eG/mj50VSd/fJ
EXrCVFsb/o9BJPKpc/ZbVAVlWnXkTCjeIZw9sw0MXTI/BGV2WoAKpkUTS/NLTZ4N5bLDRukeRtsw
KSUuMIloR0fsGDLTccferELOPkLB05en82zBQ8MSbca+O7Z0yNHKK/NnEis2XUJerrtDdTyYJYfh
pKW3aOWFwcLib90lng9NgJA/OGSR2mgRR//qoiVAfZKhJC+GkOjEdyeiYzuPeCiYI6oA2/HlUuK1
AXuB6oMwsIiSuJvbcp3N3O/kyavT//34FsOD9fWwdKhp84HbdXp+2mfid5qg5OkOJ+s3lMSLCtxL
n58aPT5e5q0e/yr+EHj5sbqtTiq6MtRcMhvlshGzHOlF0NrFC3ce2U5TTSpF2LCaNuftCWK5CjKW
+lAS6x/sRUZL3aQJ9+a6LR72SqpOCq/VxuP0WjvyY3LxFyuXYrr1ae2fspqg57eDV+A64QapIU6S
n9oKLAYwx1Hl3H30dNhmUB7jM4bHFu4Vs8x89re7MIn3/itbV+SpXeTXU6vFRJIM7nUqHpV96t/M
pCZ2ULZ5XGZrteKDlfh+KC4h5O+fg3m9ofue+GSTHTRLrRFjcrztfdJzvWAmoe6Dk6P/VX9bwpyw
NR1YMFPP+hZ8OweYFvy97m7ybVsbSn83GLKUNhpqoNPLRG+QTHeV/wNdzdRFodX2eNs1OixYfh+l
39ZGNfDV49VDEsixTQRGeV1t1j4SDEX/4Trpy3W8jkLiaH5NHKDpfW35VxzzCoTont1cMeEd30ux
Rf0fUTLMNLdwevX2yx6Te7aMQGg2idYiHDzPlQ65k1nUMZHeDhYbHXS4hqR8s3BcWhtJaggXQL64
TlQG0HZ+hkfmw3JqTv0iWgOaFsXlKbMSf6DOyuO4XvQTgWZqER+yq+NSf47AL3MGIX8ZfNtLgCct
QRQwISLrRZIaTBlDsGljmEC8ouRy4Dg1kHaegbqZN+N/76ehignggIGEQPm/wswVKAY8njkBeNeh
h2mWVptChm3ib2FjXQGek+JFB8NC+gsivv3hPV9gEF0A+yR76M+/OZIs7VEpaftQy8tyj+rIGCJJ
I2+rKuuH+/WLZvuMLWh8HtxM3bwVbL3Tv1RLOWrG18gKrcEjFVJGDrLYwDHoEp1hS/hSphnBeMGW
yRq1SYIweP3ODeRfEje9oYpUnOd8WWdELjC28YNtmvQZg1jiFtx1pNyPDeLVMpmkc9SfdOs1Mx/o
lyaqYx/unoIifghj8tbQmC+addcS6VyMSsvCd/4GztFttklaeT79gp56vBOaDpK1Toj6PEnUB82j
bnc04M55sJDRBTC4LIggE2Q0cFY2/hYZizFxtuG9JNYiXoK22uuJ9XMfL32s4uL8Q3kDaTIUooGG
c7OUi6C7+rXeP3YsLeNnCQ/FHkP2zZg6z1ydWJrJXORH5Ff7iw/BqagdbBYHjVzN/LRVjZRKJcNx
/QKpxOYq/QWvHuhaVISr+ksRgsN8VzQIdCB1/3C7ndyD6EEe5EgoIlXU+q4LurUN3sVbna5xyTJf
X371ZtVzCSIyxuJF5OKxlawDCE6F1C+5S02t4lqzsq4R6gsVxiYEzsTHWA6V6w0F/HngqaGmOmUF
go4ZGXVxaWw4aJjHPk4raf/pTayxPI3ehbDL/PF6FHTscFt2ymZyM5XXbwcK3URM280vJuKy002B
/ffn1uWoEiOltDVK/wB7oS5Q8GW0nH1LLD7WRbYUCgJUUkAtpv7o5w017AqXZXiijBlQULg8KvJn
AJAhUuW+SPwoyqaRjY89DH+zztk8hRgmmLyQvdjDhS494rY8X20ud9gJyzQo6aSPaEbh1ZdA7uZg
6aN+vp4euiU7YHUS5xSmi8bcB7WwjWnwkthVW++Qog8prNsoo25UtewgNg26Ii4wGR6c+QW+uFKq
/7/4jgQZktVTf/IY+rWGmMUwhVT4pHGIhDaQJY1FMPWudoxORgL5Xs25jeUqJHY361iJdOKtaifn
788XvoO2dnhuHwUxzTUJHnmPdRs8K2gmEkkPOuWh/DnNKoRq7AZkurlLbm4vjoNd0iV7Y4Kvbdun
NLLiAOvey+e5K3oLbX47NN9aJ33to+Gq8xDGzQn7Mm3JnH5n9sqOh3say9m/P6eXEHyJ8D/FoEgl
288U4DDr2N+2yaS3cZyYmR0HEALMfTuMlFH9lVeInpRm0VNAuZonSEAbTN693uF3+otyqZnzwahX
VomzBJnOsxCiyDg+QcKhQg0CqaMWRiqDzjdwkZpT/hLPVdWKAYlpSGqc5/om5RnaFg355LtbnEB/
dF9KDTjl1y2rgd7UNMGbhhLpH5kBFVEd2P6Nr3WZCXJj2MPuYr5rFzydhDXlDB8kU8xp0hal/q9h
zl4T2frl8XkeiFioM+EBASa7jupMtZaXnv657vs5PBGc94YMhNlXdkbCLYo3/CWndvVad66TCdgn
BpNEhKr49Pax/2jjQzRElLDLxe0kIVa8c1D8idwdpvRDRR3zQ4VU9Sjc+pvFcqV1TtXQZzeeNmmb
hp5OV9aX61ymhgskW1lanjNyaJW78DkidH5Wxv/buTTSNrvkcSDOmQPnJjjN9x44GLFJNNMTDCaC
J/9WigCUNZzqGYHc8QeEZZ2/eoxVa0VrdHjjF0Dx/QdaK2lGEa/w/6Mpf3uCMuQ08D4eTpxXfP7X
mYDxtJ2f2Ok8d+ip0pZZoDgh3ppILMNo6otkLQlJRCkuVBugtSMBx3KJOMrwzzOQcaYFddHXUat/
wdO4K6fLhgd9TnEEhNWb9wPM/hoEOWmUwB9+35xS1nSjEEYOYFv47x9G9y5l2kxAfuX4VvtuFr24
1UTCb37FI1ZDhXZhnZgQQ6Kx03NHNxC7oC5dZJimv+wMroxGsz29DmtUeUieAdNjYnAmVv6kv0uO
pRUiZ/KQJCNU2SpRsINjkFt09tDgExl0OEF3yTLQQZA8s5R813Y7bqLhVZE2GP5p3CQ29XeiMQSd
21E7g2MzSkCjFFzMF8Qjo52eiuO/gqA9JugPVy8EqH/NsV+rExnCxvlzYQXCVAKhkLtudyQS3R6t
1d83mqoWQsIb9BP5jTt5z2HoSn3+dGjLdHz5X+TY7HreS7C9k/EfnPWF5bJfYiD6Hkyn1k4ceGHW
wXw+4tqSUtNM6xI3KxZmHF7nGqI+P4Wy8x9Le5td6LPqP90aJYcuD04UbKxg5EhR49TGJ4+Yi1c6
iBvnu1R84OcP/ATJOsIBtHlhQdPbMGfbQhcmoE/XzTJJYMiJ1OUChFf+KAxnwE2Remt5cy99Y3Or
MWQpoCHqlXwhLyVrFpeBeoJHoNl1jP9QMavUlcz0Q8W5gHZ0gJ4fNYI1f8xOOXNOxajsroVAF2jy
CSYt7yo8mceQnYx61ZNA3uFQVC1c/P3VxA3gHasYNumQEjFfCxmdsI1j78UTeorojPlbuSl8BQqb
8cHRJLtMykRzdR5LDy2v+Qvry7k9HC/J1AxE5aWf1Dk1Vsf7tS6ViS/ttby+0BvgxJYyosim6r8y
c26TsO2CqcRe8vNFB1xuyYLXM8NO3bc8btsq2Vj7IQnodzlKRxlXCDzxMI/sro3PzjJg2dFfRZRr
0hABeKzGLDWkqKDFeShLtIf6sMNaC7ba0Gd3/sHqHuQpCdeTjmoIxHroRys7ubAQl8TpKk+oa7fH
X/jcjL2DyZTPJA/4Pc9obwCG75H8KJNttgcslUzb1QNhKv6lnKtw6mRQVuE0qapbWdroFjHSYaY8
nABzNYp1J04ekTX9cV6vW2X+IPQQEHJJ+gArD2XF13sNR1kw20E8AQAux9ENEmk1NdVdY9ilyJ2B
zXxFy1iYT6X2P9slO0RYu1QBA9wfwcgAG1R6wBrI0/PZo5h5PCXS3q25cLHm/3Stb9cu6b7VrVDe
VNuCq36Pwr/evM3uMPE+Q8aKv5XBYnuCKxroNxQzoPRoXnQBjDqarAPtCvirNaqNX7aal9UaS+VB
D+XqAvcWDi20IhBNyLM7zeNTOes88modDBfHAFPA25Cfj2WUO/qqnby/b65V4Q3sIZOWpj/PdUl8
uFx5rjtFVu3FxHiP3/KcalN1pWKwfIgl04PLEUtqMn+yoF3MX0QoSvnsJY+XwA++MYH3FVavT965
FuRe92YN/C1Fn1J9W5UVvuparkKh9sDaTTSJb5LeE49zRU172leHHSdYoyP6ra1MpbG/G4lwJws5
6AmDo1IgZeYw7tTlXDoNmbFuOXGIpg4lu57P9y3buQeKdOF+RxRrPSO6SfTnH183NRPHgK7pJGor
on2vhWNmicQHkpYb/v84MFcmDsuzUXrT7DoilItCSaRSY5+Ql8vJ8f0H1sY5o/AL1Toz4LLiNRPf
r4oiN818ryIaWo9Rhzwn59p2q1/MgrHa5zZxOIN2pTvyC/rpdyh0oUqWyb7sl0rsEe0PsBO+9GQa
US/qj2anDNMXImRhfk7G8fBG4oFnLJhALs9AAeOhcNjnuyntD5LQ1nAzf69K+SxgSt8MQzOkth8+
AZ9oAGww/6K1BCO9Kd+LQ8ZpAszwUdMmoy6IeGjURyKnvTK+Jc6cJ0maJzC6IgvmcQO2tl5qlwG2
4f//RN4VQ6pUvz9nW5xkS99XbaJ5hyhxxip5SWpJMNQzQ16ep55cvHCTZDAo8MAIcZfDENH72Us2
5zYnRQ4LU5FE/TcrXELJHf/ZQG3f1VDSqkBTXID8q8afSAHEbca2xbvNvK555RUmrpcGgfNZCf5e
HCCGyRTpS9x+Ol5JNLKXeVFHJZ1+CgiJaAbNhqIeozMeErw4dalqAHVx5Ika1AgHvMdPndaOVHU8
VLKsQ/gfyNjtCEECy1l1mdmj/p8Kk7v14cSei+0y5sBiVNa5ZXFc3mW1FJd4Khh6Sc05G2KYRvkz
UBcwezxDDLQ/M3NdAF16ySfWXAzH2Br+IgX/KfdZjhn20riwnyVPHkB6EU3OGZhjqgQxVTbRtHfL
tg6qx3EAnud00GLYcvG1Oqv0oPxoLB6nKR9juKNLUoFwUoiab93e1pFO33z5ceIoFT66bF515UFE
/HEexYBFVNW9BGpO9NmvrtpmvuHAjNZSgTTbotdRMdcYKY1nmCxooPufj9Cl4vDQmMvLYO1znjwh
f9KndwgMOFFwCD654pTIXKcVRL1nMksl9X38wLr3dlMKMOn0NKPLyCMDp3luNxt5YmBPiP2ajiUK
XCPsGt7GXA42+Q8YjkA9h0lRkyUicuI5v3SuY8ftlWDe++zEK0M4xaEAjt1mBYetyUwvsFC6U1i0
JLmZTcuRJFLNaUnb1hWYhjPb4msJOrb6IgwcuYMUGrfzivBl4/MxZDTOuwLCprvdO0SmN3I8bpCR
GL4N9yOeXPva8aeGSGW6VJrKCl4psZAmIZtQvxWwl1t5895MRV3JvTN8PNo+j9fsHS8++6fIg29L
PL1eZqEYD6q631mD/EH5fYeV9BLCBKIFZ3MSSVcGV58lGkzsiNqv+Wk3uftxXL1I8/q8wxaIdKqq
ncAPAx3RUPbxC7v11i6t72ReHq4nFctFB6ANAKqEIb6494Ltk9SrveDv34KFceoJroeSzwdL/xOw
SSUZ6xZ7lCCS5HmyPaXXA70/zbU7cYP3nKe5tBiPOMUB9z944ihsfggK0tA0oIw6+HHMXU7As2/2
deJ/4nvPK7eeFfdGUBz2GxdRO3G71S9cXBxA+KegxhxV14I5R9f5fQjtaOyurpWPN4vZZSiwUgS6
zS+reHIHTbXH8ah7jyUUnMEAz9S0rNmpNUSv/V/innE16UNCk3rofVM26FoyLcO37+p8jru+7APf
LJDEKT4eYh7+5vP5itnsi0N1eXNs2f6q/GQpeS8pwnDWKPE9ijkEKhH60U/HV+HJFoVKm9wiZxX5
ZROVEwT6cryiczi85X+xlz1qaC9XqkeKblooasbpYJyCq0sSW3ws1DMJudQgFinJhDVAjmj+qDk0
SZWVTFxg/9ZplzyyTXanRk2fzvWouYyMdJ5Z8j2I59qAMI5yL0x/uBeUay8Jv9c8APJISEuUIKA/
15IP7wlfNKXBbeDT8+vcJNckbZabv5SWqWbbXVgE5NgUrYJXBvvZ28rtwEoKLqvhMQnfZSCfSSTt
IPWIW7HstxWJ9q4Fsssem320tGFTVtaSC9rmegpJ2o41sY9U6gEwH/qoglX7Jr21XdYLe5LuCg+O
8yUxoP2/yWkRnjPItZLvNRcpKMqf3fKnz0KDx8SgatztgBRn/azaLlpgcVzNSOM5sBgIKPs2g4Tg
65XEOi6xraGrsc6gYRTzT3KZFf29tfNMQlLd8v0Ca/4ag1b2TmCiUXwPMdoT/S6aASMLTxCBpBop
+77y3ETiT0hBkpp1fVrowAS+Ah1lz57fAVqclKxphx1ByVh3Pw5Lx9z1jx9UUbCKvKgpiMhwt3Ol
PeZx+RCvZTn1eWDYVffM4V6IspeWF9sUmB35pzio8cLASd6s5gyzVE0A6XMiVm1TCf60jBTyD0+2
9Ra53BWSuuFoYikcuGnRNHWCR02KdpPnwJDrvs3c2eYfCFM61VRMAH9JfMveFIJ+WNeYofIEtHkn
zUmCrDQiBBQ6lmQUVR2YbhUEjGHlV8VMeacHJnVrN3NEju+osbwgNJq9vY1LWs8yZOY0sS2HCfTg
77RojsxMZ3SBoSvcFohcNs2LrMrggP0RK2jtMpyd4VRzEZzL19rUKvzA/E5BoYYkUhIBLxBNvd+2
hSXmeAoizZXyxV4jQWIxGa5UB1W41KYZt9F0H6HTC7LsI6KIwvT3WNqM5vtL2sxQJJi/v1euzYQ5
AcgEXahX7YzbVGAEwOJCOK90GoDiMLtiJCJ2eMfCuiQnLm40aZoOGExIv2+14m0UK8wl0oIJJKkj
HwpXT96MSXcpLK11wxM/15qbNNCjvHg9nT8IBQPLWEQxRElFdbi3r/JUzPfUTdWIJB86Xvr5RlT4
6O8QCKN1mjeTNUu+UzAC7cmY6tv59VEBGbJCHj3n+A17EgztW0ZAb492xtAgzjPuWLdRnsyWJ5yx
jw2W4z4baFHtGaLcxmKStSvhRbEP5JXBtUN48ZGTRTpc2LzN1fbsv99PUzZc3RmgU2ij0zWqZm93
A1vXuj4MZb+a3pqSQP/Qfw75CDiRKQH3t8/8wpSjw8BAjvJuisLetOl57WM4kREh+swxYl8Fy6bY
K8CJR4h45BsQQ7nhhndfDR+yvhQXCz3enmiOXS4+mZIDdz9L5YFSO3E0XSphBu7Lyr1FGRa3rPSw
WXx7SV23LTU5H5V8R2kyVDm2psHOSibsvdj+SvKA+cMKnNyv+iRJdcmEkhwwPZo0tW1yGd0Dri3X
1H/ELj9GD6HXWlodlCyA+naYnfI6RJoIJNspF++iYT2xuJF0jU3I2QcuZu9crYEtuIdiME1KjnHH
JvAeTa3VbR9+s5mkYo2NKqLUP0vz+ZA5KdG2DFuA71agr0dDJwtDX/3RYOtXOKolhAs7tbw9KCNV
PFMKVribE7ve2zkqwG9owk+M8yFRrFrpEHZnpwEW3JS/P/iaGUxyI05kUDZPZJzUYu7rdHIkKhTW
C21j69cOy5E5w4kMd2mbVEAIDclI//0eOlD3nBSrOUQDv9YTbemiaWDVlKvUC2dUTsLg240buvIZ
grm0wl31O58Zx+Kh4lj281bo/o4Vihj1JmPzNGIgfrCr6jduXysT1NhJNUYQR2ek5dIZXwy9ss7D
fYA9gtNGGjIKISrd6ttCCWzXG981pT0ZNIo8IiLWJC2mMuqDAIm9GgA69lPGddOXgVKhMjjI5tbJ
xeA+G4UbtVvbG/2LPJ+KOqpoD/bfl5Voor3b+T8UiDPSQlE0HUitM1lIeNYCeL/XEEBN8MFwORzr
D9XJ1J1qXX1OLJqTsyoQQilHJwuPU6JZuzmff0Cx0WCqy+6x3Of3sKunAbEmqXCSuB9CGbdUuPA8
b4pjsZkeN0qqQhHlDTZolnNOghwRbtsniCAOgg7JCjDqc9eYn+Gh/56rT/wGuGrDw1Odni/IlReo
fsOkb/KbF0LgRv//BJkYthhL7DBa5JwWINV2vLLGCFXbczUmfLBAXcZMna7N0I+cFnvj4faXyz77
Xa2tMjyht/Q/NgPKOOhgdmSyF79IxJyNyWHCnTlt43SE6id/TP8DaVLHf2TLg7BXq3VxChbbtK7s
+rmGvoDNVye7WcH7K5qLYXz8dfnKqloCkgWRn73BzfKmByJjyt1J45FSAIsT2NYYM022ZxsyA6Eo
IHC3v/AcvlGg4vUQPU7zIMjAEgjVTwWy3WEt4/2DeMr6bQ2/c9H55U9+XiHDrodopkZ2g9PUP2Gh
EdbpEnyoulUbOoOgEqn41sFPvMQz94Ffsn200d62evoO987ZeBkiUBO+n/ClPRqdb278glsk/iPY
ElhIIvljze6XrrvHkDhg+D9QLzauIW/3qOB7X8ih/zTlPFbDjcV7aLm4fGqLsryZ6UMoUOSEvqSD
dCUS3PYgQPK3ST338Tw1GWufgqBcw+NfzMt3OchPH4nBCAUUy4wwaCEBsAaInQ0AnKc0zVXybEXW
QCR6gHeSLKoZTp97Uf4pGihwF2NhrzjpdPFrQKfrAXxE4/h/IR7uCUZJLUsVW1Y9h6KhflfOaky7
XZ2lOz5J1fhO3yL6PbsS+lRGVDZN7tV+z3WTW+idAqx343GbrTwqozF4X+PyjxIQXzLP/ecLK2j/
NiPrMpCZ0z3BlFk98t89zDEV6eeZazPpSu+00KWZ7VA81beR+DLee48cojOaIUxsIdnlZzSPRgYs
TRacJXhVBgtaRSBBGzTAYzX09pEfAVdyV4n9AtpbH4u3s8yvBeMX/2owR/TxRqWNO+MYPBGNaEs1
x2V2NH22M6Fu4doXLThnhjzsOlpV577cVzm9uOhRmHYr6koLqeNs+yQoyRE6gxZKGHIlYh/KdLgP
6W8DFWJ3VS46l7+pFkQYO6URlajkP8TwLKocFRawrbmMPvPnygbaYycK6aaEXhKmshXqx+qDSsyY
pTOlxJmiegWloozMC6B8S0Z87FOz5KQJP0Yq+R71e5KsfezyykJs53qgypzCbgOz7lKPe9Y1lGt8
kVz6gUbgJw8Pmn5iBVGMDoX6JPvtBHFlZsBAjp35JuWjUqrpUPQeiHKF1Gj1HySpEet7PKYXojCu
o4ukO8htUuR6jBiQPMDFUueZtOx3T6mQqCQbdN+gJ9BeqhFrJujIrDgPODVFYpfPKyM0HzbSpEw/
eBobvtEPppin6DxnWpbOd3pAc9CkAZCQvLvnQFRqkSx/a8tp3Yy9U3ICoBSfbF14/VVjSt7dkefG
Gc+uiybXjxD7DPkV+BRU0sAmefD8Yyaz4uJW+oHbN2bhI03fci9Cm0t/CI8kCa7u4uRohQuM+Spp
rOM+AflQjX5qDByWUseO9CzCSdDdQwBDFptxtscEMesHEZm36sI9X1G+fH3qSEOqvjrHnhhiorVw
o1sV0+zW0O6AOLb0p9fTPUlxm0e6Jvu80LEEjZVnuYPZVnrhsq1b2b4hqoGmTfPGJOxiVqPn4+UM
slFNzGcvz499dFP2RBqFphbtEg9OxXNotU7OizgcDtOOKOZWU4EltsqsRDETwnUh9rwQCSgJWnMu
6e0rzQXE+XabRxJ85G+1z2vnIgfKlsVyVB4ePkhk2w9h2J+yUFXzhGuHXD5Zza+b21sRCA5QPPv3
B5OM61GrcyxH2+muIvAKK49NJGNeN+YALcSRuJv5QCko/8P7/FTOaswYDWM+2rceb+FCr2yWTDM8
Tb7OSqB13rn7BOawgMz9wtdU+NVnlcxIue9RpzsOO0UTD/E/lCjki4oV84xtBkH6qoh7Z4g6McQg
NtpCtfIFntNALVL7o8Fe63+jFgYCrjjYO+Z9hvv69MDriqgcusqAMQ4gc4TCwkGVYtoB4RUbqSV3
X3MYSJDQ4SXLcAktMWEvpEY+cR9Cy3ba7bObMc9qkBUMUZXR0p5o6inTOjUaTnqRAjJfjg01D4/5
9GfEBxeWeG2E144ORw+2zJBk+7WzQ3eNpJ38j3W1gPXd2HK60RiFagVDu1dACj9R+cTgsscqoepN
NDAkLL8t1npT9kPdMqLONrK8t105WT8MM798t00mNekofVAo49qDj1yWWIWpNmdpNfS3yA23wcl5
yJ26s39KuKX4LnKO6Y3pn9hRYfz7O6b537WDsZZ53bXQJGGi1LOdeb+IOhN433zSc9t1r0oZ1YJG
whgFMS7c+/OiIKE0u/C/wy4hEbb1vkfJzfHCoP36dZ6C1zPiYkP6UUITKcPXRd5L2HePpjWOuW7I
0WQg4XNjfrx3EHFQ4vmsA3BdFXyFOJAci6wYjkHk6xGzNE+nacXqFize8c913K9RNDlhqIzbbXnB
+rDphEmOs4I7v9zs30Dp+ljQfkokWukZpfXPZGSwjptohuU2U9mBHmeD9+WUqRs22Uv3zZjPE2ba
ksL1sGSAxFjsnsbXAB13bGe6ocX52i/rdgKBYuOY+ONG87XB/6WP0lalT/ft5amgHeX0NMqm3aAt
zGwrdz4/fDYaNjhTPsKAxnXcbGkWb/BKZbO2ETfQPH3xVg1xSOaf0RfUpAKf+yMzwKFi3jhuJNN2
eTi1smhOfvZKqUyfNhNvIYIkEqMO3/5QiXQ0NVuc1cope0sb4ZmLONyRm593Eqyii+iYNp9MzZmB
8cpwkCpvUPanRUbfS5Fq79dLAEgQkTeRBxWfI+eFqug67951WeIxiprBLlqgsS/fcciswXPmy6X/
7oYUIfnlBiq76JixCk03++H3SFfSgE9vyYn6QMdm6Cr9OkBQN6CXWV1QQdliXcpjrmQwrf+1kgse
BxLiFE2a/Cv4ZfR9J6crDbSX5stvcbpDN9lkw0Ubjq16sAWgNGZ42yfVH1a0lS+0cF4QF94gGXwb
iQi6KSCaLDI5uAjNfCNUS2BJSR4EWZ4ZPIxEmPMfG9mxhN3CuFaXSLl/VtzxKJ1Q8qcUuGvlVu+R
JWuKKSd2By2/cdJ3DehrqqZlpGZvSzMtJI31LduNomIdqZGIdTj/vpPxd6zpg/LdYKNYGTXl2ItR
u6hrbqTIFKhrvvccWy8umWpneqwBv108v4MKdZIBDqQMU2VmxwHCYiF2uvfpcuUOlT0ZzvdI/yaS
4U94tCBNYq4A8kN1ot1N69Lh1HkJc+LgwLK6QIH2aP5KIk3/hOJ8wAnSiLTD6/r0eG/Y433/rQJI
YjjPj8yNEQbzz2zaWlFPLGtwN+8zYJ5pOkwZanLoZRfN+D7Vi4Q7Z+f3/H6Mypm2+sqycL1lAxmJ
O5XsQU5LN5mq6AbNbRz9Imf0HO43SX9txs2KOXAT6nf+u9Yn1KFJGwgdmCdfK7wOsEo7Ul8FhPiv
EH2lS7QaXai+PL0Ru22epUqohDqtXgfdlNk7ERSlyXs1tSZbub/+zNWkWCIxQxZ+LCmt8oNsYe2A
6/hzjqpvcFEZgdyAvHveTZa0gpZ2bSkziOqVQaAVqbLnoeo2cQFz58d5NJJJt0d67LFvEE4D6dgI
TEjmGxYY/BeCnEDh1f4AKjKTAqIAm575eNYZ/mbbOjLcfZWT58fLFxSU9BWyO4Jab44ww7j96Ky2
OCb7wSg7x/bVGpEo7+vQVIqEod4CuZN1bFdg4AQLDN6VSHZB5DPQaMBgNTWbj8R//cPjSIF89PkU
DDkFgW/173CZdCzBRRxRXAT7eeXW259oKjeAJj6Q6qOYdVoUQG/9AM31VwGYukxmOB6bwpuVCWGn
tTruoKhYSz82GXPIsBdjU0EbMX1dMVydPPPK8+Btme8cAcxHLpvV8V/747iYpcgIdZVF/ExPaEgk
tZYwIOjFmAxgUnDEaaV8ahohEmObYfL+g3uZoztZfi9U4LhdfzmEpDlEU7BX/9dRyOGHBDrNwi6u
58I7C4pw0QJFGRfm6qPStsaTaiyR9o+m+cGvPBu5/mJgdlD23gGtSx+8fehFcBvQuguXPKqki+7H
iMVSy0RSiVAiHQgoHywrhnYBYv85/43XuMYkRpe4AqTJRzn4LLGUooP7XmSeniklF90QJXXXgb9/
LOtSS6SmMn/xQnLSH3mKfkbK0fRDxLQGCdSlh0DlMF3sh59D6zmsqbNAnR2MWd+3nylL9kz18N1H
peUnOb4rJSaYVUXC9Y+Mf0NV0JopwhyIznhCoIsBK5IXQeDelAB8K9bxtSpLi+tOSK30W6aNUDbW
83OOdF59XzQ6CKnCqkg0m6eEcqT3FFZqYHq0iYIip3iEc72YTya01obRv1RfipWmq8UvkRjZO4lL
GWaQP7da4tktGRtrASLeVcrK2jJiMqKd2O6rKAVbSMjVuHvvuBWeJUeGoD4CelgJubGn8SRpmYMZ
/8HHOQbBupegMVJ/MtnrhLP3XVIlGAmJDPIvw/YlGRKJugyW5tnUF7GPAJzhjiCsXe3TxviHTDoO
4IhqIgeAo0m32pGylHtzAj2RKc78uHyo/pZ6GwYJ9aso2Ri44CUjumzjmqyNNbqG0GrHP8zPaLTo
WW7gvZfvx9eTfMFgE9usgqiTssPqX/XXrsJWbwJdeT7oT3Awni4icrG6XWp/imr63HnLWk5pN+Ae
unBJD8MjHOUOJOVP/6DZZ2dxILQmHjD4E1gkevCvt4od4fWfBWhGtZoVjJQZNxfoUOWq5HgXSs1I
sJLPzEWOvcMVLFOp7dn8E3rRjWxSpibllKe51VeN8jKSwytN3egbkS7gjv0pXlc00lIARD2Y/TRf
qFyKzpDwdYJIMao8aFHHGGZKyIDRv6q4bgVgUVqqq1n7SW/V6DR0PYQYJw9qJiTGGc46IshFV7s3
KncmbvhXraqtNdNOPAOTek2wgRyBJ70qnBcfULaXGqRL25+ADsk2XEIpjqZ3zb9j5m+ye/oasJlK
WfocnXJFS2Tow2DAL5QYV/Nb1Ncfqa1EMjOOznogpiIav7cr/gNNu87j/0xxki1Rqn1DvzF6WEsp
rI9GRlgR/uGl+o3p4FYKrQTcL0PeGeM+WnNkbXX4AqPxRiYYydeo2N/SF0h7Z/HJ9SRg0EPCMy/o
Xw2XfiYaQPCaL4QPc0qLaWeAA7lbsmWxQh4qYJ/XrQCDXlT4TAFqRKIolyF8/nWMtrht2mtyi/Db
5qscm9rtnJsFpO0NHp5BFnwUlzNxlaQDTwC/JE+oZa6ygHvFiF9ClMhgV6eEewwQJpcaxy0BJT3C
QLDzOPgIl9w4ckV6wfCRLqrEEyRrlWnXCtL2VRDtdcivkVGHoEdxg+86RYzdOh2I/wYKsJz/1ITb
BD/f9iOBHdQo5voDm3jfKbWB85rdKwSyyNGE9aETgjZa4+rEBEJj8Q90YQ+rD/2z44KRLNoq2S8U
MbIe0t2Qizmt1tuLWTcQ5NC3g2hRWM0NKHazHDuisWzTZQ+yNVvG+HSoeDlJQX7xLmHB+VTwSxj3
PcG5Vd1/xyRlFiL/qju/sUkyta+nC2JxfjBVn139cu0WZHRUTnc6c3HYFQNzFzuX25ocK/6JqYBH
MO99bdFQ/J+Xegn4EnZIrU2qQdJpZUPEdapEt3GPvkdc8KHsEC9WGIsUmzMgmD73upxNbgutGnXQ
78663/QgrGb2ayWmTJU6HDWAzyJzQv+LPFqOFMMeVfKQhUvioFxQ6muIdQV13/LBpC5izQB9GmTe
xONA2ZqgzoMmfxXFUBcffrqRwyz7YKwqw1JzPx0V3bCyfhf4+c50cPg6vCbWylyqgvffMDmYeX08
MXcyOBY1gNfe0bsSXP8sTjLHjNhxQeRpHbM8WU11Bx0mqgXEBXikFvoykqHpqig8tLA+gwRZlbWM
HxR7jm8RpR4vgUAll3cSpiF+8dCG6fa/d93cOS7UWSqq2RsRu+wSoSwfflxhscocgXieWFarlzrL
7KQGtLId492CSu4OM49EmgJcOyUwvaFACs8t8vighsmpWV8y31MxGHVV51LYXNSDgCWljeHlsxLh
Ms0pshUHxblY98t8nMacFJw/kFYq4+TJDD4bgbPM5wxJ6Ob7X3MDxnqSPIwrGbP1U2NcaBqvm1wv
dFZ+BG/sDYVADYfLOLYWOcSs32X8aR1lcY14rJRs0sp4OEKXiHM1HG81ca1d1JAGmQA4oHR161EK
oLaQBDsx7O3c1fbhexYg1OKHu4O5hOz2eOoUY/8g8TrEbLuWv59nf6Ry4Y9ZR0qXKrLaor644iE1
PN44Yn+DKGO2NC98I8TBBD4FiONPRNVm1v8TkqrtXvyqJirbw+1GWj2hetnCSHyNjJ2fPWlvh2mE
bjokFz7hFnhUp91gKNm01XO3QHnxtauX3jwourNPrlQ8xf/sXujKK18poOdcRiQxDPEt30MQRNqW
XuIRNHtivwaA0aVRCT2t4Zxolc7Ag+iJhkBnoLKXRvXIr/q5Ml0JR9kFcRskJgReHm4Ex/eQcLCk
PrqSsYqzHi0k4HPnLthWof77FDG/6kX6NYB1/tm4vR8TQ/2l8xTc/nbPjzVJx88i6e5prbVLKySD
WA/jrC8DJQTNyXWQj3AiLpIewVaFZSyoZPjPiQfNKl54ve6ts6lSHZi6J03Wr/elKfkoK9czaxXD
6yk+IGmc85nPURJj/twyF8w+aS+0mZK+Sd6eTExgAOUSVM0+PRSv2BOIMHSDjwa+OF6ySpnxUbd2
EAlnJ3x9c3THQdcsC2DIvahbn6GOrLjSekrVipZk/Tys3jiEx/abjHnt1rLdZyexYI1hqtHcadD7
XkRZEzAgLp/Ecm6/u1vxFmzsJTfLDcrmdmTnIT3kOWJLSjYWKgc+2yvEcR4l9GhDb6zBEsmPb24i
sucXMyLqGN4LPmoTzOCExWZTulowo0NlTdFV4u+aECOgVvQm9OLayue2jKNQA5tyeER5f/w/fK07
iORmpURPQr14VaZc9VGIuHkrO4F9hPN0Wl5KIBue6374c7pMRUcCaRHsROekNc4+toKq6a0nRvPd
E7uhu8cHgFdeLAX5xqmfPWz6oRxb1UKMnzmmDFp3M92gqGOOYmEHNYxCny6a8JsdoH0JeuoXJ2f7
GN8mIuYEe9ZqDsaog6mPNNtIL74jDm3APwLSEm80FqF9QYe12RBXc+C1B1cLZomDNo6vYF9SWgXv
5rQnn7noW1WUZbo157H509XRuQ9YrYc2qCzlRzniRR00ld7LlXsK7XvZ3loCrq+bcQbNN8X9iy5v
Z4g3wbFGRTQ/JeFjMaQfCxjiks30g5KCzVAk1YvM6Itu6eqVywFJZkiwYDK6XrPJuA+n/u2R/jvK
2/JGed9oIxE/3hOj0RSkwA5Lp3zm/hdiNx8cKucwQVS6gBJUtkPB+dz4szia7iduLTArz0d4LgoQ
AyJ5b1XvCoPS6IgfCpyJKcsf+j+qSAp9eRP09YeAF5Xu5/VAzrMPbNCP+2+OiwQYVTFBlBmIyZ8L
NHCukeX9hnBC4ff0PtxkE1NlBHmfDhR4ev+W5GgdoQZXRB9NYQQvSR/PS+D8ury/yHZPA6YH46Jd
rguulOLDu9rKDL81pCgUdpvIFYUvWBEpezYnMb0msv7DnL1jfvLQV3aZtHeLxbl0kIKzZeVQI5yj
c8vj+GXrV+cMf3/v4hQ+bu40tUuJM4R5LMjoSM+8UehWR0xaJovfdbk0pvzI7OZJlt8uL3+Ou2W7
t1PjSXGK/L9dQzOiOJW0MIjs0+B0XtowBK1f7YBOG130BKisbc7TB94F/iH8hhzz8TYi+KTzFAWj
TFDx7q/kl1MG1MOQw4aGa/6Exrdu7Wxjlb7NilQBXAlrYKqfpDOJ2trTHo+ibx1JQpdnxYGMiH2D
LOjj/MC9FnaHmosCnzknvhpdH8SPYSxrTZl53mAaFOa0mIuCI3FSQbxrUwnv6K8/HREp+a0C77/g
qxkxf3+boZrNxnPj9GgbbY9MWeaOLXq1j5ptOcn1tGuZq9K2ldYym0LK2ePNLwxv6Cu8339cWTpG
vtRcmYkTnZUqLeUY+RyzLTmQvsOP+OTRbOqDFSVFy3CwYmYTgDeQk5gkHGEeKkgXSt4rrGO5BSic
l6Y8Flc78LxxvXZ3v/MOt1FVoQ5rcGnaXAHZpATJknx5dS+gunIs3DNUpI8NHyjszHrREqy9uTDG
l5CX35AYWfwpYbzvxEj8auPCzpFsz02Myupp9XHOgX4jzGToQ1Bxa2iOHWkzYsVb4MmxUbvq2M94
y9XbCnJDYFheYtrzBnxC1wlQcCQYwZkjK9pXe23yB3djK69Hh6KrBwT+9kmD7yXqvxRziP9fxlFl
xc4vrBh0/Lyv1egbcW2+p84GdRq+SUXEkqRw8O0fbE34Qfy3bM/rdGxeczmLeepmcYOa6cQf7UR8
mhrZ76JOKYzXTw/rDWwng2xm/4Pn5vY+6XQnR4xZMl3PEYynvl/kf1A82IRyA3Zaoc9RBYPFqhf7
Tzh7l9orISNV37jgFn33u3sMs9xOCQQu5C5ybavNZJzxEvmpUQphGGI8UP0VqT/Zf2sueAX0d9Zo
TKXVRTNXWGUpdq1/sMxCKAyOUIRWQPpvV8Qq5vBk4qAbshX54gLo77uq2VoP98RafBS/77UUQgvb
369uG3cwrneV9uVNx83w8smDnz8Po4Vh/NA2lz24e64AaDRDwfTWTktTJPJFha1e/eF3ebYPM2OA
26ht36d3y9Oh8ef1cWAvhKpy0eirF5IRZ86HrH6MApPGqcjlbR2qJ9vW4aSgCV2dYJP1nsjcCYDh
OcX1mQe+HzQCbwKIjE3l3w5KoDdISLbNzpdR7KH8wvbFRKPZTPhwLeU52MNT+g85U1pV+O2jz9sd
T+IbcwUDEWp1We+fbb+GzSS5RtyK8/Bc/uGUaNGS7xxZho2VIGsFa56n1BxAvlUQnVh9t9pv/560
IhIPX+i2jVRQEYFCifYbrwIp1XvEo+YGm5DTRp3eW5J70AkKN2duXnJS2dWN3BcH4vVatU4vD6kM
IiA2ZfMj7YlEoxqLVBC3qiyXMC+mnEHndGZIL+GImDmCF6PlKjInKKGSgPWn1e+jjGWhjWES2gT6
lXt83OpMboiYRlEdqRoMEbt8P5cYzsAZarUKsQ5WHi9cVyZos+9IhODKUYc7u0L/XA3/6yP5+pO7
EUKpaYhEj0+pyR2oHgPV9196luEz5mbiaPckpT/2h6AQ2b1zTwqe9h5v3MKdcti7MMng+gmgpNMz
X/Ye7W7EXLzWcigS3aV7shwdbwFxU9fg/gj86EtIcTc0nKkAj4lED8IZZvVi4w3+lLBPnQHAADWA
OWA4WOd+5OVFkUMB4brrage9kYTa29cAJYQAtUMlLtDAodf+Z+kQglfNN6GrwTJ7GBZB/vQsQ0jG
l5qzHtfHCSzEd7a4qpl1oUPX51YJhHkMQHa4zKtfr8X2gi8YLH4A/OT0dadL2lfuYx+ivqOMbP+O
i4CxcOB8SEvG77POjJdRVuAtWayBf3Is4nsfr2jpSK76QzVv3cmZaqbQSjBjP2KfJ9gShj6fKus6
DvJVssfMqPu41AroXMEDG8v87pVuw1yEiriMlVVMFupQ213bqpHmKvUjW9ueLNzS2T2KTla1pAvC
o7Q4YHcuIAJUoq7WAcpacnYwIE+FPa+70j5ndxHs54yA1VOYG+fyDp4KA3kRimpupKOb8XforjXS
w4kXpwyfbzccVRKJUdfgXqMkAFoCVoWTXaIW9tw0Wl5L7iNICD7LT5jxzf1TRONMprM+LVSmXxUM
xNxaHIRMf6ZPE4P09ZQy1SHOw1jPD3IFdBTJQyw2KuTZWUFnC1fegxSJcrcTGal/iD42J9HZk6T3
57Ml3owx3+TyxxqfbbPGBp2MNBqzeH/26n5EXHX27cTCbJ7y1V+4cXcZ3CYLBC8HL7IbXOHoKEEm
TC8rNhbgDnZipkXwmi+EyATRTyiDg0DddobjHH5ZK2hmGhNQWjgn1tCNbKnz1rFdO5o6G/a3Ow6d
CJ4DXNpVnxqaA8kIpJkvzWjolhRwRiizSY3gUBoilU92HXgXsRrCZWTjDfnnZIt+dpjyF+UpVHBL
puxIKxjGjKs/8pYJUCRG4XUHiQvXPEmDV95fRcbNuiRBIqFG6U7TZIFz5fcGUKWotIqaD5sMzNiG
iiiliE8T1xpXTdNLYgJsFDpZL0to+1deQ1RvCFEV3Afzga4Q6AC43pvP5nGwaDi6oR7ZJ/OKE2pL
VRkvnEorqNq0psEqsArQNW/OPeMHtIanT3AT+xsM/HRQ2jYfsnRXagw7UUpNhVXHwJf6CIjBgCrD
W5KbIHT8C3rsH7rtauUJixEQ4Lsvv8/cirUDA4qx1AG4g9XWkn9cFeG4yf1AKgYYENQambwN4KGh
JtdiG2PGEQYNRJ9JFjvcKJmVe5ieldvkScnhAyzbgyvAs/nNuVQiKuv9dzEETV9hSnXzC0InWsyj
MsObTx952V+NBgP1wv2Q/UX4pn+epVrRm/7RJrHMrwE+z1c88wmowuWf87DWKacFdyFxfdzvv/RD
p+PgBdHKE1YPaJ5T3xRA3Ro0VAEHvhYFoeWbykNo7ME46ACEI4nJ9H1P546PIYUyNYxTP8RzLSyr
MecRTCdJz7UbJLGuoKS6RQio7BbL7/AdjtV8eHUKA26uOVDf7K3t8bDrkGoWRpJqGv+Qe4QVzLSJ
agNtLE4/J/Lf/1UhmlB1/osi+DEH9g43TY9HvZ4SzUoVh1ps6h9RXPyuxf4ijz6mFfpsHVe6tPM8
FxMOhdzVqdBf95BRLBm7tJRe31XZKIlKj9ydalZahzvAoceJPV4m5SzKIWLmzT4AuVP8p0zL4X4y
sWzgW6oAUIJRNgG18r7ndbc0oaehXPYeeu2k0kjuhmjCOAfonz7NwMYXtVr4cAvkKqZAz2qdbyn/
MLSkJHAKM8LmRQQ5cdy2Jyru5Gg1kg97SjAQTZGNJomZ8WudunJ1s+48DVjT2sUK1HDImTn4OkSJ
rLO8p79Ew5tjPSBESq7jHC3Tk4aUxewmqe+hWTDU82jLkmD/BPVEJKVFvDj7QHBqbAH4WzGDuRN6
UUr/dwRtG1VwIDlrKxO+aaKToreMwg9F7RQdSphVxurDDNnloRab9zbelLMJYMiid+/77wxZnzj9
0p5TbnqhG7weZNNxso4pCxz5B/IJtkAzm5cDwrCOR0ArUdRqKOCcS9TmSajK85WJ9+PRlw3GXkj3
KOzr2aE6JRLjv7q17S6kzwkB5oE1h0weRPBB7wq5sK3ILWtLQv06w5nvGILddlURclqyMXhtiKzA
HFyU01Nf219C+gWtA19bCLmGbjFWHDfvRZvhgXhDSSbnkFBiiRsADZXNnczYt9XPb+urSXII/xA+
hH651hl+G7EFZ6w5dyLlVXzDrLAeJMwOdjMzoA4awWJaX2ZHRZzattv+sKhL2ZGGuGKiThc/6Ccl
o9UOHY6gz2337haM+O90LTnKaVJ+EGjEIGbTrTeOp4KU6u3hCiEtaBOslr6huBEhZK7+YWMREMgs
DlAeyZaGDmd70t1dYL2CoiaDNjYmnOXpeHd/GaeaV2E13D/eNbXYPqwrUWScrzUDuZIO6mWZ47hr
1ZKWp6Qqjl4piz3tElw0Gh8pjIJOFmWewj71xPBc4hF69wmaVBN9z+hoYQm9sGqewDg9AzHhtnY3
7EgwcuCeIIfOQQneI1VcaPd9rCfXJUf82iMA652ZjY5X4qiHYuaqifNCpemwWffugK5ZFB1qjjpY
JXp7OXrxGi4/x1yY6kLXcJW0PphoAg6wi9pOEkRMxzbMdn4RzUdbgIVaKayQMN4zDXbMXejpQfUX
XxfBZktGhBxZS5jFuBH5Fr+FHsMrxKvTSvVK1UjRpdgKizG/JGMlps1g5n2BoQSGhZ/+1IPyX7nv
KK1Lh18DmacINDjVDOVqHo6EQIKY/fmzXnJfTV1Z4FAt3pFXtAn+bDJ7tyzTOBnR9upEaLMWr48C
/cdOe0hB7DqzamNE/af5pvQdJG4lvrH6xoggNBai3f0bO82dFOYJxIARC5Wc7lkyPOJWeVMXHbET
pLWH8GV4VcnZ1ZXlV6S6u4opyI7ZK2PicOk0t7u2sGlEkb0Gny3EyaSgT05Lu0GKiIOK4eLgar3w
p5De2tAuWOIXe8iFZkc0NkahlVzwBIXPrCiI/XdlEWSnOwF67QhXkjBGwFLH685hh55K3sH/C7u2
pFRSeciINdA2iQVGSN8BbqFdKM1/9vp6ExbEYpckfTdGL9mZvhZ3oblvz9kvxhDNy/5rEEc8SZhC
vTm6cWoVXxerZF/uoRUa/HauhFRLSajVXmVI8cSb6seFaQcc/BCZE3FGEfK8c4iZAVhNNzR3B/ap
CyvbwtdUp8uLX5kaRGEVqJIt14V6j3B3B3e0tmfBMj8T9qPoRtZCSykS8ix9pVkbG5KFnkOMouww
fn0nxLvByFwlc8rU2jDjWCquGTHNgMEyuVP1yXYhuhDDhlGz/ThBCJCjRWwlCjjD1M0xz/n7rz7u
5NyYCy1Pwe/a+Mf10cGeh8KjRZ30SpzeVyJtiSbIs+31UjovZyMNlID2zJ+aRsbuNQhNuDezCv0t
8oROrGdgkGhX7nVvnlUwlMLbf77hZ4nOiIBcrGZ2KSEEwfnFIwpCjqGG5g3SeVUyeA1Sj39bVSVq
Vp27NrmGFIpKDhR8OM2OnUC+26FXgvki1UYMtqXInOOqZoSEnPRdZ2tk0GzG4m7y4TtH28HIKsGy
9TU1hhEKlod37A1CKzhMWpv30AurVR6fcZ+cp3Yd1o95FJ9wx16nQwz/90xFHa2f4sDAlfFirxqk
RWMgOD/PAkhrkNinnJFl+Oefbnvo8KxsyuFZqKtM1TANu/GHPX/aMrLYaYKJgxacISjFP/C2IM9T
MtW3BTT8nB5dytx0NlzcyZQEXxZtpwG2cKAitzgxSukgSK6y4/DEObInlQ1vnYsagXmxVstz6pqI
7wXWJC1f6ObTY/e/laMaf2UIKEqztI7qlb/vkPrlrdkKfd+sz3NX674rEVxdz9MhzZwhGxSnbdrN
Xd5HhQPsPSE6D2wTXm7tqjs5bNXdrw8TfZrsrHWlKMYUa/jiRrln8IfpQtb42Orjx7EZ+trY83B9
qCi8CulVZaWW/CxpOgJmVH8Q85sMNE6oIxrEJCVcEko6SMNTiRN4NdwojNI5A8NjRrjfndZJ4nSC
8AKu/s3xAUFuNbvS9UIQ+xt38WRpmk9n92k2jAvnWTLBHCg0DtZbK2ScB4CwO35FTHvobijRzZsT
OtlseG9CV5bAVN4NQQ4f2gWufPP/QwGErBqONFxvFYn6gjvCvtftcThwcNDO5NSNk/5QA4COtPFr
vq1BiiiEHdunoGd8hDSDtp4AdbIAmkTcxLRpMShYrG+ytZdiNqCg0MtF7dhx/0AZJQPU8P/QmjPA
PJHRzt2LeWDydG0ju/oDVpPwBOR7iHTXAvbJy9ScNXH7ZNaDKeKFGXg5JBOVSXeyYbNWo0DzMQsw
Z0puOjUW5zcQ5/jyNn+eQ9fINRoE0jliDgjK2jO4hO8JDUq/X9CO8CmiWhctyz02mFKIdg3f6tyB
wRMZoGGaRFUDGuUDzjXanOfuZKTNtRmDNNtcm3YlvdhwpLoSVY45HRcT1Wmh75tK6lro0cJV0Qa+
5ayHIfyyOxpsKwRrrEr69wm2nBrM7lBpme4g4v+k9isR2IbRsI3qlIJ9cQ1a9TTrxXJHLdyMH4jH
9H/M6H2CZMujkyVOSEHJKOumMwcvZpVz3pLfDHiKtYoEs7lmp8HI66WchOOHAOoAKpOgWXfJ/qHp
6c74dtbhD8IYhYRCEKPJCgN44OYr49A/VaodoUyHm+qbqASeKCnelk/wPkJYlOXe7vxovaewIxOs
Mv/ac74g+ED6s/FJ6o6rWGyhDWIvhuAasy+lHOF/ZsRfFe8TtWi18qVWzifBaCy054aOBUhQ1p9w
C2pqZ2RZqaA7xgFr2VeVSlMug1sDWX+tLcWaowt98yorY16FiULr581yRcFJuEX2Fe5vzAA1EPVm
+qbTNT8gwWyfYKUOqCHmtf8V/Laxt4pE6f/fibQR6/t+cbzpj8zLlCCbnog6Hq1kMU2jF/vpPG8H
PehyDAdsJY9insorNiYXd5cLHPZszphc3ITJIOYx9QN2cjVJiXPGwPfB2pyQ6E7Ul9lRVfe97opU
f8NpmZDzzT6KIsoG9qAM7DHxUcVrEnhtWapGzaYJ7ZkzqRNCMKNrZBHCyfr3Q1F0OVsfmSXOxqXN
LbS6jxhweD9plQY4jc6s9nAiR/jWFsBaGS0/ExBR9ji7sFIG2Rfs/koV7HTLMLSkAW0imhHpYBtZ
fqdK5GAUYQ7CsabaZ/+NHg3y7F2wLbHX4UPCxgL7H9pidQehiN0g2wgk1SrYxefhJZg/39A5vJpP
kSd05quCnYnZmR63aAkb3mf3NEqfAo1ouSKpB/DmvqSEalMRlJhZAfEcSDnT2vQPLYlp1mCg3rDW
4BuJJF2H6csteHS9TeDKzhCH1ovLBxvOrlp2tGcxUeHfd41kLqC0hBVjdwOOzcdnqukBiOX4V0lR
lNJO7BJ2TLpicdLhL1kTTAg/41WQNYwd6WuNTvMNOr+e2F4Fv+NsIxuPmK4142koLrBiqt1zPLUA
sFz71JDd1fCJe8iFWOl8PDNmhX4BWcqP3WQ4UuG8ujMbajf3SnIp+5QDT+N3Iwh+YlLmAPkw/YtW
QRL8M1BeIzkiU/IIEgcHFk6+M2LsXPiAobUzA5b6N0LERlQHkkXxOO66UpFciSOIim7/HeWbdg1T
Z4Beqcvz2+bWW70X5bufvAgtzQX16M90ge43wfFbRjKVJIwaT+/7++5QCjPeb31H2IaE4e9ucIZ5
Dsr6pcRDr1vVgSo2h6/snU6Pb0rIZ/jZGqLwI+AZhVj01eS4Bli69mcJNxgli/Xago4lMiXn0msT
peC7Q2RaGxp2oklRjHF/d/cUpY3JG9v3wmkUKxUvufCaBhJlDHT3+/WSPEDSnKRoV+ecvicHAqvA
O9CoWIes91cS903iqafygNMn1Na50mv+y6fBxxruDd8dbYR2QA8d7r8vOmxBwTRxmkfVQZ2qKLk5
0b4qgtUlm+GGbSCaIvLMTRjxYP/iAo0SGWD6tZI19AaDExxS+7rQcK2UaUyTbkTMHztKhq4J3eqV
Hd6/9VmX24HU2iuobZ4kZBC8gTf5ffqi2X+D71PzuLwU2LUQjxAq90JV5nI3j3BHoZzgLEH9X7HS
laE3N7wWAXvNGlzjSX2AsswyeiQSkcrIrdXPdapABS4Z/WsMzoHv9KWrM75JTxRlzRjcaEAkbFeB
lgR/0ENx4xHzE6DjB7pKTd1RMvpiMaVpX+9YLjjFhuaLxybAohGAU8BnvTb4mznJjq29o2RmUdDl
HaY1ExafURV5Dc6kg38JdCG8xwBv/RdeIlKfoLHlZeT61BW9jJms4pb+5NlNsdJcyy0pQUP+iSAh
9rlvQdqVPqiA+ZwVZZYqQIUH66D+kEqz+dGCA2cN/wvudIhNjAQWegztnMKKpgMXpx0+219Dz2Ma
tNg6t+XWMKN6Lr6GuudGpJZfA/T45InWnmSVCIAksC0mKEzG33OH6LOkvluuvOSOym9oDl2J0UNg
IRuFBibtQ9QMdoMbdnoc5jIMRb/YfogM1eI1V9lLsdJGPcqoZzxWZxvlCM7lYTMWB8GQdwt4zeNE
pSRrnHunfuL0jPnOw3czFrJQ4jged9UIgfs103Ny3+gYGUJuipGjlhg6q9+rdWgF7Pt2/6K6/G2m
MwLo+4mZU+qM7xplHZiLMsp0rrf1ufj7nPIXbUBuBJsDw4TY84jovyohpCFA1T4hEa97WUXSB92H
vwqxGDKV/9Ezvdcl8lVZH9iR6QS8gfUFclwGlHBW12xFOJnm2+I9KYsCo3j2JfG7yiYeunAuQ6o9
eOZ2XmmKhjDmMAzB+RApfImUjnxmrbB687loNNbm3FmzvsJCxRSka3Xq2mVAztPsXlKXjlfz2Snq
kRA7h1uGEDWAr/NwxS0JNhgmEy7lmN9fAwqQ8tlQTLseze162DcdX0ESY+QChMfYQXZa2vMcH9hv
cwhgIyAS3tw9IWP7CgZtwUgNubCF265YOjpyQ5PzvXnxHGpnZ0Dwht8AcYh+58lZP4lDDIpPPbVK
qu2iyJobBCHoAYrcs00tY63/dDJalFL8EdWKu2FQp5OpaWofTnUDdK7zZTvbkrdqfe+aWPzuDljR
n2T5y/bANEmdBQfxp1rxO7Reo7Mz2El77V2xDa392R0Zn+VS4cfq6XnZPh1dEpoELiSBrBr9eP54
by7nPvw5sBdTuzd3e+L0O172P7HxqehAMk+vKISjzgEnI4Wq6EC8bdUYFF69v+LOeYDV5iCbzKsM
DulmfSl9UyX1gXtMZ4M5cpLWgbjiIao4buaACukpSc9CvfKxPFnszcWpZkJfjuHcQ7mIeOqQ+tFT
Blq1caVTLoAgr0K8d5fiqqMc4P/dJG8VqmGimpRGlrLsLWaI1vBiFSBp7/QMqtNebeAd10qowvpK
GqWuf7hvznN3OBAOFlC2hnnQ7gZa8hqziKAknUelLNtla59JFE/Ta2kooasaf6FJaljjFQ/eORQo
8cFRQVN+avKpJZn+jEjzQlgkZUKQznGQgfmlVlTUd5pvLuzf8yN/aGBDmEpVB2X8ZvOKYfkk1VEv
ocmCJNjBSC9ZMijZgN2LrBW3oDwleSKmcXanF6O6LLbbWxU+SdkKNFUDDBAhZUzS54aNrvX8qXVl
qXnRFgLx85YSO1rmQ37gU7KPzgbHQF8XmgdtpRqh6TD6PgBLJgT5taUpknzct47fdGl/eaP58l3J
AJeiCRwsgWCO6YWfPk3druEIEbIghSR1HADyln1iPRibAftH86Ihte5XVL47cSB3++0orrCKcQKg
aEnx4HZWaudUy7K2lxzaFoCqWSWOo6lBV+kEkRxgFRZXYyuD3K2arKs6KMgM/TF6TYRU5iiMBgJH
/P/4oJkXQJ/yToDKkDTFrB2OxmVAnT4Gq/fGOMSwZCxwfvrwvQvvCUrL/IfR+qu4TZwwJhp3aq4/
fTNZFQ3wwRuJ5bXP4Qa7nx9IiLyy6vlWfXtNk8azQutG4QSjxN4DejrX/9YxTwiBF15fiNdEeRvX
eGjNQSSg6+TquMp/BiZf7tn8g2JXh3+A7fVRdkXNBhRvyjSblkgbpRgrRCBfDNr8rSUOpMuzCl45
wiXKvGMFt7ruFlqs3T3vYUWfnJTroOZpW048mtdrXQK0zrTh+RfwoR+TuHdUaG5aDISOi8h+6Kzi
vEMcCuAbL+6YW6GFfElkqRjmSMW0fvjjvs3hySd0EZudhv0IiT6zp9PMXARlApxFg2OajL59i+Bn
wy5JLGq1bLNDu+oW4HaXxxXiTnhLS/PHGFPq5DY8Www9FLgvN4Iji+ht3eIJjUB89gK4rreZ1TXT
jo/jUUScJ8sd9U05ndR5FO+CChgTT37Kbt6Hh1wKxol9v6q7nfcov12eX7gS9viaN4cpwR84RBC4
WoFNEQbLS8p/cxJOeWyDscLcPjEZLuqSV6bSJ/cDDN7kTVH2CmzkJQFIlMNIfgXC6zgQcttBEm6F
9VJvXmMnZEXhHRawE9zIrvPdn79VG59zr/yNaxONVTXjC3iCdlapWG/8/SFcSHxlPQDJYqvG6469
QDWVXYGzUJ+h5uz1msAdgbnYG4wCDzXRP71OtXelAo6pnRDiRBt/wHV5nvSRc5AqqS+2p4baS6JM
kIyghLAZhMuQd/XIyJqnEap0fZ74MYdbOdywcyLEDy+40W/b/eJiMHiVE7SHmzBYi1++eGTVNwqz
dXT1EnjK9846Yn0R3T11HLNstARKo47pq5cJpzKCnWoglhnd7BgeYo/9AAz8ChlWXMf/z80YFtgh
h/9NsS6gbd2Kjw6CyafisHURJCVknre0fRAWiEECOApFg/3R4xJaJXwQ+g51NMYys/4NIoMhIXw/
+o8EkI7BA3u1b+Su8c5QzhQNhz5Tuc2DBmiZBkN8QIlB28bLDQgVtXvcuWREr7Y9UvLPcwFttiov
37Vj7MTnGsMbnHG6IYpd/i5HXUx9r72vcu0agD1KvebopKCu34FHGW01ZOKVWOwPf5hIIglJipFu
Sx8ZRh6wClr3Oux6M/ZP6BT4gFQJqr2qubOglMmAiN5K4qP3vEm1t6LhIBKbKIRhBB7b+mlV9NoN
Bj/3ktA7N5zYkFNSyj+sHOZM2mVppQYaXAiRBOr4Gdqxg6Rx1imXkYu+RHaKLYMefS3Gf4fhRNUe
bYK41CioLcRMlH8N2cuQf113VGM7OGqtN6rNR2+p3sraMFf0P2r6CaD9Qf2LGEV/B396dny4ykdX
KOlb3AoPMacbRU6/8TBMFyrsTHX8O9P4Uy6FMtckgM8HLBU7SyR4GrgXIo8JJLcEMMHMnXcx6cZb
cCRzIK0zjadLw+OuPe9IQ1iHHrkAWZmyZCYdbndy7WrgTlMNgEl/0rWM08ps5O5vFQBJEr1GWG1N
oVYqdPVyh594Ab93hUFPNkqBtkf+UTB6a+/uNGwuPJJa+tlJvnNDQ5DWABjBGGFSTrtEHehhGxAs
SeVlKLMckcBuriJ8L3wyi06OeH+rml92/INK8a7rh+LWTKus362Gmf28Qx1suso9pMUGeKKgJrSK
BV3622N2Xwb6mpTloQYKBnwFHmdkou0eJuwqEmBhAZWt8+HH78goGwAj4ovDfUyyGHrz/nLB6rRY
RqhsPOcYbrrxPRQHBWMhb5L5PxFATPun0R2NfQPUPPglka68C16q3GzUc2NEa88FYoK9NLO7ReGP
fHx6W1ojhJ9T/RnHqfJH7XWKiaGqAxaNajEzhmoLYJYWEXtUPo4zuTYLfqdkQKA3LPsGNaiTld90
+AOiFdTrgP2hU2CBFzUGz2Y35hiP+l0guISW8zf9Hanyj3wjghO6HLc7t/ItfvGgUfoXwXzmDvkj
t8ZSk2vVUu7WU1fe5YhCDD6P4nQQHCuOCqRoxuSvDZaGMnuHLNl7bIuC7H82eVO/e2tUnzRHcruC
TSYOtIMW8PBRtms8E7UGRtUkS3r+V89znqCbwdaJMej7bla9UCCYPatOGOow4KveZtFKF7frOrv6
TD3SuaG2ysvtqEqX5E+6OFQmPV/uawJNUWQHBBsVJa4qhe9i4sl9a140MZloH2Mt6pp6iYZmjs2h
WFP5hjCdbWTpHGzW0P2t5f2TAaX9O/5Fe9QfsF2OScj8ItSs8PQCO+DvAhao0ERadya2nH4BIyS1
0qILi12YwMhiRaxNgbzuZumZxbuyDAEmE8VE9H0eeMLfJCGRPJk/5e2vOGk1j41DG8q6gzQsHc59
Zc0VjITU9jil0Cxa4um0SFncPJg+MU4zwHfX2hxFzBoL7GjF3ETLxCMyOv3wFNM+irj5aKhmyV4P
dwcrxE9Ox5FZiWJsYeOi/VwB2M94X4q8GHg80rTYYwxNf4zwcOYAnlOy9G/QgUYf4eGi/AZ1KDsr
OlIZ//rJVJuReSg+0NvDT99iQ53uPSr0r5a2/oA5EOWBePAiH/x39tDrRV9g8fNI90gq+jwsVc9L
gsG9JyJKa4Ar0qVTskJpr6KgD2hfpdWtAlvmOVWTvZeyu0svh1LsBQ94tIX8LlpLrZiL+5EfAST3
kBxS59+Gn51re/vUmx40lHAxTqFQYxWP+IhlsJAHBhcpGo0enwoI8nE7zMGsz/wmV37D2joe58XN
038N1A2KGDcegZhtckHDBSQ8DfUAPLM8ovsBBp2oYD08A5IwvfMZbfuKFw65zMvlJMhkvGCzhCIo
23pt4xLgI89kEGeendIXYED5AAkbKH3Un59DMtoWsCeh9+yTFKPk4PiUMsMNu/2pGQvHF5CEe9kE
AoM4OmD864GRcLoZeXMoJEp/oBlfclXQyiKNuk8cdtQe1kxRg6yiH39eHFXDql4EsqZ3GuGb3u+s
q7zE2FnBUOV7D6kddLlirJkHzS8GrC42//hjEf7xHrDPoS2EwWihW7s+oTyTHbD/SMQO4haz/0/M
gn0Eq0T29zvUv8NX+8ok6N1YESAj3b+kcgssgGetK9I4C7cEuyXW7bJz5C3Vvq3oIoEKncna3k+7
bXxLX0ASwsdL+YGaMKpR/ZtQGuKekCMicVhIfNeJwBn98YmOZLG/Okcoo6BvfX4rYk+z1/M8LXkY
sQZ+4I6lPhLr8VXBWeOZWGNmAFtecnW25q6Cs+d+h2Fjj7wYRC9/ONm2kBSE4h90LPWBMpeg3Jn2
8wjOlkcQJzWBdodEALfYh4Xf0SyZztOU/5ozVqjh8D6HJ8I4174LB6Oln331o6OhhkTcyH9XMQOI
cJDYbwhOGFEWgbaYOmVMljUgnZDgqyykjyIchaZtEzdO4WF3tpc5d+KIBb9bTCIHWy3xtIlkPNWW
FSMAqhwWbnwFEC2BJBL+f1KWX775DNFhSx0YABgSBeqPU/kUNr1svwfakldedJ9c9X+8CZCIsQyv
obMD80SpV1FqmtlGssUZbHhTK8B1ZsFLGOKuYNA21cr4sQ2oK/x6wLGok2I6PsXW/xtDWAuV+yAB
5ICxasGR7VLzDEOyYayTWpPq3xAUOW1TN13C9bMJBZ5bRF+j8KdZ7t/dXWh9/glhCz3mceildiee
zK1OMKEHh3ss2Ps7Y4XJTWJMpctflRNh4jcy772pAK+JarwAmJPVbLoGoaLcQJ/I/cGhg1OAWlaa
ue1IopQqy6J+NMkcJxHfOmjhYKTgrhIei94p1jysYegXkVKk+ItBriRcldnV9UD/Te/8uqVud4Dn
gO84qjTHbhHaNxAwKlnSSBu2dFrWB9q0PpqKtRhlCq71PnfvbGFLJXpkhD8CVttBjSh0DXSo3VeR
nWb2EUyzuk8TSBeAjdOaOnJuyMuwTmp6ER0yXjft+wnC9tFhhyOflDb5IT5VJGHm/p+XHCHTJgMw
F52XYs1vHwDYWO5RSbEVlrKeaJt/Gh12mqghzPeeFDYE4KotB4HFS0R5hbaH1F8B9+ym3cGt0fEJ
e5MFLrxpjsEfMhGKJsARbSsqh0eavM5CV3P8f0yqMSwSDNHNd1s2FaHKErua1ruy5XcSmrWjl6yn
y1i3UCP3T9p+RkPfOLr9xqepQvXf2cAxhJ5T+bPrLL4COuJIZFfe9A8cdRODWx9ZBy7lE/rwOuo7
Tf6UnwXr77Wfb9412PC0d6x+uNLiaQPi5jucF/tWafakUbxUj62pEIcKcfdY9jhd4IWEd3fqRHr1
gxrcELi1rZpi6f7e6NRIVlv5cBMReXoQDaXOQsoiXVJlAVi3UBUsVPLeg76SD3YKhjtw5+l+Szze
NF/8v8pbp4hQEG8Fm976Xvo6c6PANDvwKjHfUZCYs2Rhpo93FaS1yTIBac12lnxY8JIq47IRgtnX
FhgZX8Nnrxi2SkXQb6Ne7E2JHQc3o+rNyCuR7AWqhlRoGNaVQ3eHYfrnJtXMVoTLuCbZaADOajE1
0o3HVbIjiRPcMV7tkzhzq7Cr5LVr7aT12TwR69M1bmP9mi7ELLxAo55xMfKb6c7R0RSyF6PyT/ev
xqxlhyXviQM57POfcOuZOCwHyId/Rd9UadcaOapnIrVcdGxRjHy29pb2aclcLKjMqVRkzR+ufDHV
N49m88xnRF1Bhds6YZNmg6RSS5VEOCR0s5EcY94sHOD+LJFbNC+zkAKBNfgsOJiFZSmFijDy8TVF
x72u+OIJDwk/jKqDyy3xab5Xxs6qwlhU+Ee9ayIbkdFXUf5Dj0rzcDp7kZzV+bAzrcePegVTHGMg
uD9H/8XcrPS8B4TYa9qPaHAd2vJ+4eBqekMe2PFYQ0zBb/kT128FsOwwsUtuV8pHZMle2GsVsxuN
K/RhL5sZQDm4oFPDR6VNZ24wlqNMGu/1zN2ywM8ltvdVkno7ZwRg2wCh65f+iHAUsKMsbNiwP8cU
9mvk9plbBLpBadBbfcJ7Xm32YKVV0a1N6q3U3nzSV9Uidz13qshflrw2bKtsWNdTfcXlmsGSRpH1
tytg1FGn91sBT3Je/cYZar2y1BkENxPtUICvg1iWeJ+rI88grhgxnDK/D5qxFzS03LcnJsfHZu8r
M+ZEtN4KQ9L6kDcdH/PoUnUmmk84JdxDxP2llbs65V5nTfx8X4nAdZgFRrFT+P6/D2s9v836+o1b
gyXPOuHItRBEgIvUkhvBCGRSSVpglS1cxK3k2HSVxx+JtNQclf9VgVj36AabeiLTgYdZ3UEKyZQN
VIfvAnlMNKf8okyL4SnilhoKIbxSR00gPQW1mPMHDuRMxpUmO5a6t14QvHEPMSdGFFqTH1qZofne
VtbcHAGe2D3GyEa3JOCewkZmv6ChPiIm5HOJmQ7u9eADGPvWEr0gFr5ZAcBoorowGiAPd1M5NwHN
wjWDPcmzFlvqS1mEsRaiQXYaf30ga0SmEkY4cpnHxIIE4nGlloz8eSXitJfvynDrF63B9cBx8M5i
ZIQii6spZ04nx3/GBRcz2bSCV/wMo98ZhJ6wvyVXDq52wOQbQyCjkxCShNgCl9kuF6YGrM9J1eNm
ejg9g5xcCk8+49Q5De3dNaODUCuMu+FVjpcK1GwPKNeGqX1DGr9Y019L5gY8gwCq08V/r+W6kFjZ
iqKdHHhA5kJqeqfc+KdkpNhPS1HGwb09ieHwhmXQOZvHNPU1qj0gzytGqTeySrIHTvEWxxbbDh26
aEW8xczrDR3iPNEnJXvCFYzXGjCb3Yqim+v0iH4h5qPxN4bB+kvit/46jxSzJJCzdiYW29bn2BTy
M//S9yeJeO8HLXkwpoA4GdUEeVG2goR4qzuXV0qfKbxqzRpUpXQsDSBux5gPmj3+JA0SKSgvuIFu
7W0Oo8rFna61Xs2uWCziqCqstgmOjiurmIX03VU7UmwQF/Xo7clxxoGOPFbH27Eslb3jsdMxJThC
okS3RjrgAUfMTLxK2wZxPfOor9nwpeA8PlkCTv/B0nqC/yQOXWdmSWCYYKjam2pWaVv1/H3B4mLK
u4Gh6ZrmXXh3LtHdpTTcEjMJbt6ar7ojZswrcts+OZ1wC6T0DgmXlXzy0o0gRjLQ7rAqDTxEglK4
7Q7pikVR3JKVc2ih6PZdcD35noE13QnVEdxnzj6Wx5qM7beAolDlYRHpGdhmSatHOK73OxsUc0X3
6/W7E5gODcQ2hoV1u+JDnsXhxzZJbWOAFSa5+KRriMJIili8FlGQwA7bgSGfsNgeVkBzCYk+sUs4
UqkZDu7okSFXo/VnosQP9Vtsk27fGLuPQPutW2txx8fEliiUf40JwLIeWczbZWHnJQHPubRjtrEv
ow9opbxOxVFlcT9O6Xsjg0uwXrCBnQrn1YET1zv7ZBuEpcZgBoJ9X73eFS2NFAp6lV48fcMSd07d
nNAk6jwoJ71OFKDpKHpNNhMYf7pqBnh8ufqk008MszdqRPTpIHOZk7Kt/tkn1m5U2wGQh5Baciz+
2vnY1HGKG+S3fSvPQn0hT2Nd2emir5HBqtDIDQWSYUidLOuG5E2u2kSeCwLRBruEfbQZ8L3oA7aG
eQAoImDv3j2TSmBRHQW+VKDW9OPd2eP0u7ry4/4jOQ2q8HlffeIq3zSlgXfmdXHQVknlu9F+nPF1
LAFevLxmL6MxK5wfcGqc79GvDjEJ9kev2ES0nEKaL9tpDhlBXF/GHFJ/1hIPDjEc/3EWw0DIJnjc
n5DM5KGib5GCeKJz3zONa08Fymqlm4haTLJiNeE4qWGe8mJu/m6na7EjdQtWIxXY9KjzHv+pc44q
FxWEnc/TjnBOk9xPhIGIBB0xpT0a+Beu7e+XqbweDzPvAyu3FYxS5kzPfP0Zhw8WhOcI7NsYoUql
dxTuUrzndrTRFryw7Eu1YdEd1zt7bHL2XqQ5qWpPKDnX0Rx6dLuT1k5EPjnwRTQzJW4jOUHpwEVE
VZRIclMEbQKLXd+EhVLryK8o3K7X31/dQOI644I1EXeJ39O8r+y153mqP/e9Q3d4mvnBFeEYKR+m
3Swsh35ocXKlKu2NKl5GSQTDcbaTlShsSeTsbtsEWZ9ikblpxgy0xAwum6vLsxPtyPZtqajyb9Es
uNV9sC1NeNEiMFzhk3KQ+xfuIiDaNmCGtEdu08rhEoSkXPnxzPJK6+8DicO2GJfbCFdJ75LXNexv
Tebdu6KDaFAOGviTZuHaciTwCF758Iu8ZwPqJdXVyduXU9Ivz7vbfB+kJirUDXcMgmkQNV/xbW3t
9M7b+PBUz16kS3AC5COgyHqdlpee1F8uQ2vVLCcCm+GmVcIcxyuGXksLMqH1hAg2ouaCS0oB05s2
ULugMkEiksx8CgV905Nk9QuQclvh1cI+PidaSk8duEv6FwS9hd88jISKg20NJjS0NOcaCiPcfREC
QV74i6zFtVwPbgXUnDg3AnQNm/KjsK606R2NEmueyfWHZjnAZm9DWBcojCWiWOJPX+9ew+WHO/3y
iDfhveY55wONG8EHyDmOnfEyg82VS/E8kFTb74y8hqfT1BhVsbxNXGgNLu8Rmd2PIJS/2jMFYZmV
9XleY6fBKxVMs57vhzd4Do1vP9sZiBDdU/QrdfANO8zJOhBIbed3152E4zM1I0M9u7/kzh7apSP8
pkqvuVBpTfoQGtHU2DcPgseH3Pa5PrbCuNEnuEayfHKEzW7lhAyBCWmGatDm1YYdgNssCkovRKv7
aDnFDLicW7X6AKqEa8m2g5l/1WZZnAe0wrZmaAJGqlYozfh8q8shaVYh1uyBDNewQ+2wMuc2MJO6
fMJMoycr8ixs1omRwuqY2mBFPTLqgpNoNgZaO+WUP7aQc77nRedogV87RHMTsweV55RWsy51Szo4
bebOALAOG+NPT7fOAXXUKiPF9uQuu9SQDcrnzVGVbOF77zOh8uyqOLD1nbAj9LncVpDrjfqKtzs/
5Z4C/ou6irFgVI17SiHYpukfY0T3uGOMDmP35M9mEXSClDN9wpm+BfvHOTSzDjpF6Jlc66wfsZD5
H5ZD+adeJqnKRnX2oqkJg4+vldFQqzqChMf/C6VEqigJZd7hMvjxYYPhRrkfjR86dtLuT5hqkYjs
L6mWKjC/tpZczoObOYq5Bnt8kHqa0qUFmwNEBsWdhMpYZ3RF7wEqmNro+Ze+MObK2eXo/FLC19Bj
pM8InmAm1JNsIdJPMjQJoMdpJRMSGIQp9T7oBJTLVc7OyiUZHusBm3dbZJ2drejHccB1YUAq6lCT
R0GQ2lvNqgyrZI1BvPzA46NceV68oZZJbdWd7kW7SxKl5L39se4y7S7pcyoKwT4U7C5/cgzY065y
AI7OE8NPNTNS/E3qt9VuPA3Tq3Tss0VYsxLOaCCaE5lI3yvMZL1GznpRL46IdO6DGbkQfHIwdLE0
P9QN/Buqxw5GY8lkdL5mQU/yFf2bCWuFdyGNe518YEYDF4G8GBke4AUSJmXJJTPGDrIRg/M70Q6T
uvFebUX7QdD7qIAWwAQEuhpVSi3rh9TAKlWjrA9AbssyKOaKo3PXLqdwBapPC09wl/wNDhI4YGXy
384GcgU6XUGIP2mI3pK8d+R4IadttVSNJK8r1CS8dhITZLO6MPrQ25lwg3zRtvrBQBko6PfW8B57
7CAj7A+S4B98kvu2EE6eeTTkihSglMwiwvj7bdUag3eNG0tbmwi9OQM04Axy1bNe3s7zqN2o5jP4
ODOKdZk5BXun9wJ4N6f+xTaRoDMgsHmFPjmO+GEMYPNvJLT4xqNWKUP9CmtYLWckOaDOJoVf8WL3
ZOyrUFqSaXa+gV7VN7rFrGHa2LjtDhGXUzXTghjDCXSe2I978jyQfhUM/DGc2Lrg2Jt4A8bjuznm
zfrhcgmy2HPd4C8W2hyA+Gd07IvR2wIP3XqGzzqjf+yvPcAGE2/ahfHwxIkgsPWVTjfEQUIwd+MW
BhL2fdvFgFJ5J1OOpFF6ZDhY5h9Ta9yYcuBp6xzaGJKBjIQuOOBjZlU0hwrTaUcJBi/UQk0mu6yx
W4GE/es4erBlZx9+G4dC80VvKJGstZeqFPE+Gyoc4Bv2WrkQVFO5UeG/Ihe0w2PYWx9UeZqmBT7X
WnWl79NE522mRhnZSRSMSL3UofCiBkWm+SQRssYjAzqWwIqtcY0KYEutGYCXNlADCFM5jBKdKhA+
Ko+FtKLglcns6uERHqnn65TT3fT/NhBAIbm4TQBZ7gm/4U4rERSpEtvgSaDKx8GzbNicTaHCj0Zw
Ko7l6vTIvwyVbG7kxFnf+/8gCr6Q6ocieAMNFQotw3/otZaPnXdEafAk0zGaJcqqQVbmd/moJNpW
1cB66J56FBaKeXqrT8s0AjFGolfaWYaRJ8cEw+ofBfjP4YMyzne3ERoJbJ/b7opg/u97a2zCmUWL
TNmBLKp830YswaVt2pTEmA97BMbJYLLMn8aZS4ma5ahHJQwjKOi0cELwfEViJxiJGYW2ubw8LjsO
VBjsCaw05MA3/6hRPCg71BYKVZASBY4g9eltNdvnmbwV9UnG8ykGxsm7Q83aT3zAIFEj7ePwVLUQ
etRsEztDcbBCUGjVX5Oam4EuzaKRYyqAv3sIydK9no8vjFqhflTbs90cCQfNEfykVOd/e1yDsXeP
eXrbbphKnHDack/uTtzsdOWCsLNThu2zr+bYwS2/THPYFVhk19Z8BVpBdbzlA5EqTHgmB/WezS4P
AgeZVVYSE+kHm1dJ7j9xDI6CEN70zj0kUC3rd15FLH96sSMmoN/uFywxJF6JHrv8t4eAslRENzQ/
XZhI73Dn4kfN7dipn5pCCOgZ9/9ha/JbeY2x9bkgGeMsiVUHYPw9txJ++s98BgEwxM6uyEAurvlJ
PMTHJXlFgK9sZn7cxHEKaA/YWRMpS/xmzj5+70ccoXyywV+JAIpJfVRL9gbFh5bDU5aOiw+Hskdl
9v9bx6QPBGmVTMigKwj22ba4ZjULAJ9NBjGMEk4jcxIiqgOW/WzEvAy0ZCerI2ioHjFd+6YzJ6mE
lPfmfS8awBNmE8bNUxivyG1Ej3CTmHzq/d16GxnVM8fbKcSJAL+8+y5AyzH55y1xng39+NczELqP
HhoPLFTwUcHjlnxtwosFmesn+rjmZoHk4hNpDOxzO07ShhFFgOnMmpz/tEfkEXhEAel5Us79y5ap
xOVGR3PuE/dyP0V2+4r03o0aZHSQLFCgyoNiHGbkwqOl8dMT7Rcw5AOA21jYPRHel3yimEx2yejM
T3F31rw/MJKZVHkcYejMJKnSUoGZhDYBBpD5pDhygyT+2R5IW+9xV1ImE2jZ9KTMEUqAogVZ43Uj
hOt8wdX3qbJDdK82P1WGKlH7kxfB7Xe8PpkUK6ySqQUOpG5D1qlaYdSwRuPc9dPkMGwMDU5k+y0V
Rn0hKWJOF4aeBycvnbHvQzUkFmLhEae5XHBzba5F1f49OKcn5nHznk/ZdeqCXJhqN3oMUmHRYnlq
oWA/uPtfdXZGqxChFPl3V0qTY28TtIHUey6rm8QdFc1O4enaLkELn54VcDod9leHiPDoF+sjYef5
yPEJT8Q1hXkVTWLwj40wrSrOoNQivPDbagGyRpKzvm7QAB1wo/1sq64sKyv4IYH+PT6deTyZT7MS
TctuF7nfvvkayOPO1TiXsvFRb2uTRDK70dsTjjm2CNtjwU635tSbfPtDkAuQZ6azFE7KflokmKOu
y5xq0noeRR1oYkYUYNTKc/ulsVf2lTjTIy+4HCUtzXv8HT6u1qQ/ALHLhHn5OYpfPK488biLCSpY
IvtD7BRxDiDMV2zQyFKXqrxSQTSozFP+0GKtsIKFUH7TDc/gGQeUn/6f2zIYGKB5M6Pj4ViNVe+m
RLkX747kbtwwPalNJ0VAmZjFVxtRk+qPlkBod/cezj5/bLztNFjXf3qJNgwFgno9cvwN7N6R9qdg
wiqq7fSYWbWd9xv7oog/oIC/sgElDt3a/w+Kc5G64gWJOIiN+c6SP001jI3LGltUSls2ocDwS0OG
j+VeD2PntDAIfmI2s0EUvJmNsqh0OPaUghjRCbTXg/+EJprCB2mGiqu+/iOqnOz9GKsG2mc61kDI
ebIIMKx+D6hLdUlZkNVA4WoREapAOnVThTmYsaCxNEndXpCDiH23gw4XNWJngTqV2hZeONXYa9pr
tGxgaQsb2Yztpsp89b0zTXUbWAIEBZHnNohDlRMkm/z0YE2Yo5DQVz19+kGNixu3/xRhhmvp1OGe
fnCxAfJZmA573P1X+0eLr0zS1yl0pdAMXHRQciZLozjrcEBHj+H+PWnj94FBdDJDoYE/YbIx+xyv
XwA4k8kXYTmWzw07V5oPpOt5GliJMqQ+E4ETEzVd+ajopY4tb/v7lkVeEmNc0Lrr1g30fCWxHQMT
oiVCRs9/m+2cvpxzP17VzbX0tefg+L3UQIKCdf6SBmD0M9g48MYPih8xYOLuT4PwTZNTpWgzRCcZ
DTOVT5WnpHtJkBB5C1fIIR35efzM8PTUp/X4EcqFxVnFO0h/ozJyDff4ZA0w9w5gvEz1ifPnHdap
lUZr8bllClJxK3n+w3tsHJ3nyRkQLOh0akWuYWxcbeptw0c7GrWeb5weAEpPRe33E5zVgtmKzl5k
W3vbaHCW0uqN6eDzatG3qrTiN4xvUugRFD6db+MTSWStxx3c7sjgCXdvQN0Z2jCZ3QmXkyYPrerG
bzDRMUy0pTSUp0zI20XIqv+bs766ucfVQkKu6xAMyeK+CDdZ+GHc8XiUTH6HNi7MdhZSM3cBg5Ud
TrfVkRjNXmSV62dZ+jzyqrBcddOfQHuscOqVMGokkktPD90nuApQkO17gG8bB0S8wDjNzCq0n3eh
RvVowgG52cucCLhpzDRZrDWOaEgn6bEkKMdVWybQxzC//ZsSYfjb9Q4SFG89qnBnLZ2sqNrqjVnt
/iQZikektSx+q83MFOm8bozzgnVHPwJGSo8feb80zEi0sQ919bt0CZTr7e1PmT4/zWhjVxTUS1tb
QOZk7cJs2i7DtPdUrDNhfBxLXUQcyoy21PIIyLPWVHJKYL2R5yp9naF6n9tlmurwgZe6kwDrIgNh
hX7FX/yCjJXtIbh5B2FWIbbQ1ikUnx48nqF8oKNNt49jVRoMwOSWli2YBBUbq3/xfdwoJCW43kck
lZyXyQN9bUEXeoNE4v6mvd3BDHntv1UI07dRGCRPp3DoWwfBGEvyBZIeIcH70U11ZgA/zZCqwzLo
Mp3V89NBarWW+xWIwGEKZgQAPnDaBoXlrQUOUqha7rmXYJMxzWRl03SyG6qNkjxpdTaKU54Y9k8T
AXF91DLfhk6ETyiNyTcAdRzYHx/wE6aMpMzgOCtBoklNozDrrPNjRNMvp35w1ZJD3uDFvg8LkI02
eyL0vvtBmdT2MA21R4r3vG0CP0HWTiwOdk8I1o7B5M0iDpIfNjXErUYEpfw1N7VmjglwkFJ97EZY
zVul6yr1daqYMr4OzpLho2K6dQj/kVRZnEfJ5p/guXtox8RXI+4xvCGsnoAw5RJoQoTG+T0b8Sle
5kg1TVZEt998BIltAIw2mjBmmxGduXSzOpWhZfuvnPPu6kBIb6XmERtaEKIKiN0vStR2cpZ8lLhL
lKtnfUkY1eT51vg9MDUTYqowcmwPCOEctrj91QgypzHWNClqqFr7u1R5YDk/WveF82qA93m6+JzH
XJX5z0kpjocoi5Ya5eC3AeshnMF+IX/uixPqS6iQZlm57LZ7k1ZQt7brLoyFwElKessaX/UrZ9HX
/ii8QQHapGClGgDvx/UmtMPPbt82PqTDhdXnUC6JfMTAD4lAz7SVFmby19rpesVtHy1ctsMCEMlg
gvSwa3eQ3Qqr1v34DeI1YwhTkFr1/rpOheMDjnwTJD7ecahDlbp0NWpx4kKoTwOEbVUezP6C8NdZ
2KSEiv0RxOThgbK1OmQcKZB3gI7AJDd76eteG0AMFbeJAkVwodoQxY2Wza8ouF2EAAnZQ8LJI2C8
FgmYygYrA1fTSBFMUIVULXjqotffRiufLLhcthjkPt4TU1D1m8a1UBVfc/VYraCehFAMJvHLnGPl
1VvBCbAx9YNtlI9FfqBwpWssqIa+59nfNC8Dsxnu5NXCw0od1uztPYofIwZP1lcYhmZ++GHL+hsD
TlrCIw39MJ+dBE29mrqtvrEmrOlCYDgcaKptR7YHgcotHBXdmf157a11JRJxCa7AoLs26ScBCrAJ
ZV3DW8GToKW2BYpE44hA6j6EM76UBY/KpKiriK7gnssOSg64YP9b5NKY0b5vWhc/Sm1/6cUs00uv
+NRABOaK3bT5eurm7IMnWGi7AY2WusSfU8qNmUKGsOdOf2zoiCngAAfUQkb24Ah+zVP4JwO8AASC
MXPHKugn/fGrby00MqiPuuoF5CQC5vdjipevG5eUy3A24V0PxQdE8tn/Y+65NNOWrE6gCwTUQxYD
ddUwvaoxaja+qRoqFLOCKuaIbWlTVSHvCbom5tLgeRknjUsbZYtHWbmyjpwNCP+WaJfts3kq5Aw0
vfWmM1YbaSMRYrfTFGoMHPS2iE6fNhh9OmaSK+xNgxxHjcpfTqUUSuu1ReVVzaI1JSoglwBx0ljG
K9Rmks7woBRIVgOLEz3nua+0LzARteBRNIpFIHOK+nKdQzP0BKL4hF2diHVLmJf6qIivYwyOdHze
aWgOy3WQZ1zVwEQ313sx82RlNWOpGKbpkU9t67weWMcLBcFSsz8/w9Q64UfP9NzAjb9dOfqItXc0
Vm+UVKIqCDnjXm61wHaK6V+UX3PhfcsubGy7BZzdtx0Hv7ZHvqq1r5yGtV4OEOMLqb1PE0xCqP83
oHm73r2U95uac/AFLUQheijgM1S9CG9TH8LhvERjyHwHUompKO5SHQQBFULsodgLSpNnLwy6Nsup
ymR637zxnW6fzFs1MunrR7vQRTMIrJbLdVJbFDPNL9QPFJzp2gsmNdoHzbKGiwEtmWybLT7H6VQ9
r8VfMIBjbSYRJBK24cPxeUC5Jri5JPllXv9MXmwS27QB7LCpw1Ag3waCvbEELniYcy/VtuffyQN7
UGHtb+xLtSD/Q7QSo3NZUh4UREF056MGlxWF/a4N5oPihNH0fgh62AyaZmGKwizBV+N0VqzGeCmX
78UDaHncxdCJefxfcy3rLTYVEvJTieXYap5oKasxMbXVjF/Nj7UQWVPzFoMkIk9Qe2WEp+/gRvhc
dw4HUGGg/EGkoXIyeluks8az8oUuFx44CvXGXdJJhiSJyzXJDIwo1yBrnpyjxK2SHO3v2lBCjLsQ
UQUF8KWEqU51qGc4zJf7Fhqvic2zjdionL2RZbCL5Xshak5JFaF9T6Yh3KLDVCasQUgj3ZnigLCi
N9NZgk5POroeMUR3xR1LGc7ftxpvhYkspYBY2uVMQOkNdb9NZwWpvsH6Gzn45KXgyl5uXtmcBcli
bFmolwnSlVRqMJ8Nl61simw+P6OWv3qgDLK6Bcaxw8jLqL73yvkLmhsSKNiQyWT5fwKcLHSXqdSm
GbaSGAypIchj4m1o+TGDrddGZJZCSJM4mUfm6TwXUCWL23j5PiS4+YFWZga5hql1i2zD1Q4TQpto
VvHNw9B+D6iXZ7kMrC0LvAZS0gKVgI19ccw86INSl+F/qf3M8r1RoFfZ7SgJVboshAIdFdo+A4a7
46L9EMQh8u52UGug1tl1lx5tXuoMK7hh548cTQkUlP89VEhPiUWZGIQOv8w5BPUR2pRDNpkUEXTc
Yt+a2bmx0OiMJ1OdfN0Y8bcUPNuxF5nwFX/+mosMLbOXb+WE4Q9EL3H+yaTZxqJtdH7Uc8s8yRVM
bh8jXFkKfWnl4kpYNS5RqnU6fMK6XGeFlbhErVj49/kbZGMKZ1wr+nsgZfVNzDyR0uA3d6igC8Mu
/rYOEvh3tKM6+GpaCVNnic21dsmS2/sjy1+0XpPi3z6Q9cQmMwEokZbDMrlhRVDowsm130XUFFGr
6YxyNIED0ne3iPsFLRXEos1qnN8fBmmymXQiNPxFy0rTjfyGhXnF+ULRiUqA1murTR4px5Jf96ew
08MPIBGtxINze65CDXSUpCGuh6mvZYWOzfv9HF0f01syVT7+w7M04l2Z30JsabaO1QboTOiHDs6a
Vq5uF+6SMOx7lbpygaISKVXxRLu0s3pPlqRQjPXk+YcuQzUBfmM14ZVNu1tEpbKiXpwEoLvqYcDB
cuppqUTAIGD1wdimw2K//ZfqeCdMQMHzhX6ttN4xfx11jaxF20zkzUuWTEqoiUrZnKl/xWGodY8m
uMMkVogK+AHZVmz1hfCbMBSFdR/4Drq1RPVRr/2GYUk0ONfK5UVxB2h7RpPvXFppmlB9Igi6/s+A
T59wdF9d6LOffVxUvtSF3W+9TCk1LX4TT2mKAg7r6IbmaBhvIkiLs6d5NbK085bDqHHPLK2MlZWL
VTbu2TgudpZVxZIgXiWZ7WFkQ9pM8LG/E0/E+Y/jqBmkqUfSrg30GeOCRLKqAyxXqjhup+VcUk8r
RSNEzhfMRHrIoAV8K7E7QmfsqupM9o7YcFSpK6cokipEPWgmxbd3F5yV9+hYsGlmbhlnufzTZh8p
DwrTh44U7ja7yNIqckRbcYGob83kVru7SkAf5TyibPLwk+RqMcVOFcUyxShlrfuoRj0h02bh14ur
BnXrgX3LW5mJqyI07jIrh8uhU2+QtjiTaluYhRJNzQ/S0tCYGnq5KI6yHCjcIAfJwzWhIegOisaj
aH+aikxfSKAZ8ZaV7/xIWKlDcCtMe9/h2Db1hzVJTTncDJUY7hlH5PRBFA20PCOk86NE1QUY+eoQ
S6+XHJP+Kk/mJekKIkIk4ag+LYwlmOcaKddcZ/3gTnW8GfB5xBFc+e0YFpFimiPnlRRV0E5PKaJl
iwWSczqHXrLwX65RS3fN9UgUmhIDQHCcg4LIv9Akob/Yj4yUAIgMJHB0Pyu0XQs6FXBW24HSLWhy
q4tICvsgU9ge4u/tfuhHctCTaEI3GMSwaSuBUXaYOOQ0dc0fZKMf9izMLsEeEocu4YK+wylwQyZb
v8Cwvf0BhdjyjYFaCvkk3XtDsutGDlKYh5+hcDjQui310bhGUbXnL6X27c1OzT5OyBTCwWJr7KJK
alvhMVH5m9InwXE6Fq0gtxmd5FDW7X74wnx30l42tqO2GViRWdv+jDY6P0NtPL0p7s3YpChUYib6
7YZSxn0uCLG+4Af3ZyK8hZC3WiXpsVXp/tnAvIJf8vPmstYdWotFN2vmpqAd2dVDsGhxBUAq7fVx
rdH0FFnn6zICxarCVBSQwIK4w9i6pBNREwfj8iHlYUfwJRTrVz/zbOVi+WSAswR/QGZPr6HP4fms
gJasQPfl9s0rwc3er/k75GhkYixPYK38f2RHF831mGBaniSnVd7qkOFvD+OC0a+EN+8S4kYHRWyo
/1Uc7Nz8CYPEa3iMniaeTE/nim5ZMiLiYmeiUz+ZNEI+GI7XIqHkutI3rH9ZOctc9HhJfTYAr4v9
WgO87hdzR5hnfgtySD5UEFRqmhZ/+Z9GNqjSEs4TCoZIhP2SitM30QJvvv40IANUYuT7UAlGYkMI
XWjFsXYukrat8I0/fESX+bLphADTJL6XA7hwRcClp4TH5W+bw/7dUk6uktMhgoQxlPlcwPytlekh
McCMAAMupizaqwhL1l5iilxUV4SkH/ETfAw5TKcOSEehatkmQihLElaqjsy+in9SzxjA+i+pTi5q
YTDnPk1rg4TFy83MW0kfDR2Hh7WBqJd9x+7dJqfijpMhE9SsrLxaTA3M7z4bUaxhy0YOeHFO+7wB
nBRRN2aTF4m3bHbIVkgCgRXh96D3dQ3zGKfFyYHrOflBs2GEOyVHozX6lM+/Xtuo+Ljgv8YccHSB
+8P/4GO5QKBG/AXpsVtTdc2KkmemGujAYFEAIjvqiOGLLmkDfsiyQUfN7U+Xh2qOhz/np6RL6GVr
1rZjejUQPu3b8wzP2PuDbKZppajKctV7IoPpRTwiT4AAF888rGX7xEqCivWWJPQ27OP+nPUqdYnr
1YGCJOzMcQVL+P5i3nn+jZUkan3377P3L5I5FyfmKlpQdbVHqXgUiUQajx79CMjvGk5zflS/FzGs
paGNsTc4qpuZpNB9q9FORHLD74WIde3bCvU0ZvTbEpzuSsQ7JUqAqxixQj6M7xcBxu/Z3N5V1kUh
G9VzC/w0IhOlLLH2DhuBsRPHP6mWhkA0EoRBXZWnp/bHLn2lzsyDO5CVRBfH4C1F4fDTAjW7l0c1
nQEHunKuCVnOuXixpGBvnyT2cIDLmmdiZP+5T12vPEafdPgzknd5a3JEYjg9gA6yxcIZLv2Ys6+o
BMS9m+LJCY9YqDo1ODstyqFTvJCVT2aYFLL48AOtZ0ugo21W2lRAzh4yix77dxnkymgw8sNGL9ci
ngo6Q6jcK/KpreisFraA7vR0mBk9+IoELrhDCHTu8TCHX0O9e1AgONP2MwP4GCtVqTAEBWqH4M36
5uMiWq6Z1bzcAlYJDtiz0sZXGhGSKg/8cw1CM2QW9SpotWAo/FGgoRsHJFNWMVqV2zT7ZbNseBm4
OxQuDeqOnEJkiLr4BwL/4Mwl/SUu25uI3H0jqbBlSOoWFU2A9Bq0kgoKphRSOBe1/YzT17IyO493
fwRyc5K1CpY8XWv2y2Z9cp9VXfMssigcEOsrS8bgep4jl+eHUleiTHleQ/8mpKhrIwVhK+/mtH+B
r4UHpWZpimOUyvg9a/sca+5JYVK6z+/iY6TzRr9Fa8BiPf1/pyip1HKtWXtY6JXAepfyk98II97y
28UclcHAcPxUTdDoJxBdivropJZO6ClfsFOX3bWbymMf4LaCi8PGmd9L5g0PY1a8sZFLeGK20L6o
ql7ExE0AoJjQ1bG0bEV9fL4uKOnj+sa9N/ombAxaj73JQy1FOQEB8VAPmkNcb0AikofqOnXb5hrj
Vq4cOhiLcyFH0KLX2pr61bI1G68xV6BEsRHRuBc19z8xjrqiF5+J2OP0HhtyBVvNOOKieJBZCiCC
8wmaxijOEWWk+LY9iEGoTy66pilEznxfTXXXwGMdPELsBvNBauRV3CyrgDHD9yFuGHGy3xESlz5e
IoqrqWR39HmJn1S1P48Ganbk4OcLc6NFt9PlKrkFmEHBzGbR2sWgC++OjByxavEmov2LF7fabdHO
w3qHyK/aNX6XnPmoUohsvshubqbMZdBIyQhIOB98q7EwL6fRPXDu6qSdy+p7n7kEea/uZ8MxDjfH
uQ6VMip8m4UjNvh4G0xXupfyM+jT3Xfd1dOqgovycXURUVVkJ1i1CODPVwoThBsiMy5VPpl4Pgn7
bUBCxni8D6x30nRdmC69p0RPwpKQG81APiWc4nY7GwKjCAc3zrJFjnMB9hVUvpG1wyzG3dJ9g5uW
kxrm6qRVrhbXO6RNEdG7bgCiD1NLlnaErlIn/u+QDtsGEfpzI3WgZirqvd8m0R7f3iPQc2I3g72x
xzBAKgheSfEaTX4FjNGIkp2DWO691xz0dhFrbDQ/bfRjmXHJgnDbq38vyWWE6aw01ObDL+hif0PX
ju5+Fl8Y0JFbWp5HyoA3mPMDjWThpG+6RNbuIT+B6I9YphfT0ufrbPiJH5zsPb7Pv5u2v/bot6FC
E7cUzGCA9RMvN7oKiqgQRjih/VXcWWNukATJSi8ut3yFA7EwyPQoXU9AhY+QI/LruJoy6m5k7X6b
Z1N5dbgJ8l7uOT/pGy86S9VuHjWd9AQSnzxqPP9ikTqFbdTuw9th1HBpJkaGclQLfuuJvSl05XAZ
TsOYAja8FzbezDjc6tei42mEipOqxqjYLQF5VQn1erlHxlO3YgTmtVmLIuCDfpTaUC80yGrNLT5t
Zyg/q5jvE4FQciVucznnWATWv9hwRTTauWmBVJVhiRIxzZSAJGrRENVee9R4dq9fX+uryRrai+Ff
dDYap8l8dl+joFCJDIUvM1SJRb+rjSvfjgiXVE8CnPtbRvdQJxjtN9X49QYM8DxQVg80fdXNaozu
KfBKOdmpPIId/YqoA04jPmjxaUzwBu+bkRiJ67xDHt5gFpVsJcto2HAEZn9Ws4KjaBu+gUXoJp/i
c3CPe27oeVydMD35xqIFqe89/jqss0pfiM0RG07lrX8R+amSUBSkF0b8LDfopaic136uWH4Xwrdt
MNYg+OcFxGt7+hZa8rKhTJelmVcBwRfqrqRoRX2OLtt9RhsXhWSVZLagJSOcH8mr8C9bym15pt+S
X3U2llxS0b2YL/jj/ETLpQBydCDoDsoMNOY8IIUIcufIy0YmMxuBahD3azvKfUrCjY+CwKvbZbgi
/nB3KjKnL5wiwwSIL9wSLGaEFYMxTMceROr3r7UYyV80Y/Ygm9aL2bII9VmClLo0LMsHpBPFwdrV
dFgtxDk+jrjXfV3xbBYgYF8UaEWkJtpzsIHq1acv041RW5wXosCksKKB0MR3oG6nvcNePv7u99EO
BOC4H6BYsl+J5xgliRY8WhymIfg1gb4CnNhtAHaLDDMDpVZ2dppG+Pg97KTSIQFmmJdYHRTLUD2K
1Z1J0ux9YxA7lZH3D+gSh2aim0UjAdR2a9jYe57oAP3n0TJOAv69tFWZYVcZAa4K5OBYlaonY125
7xoCi9wu3lnqPuA3gwZgoMfe7aBUIJPylNCANrN8F9ULciLYAuMD7SxbpC8iB3OiitTjyA5nf0nM
km6AybMLtW0Y6rVmLpnvHLoB1F5nwhXx12F0lcxRrtAstRa3HTDbuTeNXCWbHqn9Cpw0p5NZyDGF
XhLkv/DirqDIkZmamD/vnX5XJvj4sRI2jvJMhkmRS/fiKWtffQVKkaHudHw+ej+VINyzCxBcJG85
mkBPjDJKTf3qErLoDUY+6PT8D+5aqwKlihgiM61NE8hxG+vxK8M/bGLYLBtLbWvJSnl53YFh70qR
sE8SJ762kVWGMbEXq0TJjQKFErFGor9RS3Md71Ci1Mn0d2o3So1j/SaTVlEY497xEtBzIZ+I3rhm
nsjC2Wh24LnC/gWwrtiBStlflm5U1liEoam4aI2WNshissNfPY9sBj5CsszBd3IDoSNTXvWGSJf6
BjmaUERtE2Y4KBiEKUkl4yi6ipSDnKz42VZkWseHFuOgYJk/f/5+XILWk+NnPOOGcTzEkU8fggQ+
6nHtshri093KghMcmXNOE2xPeB8jpkqy+vqXNZDYH6d0y/RAkVILbP8bud7ym3pWmVcFrNLE8Q0W
zJOOEN3ewVs16eh3GYDsvfdeVL7Tnvc/YauMtI+vbnU7/ofy9bHnHHWB8Ft0MNnGQafsWm5JT5w/
3jC3dfxG33d47jj0xrdtv6ALMZ3LclsUMgh7lE2f62zHIyZKEDWd2wPpKw/C8zCxyzXMa9IDe6Cq
Ep+uCEAmluigg+3CuRp+eoRhaCtFFWJ2vvDfTVyg5d5tmcoV6VrqAXnVOR/uSc+/mjMrtbruj76S
spXjWqXfd+MGOaAqBWnoa6a4Sg10tR93P6p0zsEBxFIzfr5rDLBg/L26LLMwWNgt44v6I9A48xFA
C5CWrWZFN7Dn/O3mSQxJgQnHcgBEVXRlIs3ATKmfx8ttXoPfiwtMPpkMED+W1LgN9t4QDRIzQLIT
EdJs7XfMHfIxCYsnYOpuDXXcLxXU7Wz0Q5ScvyxQnYqDvBBOZ/EeyAaagNjGTpdwWYK0tKQaeOwC
aIfSwYlKla58zXSRgER0oBclDW88SYSE5KFM5NXDQD0wEsAHUQxwKp2z7LiPMLsTCh4X2udiT6vU
Mck7dn/yEnwfj1kN16gvdz8NVrYvo2es6ByYbO6CHMk7ldhHpR0s6So/KAwwTTAlY3EnmGeyXE7s
kdOIb6J1FD3yN8g2plQ7x0rdCTGKb6swAvEnnVkEbI2zWYx6nRwY12eyaJCAH7rWK6O6+pHP3nhS
G+6zqeUU7ZTMG491AsqjGebepHMXzrDOa2Rs18YoiPkaivC0BmxZgy1heEY3USoNVObeoAfzcOt7
IXStHahOTEMZiQQ6btQFuG3hhxBTWd6scbsgYs5XhbUopMe4dQjvIbAKAgOc+sTsbp/rr9qV+Vkk
Tb4VrxYE1Y9uLE8Ha19+MN3DuVX4MWMQYRamK3GNIH0wTOrXAmcPTdIOfEtGY2WsBcxvgSVDZXzt
4KkGK/YBPKKcdjIbAg9QQ3o52st4ejRnmv7tgmg02QggW49PlbjPjT0A91lPzoi7hKTZTS49WBGA
frZPNiBKtJVisnzM3v+zDXoDbXQpONSz+b3TgY8ZYjwuNs3uz06zMBUK80oWJ68iAFi3+ndxIkVN
XLUCdbDoS2geiFcQZ8pAwq3dgxJF7j7NB8I+O2uP2y5MVcLp/OHJtmhXgGXL1lXQwBzgLI7PQsUi
rQXQbVIIGGPMGouu/SsLKodWW2YGGAKZHMVyHMijmykPMMd2XA0MF5BdgvIqV4DU5lwa9Js8fgFB
9wokgqwhMaeQPC1Se0MGhDn7Yfy+EcuxQHGtkKnhimNlOklB28piSOFW1xjgZ8KLIfhl4l5u64U6
Xcrau+wpNNsuQOdF6LQzmxIJjA4lvD/NNFiwQ4qERe058b7Vm7Y59iDBdG7kX1M9aoHU9wbdpgiw
TpUW4rhMfuYVmGWBJNxc1U+upjVMUPuXsNjp9MyddBk3hfD9e7JkcGbU1zMMTp97GRylEXqfvDRO
Mw4ky4sVy8UIj6jS+68rWTk6vaHIv8GiW1mJXu8I+lDXAQy9hyIA0sPSvSHG3sfxWwSlLgePke2U
MP9maDSyXitHZ5fvoW5JlZgmBloHz+tdevfni1+Qtydzwc7tQTcOCw47vsec64S8LzviF5IiXnYB
72hlvgJCmqTvfqdXcLcT/41ymRlY5KTGn1ROju2IWnzy4djhO0wS7vwvq/Fdir8djs2h+NESa/5r
H2tkS88Xn0Q/jxh0VAg/6FdkIouddHPc63utGrB8hcaq+TQalLm6pTgUrzOpG/oQ3O/3C2Om7mgH
ir2OZg/mukn2VrUjCF0NghbuI2dV52ybB23MbAJNSoFsvcSGxf1vyVdge1bj3DBCwGTL7dIcJzbu
yhsjism83BwXZPYXHp1kRa+ZZSu3wGNUNEr3fYtpOC7D7IITFZ9soIGlf7kfZjUGaeg+n+OgXcgg
cIFDT/2As4A5QO8KbgWdsn9EbUcK3voLeXkNtRVkjXUVFjedVHL1lFFDgh6W3D4YdMeYIuF1LMVK
ytd0LG6NXHuvHzsFnssEZ3xAy5YNzGiKZz+jhscbGsJ5ZqcZaf7I/P15gMGRmPGAEMsz4dBS4RTu
mGOWB18uMSDgpTLidQbbkD3oIugMls9Oc39TYFq77Up/CKa0xUaXfBl+GCS/Zvv2+mKABioiJEjx
B2HsCf4oHNnz9/G6EOkJ+zysRlGfIn5H9s9iRkKznAUgV/3I6o9rT598kJHk8E14chuUHNuwK47K
ZzAnWVAtl7L3lp4uZjuiJ7tFqQtsfPgvW1xCoRG3CeUSjHfRR4S6W2/MC3CWr2LlJVMFeHkNV8sO
7vDE0DvPk1THJYzkkx5468pK8ZRnV5i4rNrSf2giT+OK0wteH6Dfuyr43xAuo+JUnmgQxVlbauus
15Xd4Q231zK3IYVzPWlKx1sNwbIxFQ0owzLEsH3BHtMQliDNrZKcFQUq7jEvXTh7W6ffzKJUO5wO
s/AoIBtKo2vMrN60Gy+TRveLJOF40LYKQ/M8HofyBzWZvAtcx4Ro+kLgN3A8+DrYni/pvSHakACY
Pfdlxd7zemUOL5fHn/rQd9LcTobl7GdZ+hhYPGtCZVHHUJN0t8rnElk+kOQ2nO4WZq+KcDfyr/9R
UwwCApHvggg3ZuesSIiRyGE69quDTJZoLV8Bhcv8iLAw7WczZColHMPQR6rnEX0MTtR0l329HxHh
QLMBwO2Q3rBYVzBaS2n/138+HrX3ipPUDnGFhByJttXswhjsHSdhN4ILSFuw9mBCbAO949/m+tLY
lcPIZGbytnthtJleujTDkg5GIpQ1hoFLqRHf4IfaGAMjvZZr7HxcTuA6iRJdqtpGxatq5UkPjqWB
zLu9u6zncnah59P/jM3viJ1Eu6nstf7MYtXsgoVBz1OPkEzbb/zCGkFhzNs09scHF31IlG1SUj6F
hdHvzqapjWR7ySijLPo1JzAw/WftiO8eFERGqSr9200B0lptdXjlQ5nRS0zavRn4SaU2eB2OKqD5
8Mwgb2NNO2ATK2ZRt8+wqa6a0kfJbf0xAFO+oszMg0VIwKsXTgBBm2WUqlOnlHe8khO9Qj10vGSN
rVR3wdEsi2vIm+fpqatnj8uzbgqLa08cSLqUEaJpPfw5PMNWav0qI7ktxIikOwoPclB3ZfxQksa6
fxcp+HxfFc304PAgfLnKIkhHrMFt0UtCHluZB5XFTNzPXud5+Gf9C9yyf8/jSptkwcpQPseIPE69
hagH/jcjxgUmlPERQskiXL/YuFtu40GUp996qlZ3qP4jKCg0hu5B60YFVk5hdB0b5gFViRPs+BF/
jPIzwwNEG+Qca38bH/k/uTKrkDBdsgFkHWejz2kdzmI7cYyaptOv7RqrCHWbDnfFPa6QvpM6f+g0
16jpJj5LfEXN3vFy6Vhb5eL614PhPcz+8JV5evTvvjXeZsS/7yazPDlc0ZY6QWsZIbOUcR9uXbDX
70EjAUNvU6o40wPJ9uiFeoVynY3ALiS0UcvClla7n5rI0hV8PcTkaRUSkqIaefuz0a6LQnp6hViT
uG4qMLYnUEK7AdyHFPfi9GvYfUtrcVPiYsb04n8jE+NLO8WuRIyrTsIQ/AdAiFuG0j0ziSCU8V8Q
E+iCo6iGbAx2BvOX7gm560SZ9AJCaV3ivNbyniWfZETx8M9uI751hPUTdypR8ozPXwJ3gymWEMxa
8fCBhnn6RCm5DeB5zsWYf8bd+whZfqRBLr7qUNSYA0U87o/mSGcUSVCj8YS1jWdtzfNLSeJ6fyVX
7JBhIGUZLa3iKbRi005Uz5XMtoaG9eOEVmpwCIkEKhXJ/AXsDly//G9lnP8Arx3JinKByVN8IsCN
ZV67zuxvnY3v1gC9kJiZfP8I41JscAaLOT63F3+Tmk3b8cJxVpl1HAD+kDqF9NRhqVuulBOGHPnG
vvTfAZ7tYImTtlIQqJhfmwyCuaBBhVOYG089pF7g44e8BRDuItVK25ylj6rBS/tmZMnkHL0WIyoH
txyJvph4Pto4pu4y7gG6qtkyR9bCbTKw/vpwjVyS9+oCnDrqsO+DzZmY16wGw7pl9hoVm3lcxCDI
ETtB4VmshtOFRa0G3QNRpNW4km99LxYuAJ9ynG5U9JGgCjxQ1MiHC5Utun9RuxN1bbCPIcKcASi3
IyCMqKAz0vON6gMgbOh+UwXWH5jQKHuPKefGXm/POAUktAMGkt99GcxZzlucoRq8uxs0N+ZEPxCz
MqTr+baRTNjmZVSMKKEorlfbSaHbRypuaD5ZtV3zVCOJJfacZ0TYSuF2AIWR++fA10N1wRIE3oHY
/t3MX4CDbl+xx8o47MxIapx5KBq+0EUXkMO06QUHQiPbieQcLcEPifPNphQ4r1zQ3HJWDHs1ZqkY
QdP3p1shv//EwWvXpYCJeM86tcGYvOhXGHRpST0SCidQ4e76UEbxk53pMT3PIcoF2Bk2pBZsyLMg
sdS3eB0LHfWRXIJHLlHtA1WrzUdpj+jA29fJWxI41xv16VpVDWcL6E1oxW79Tf74zRDNURuunm3F
p9NKVOKPohbcCiQO95ykVvb9fS/xjWUIoCf0LlFO/UAlRXoNFZho7ray4eJNqExpB0VUyVrwXDDC
g+uOmjbgIt55bX8BZu0Mx+JMj/GkyLno8mQ+cKKbGIljEE154WWHFe2g/j9cbDQEd0vNvT6J6YaX
DtGxYMBnci5gAYGb+Bam3q742v068wLhyA4oUoOAm5zTdH0oP2Y7OaYKYlq9toxcJFWyjwnNTU5A
s2qeOSsiIT51kfdrhGO6qQ11pKggUUnUsz0xTfqgoxJ1AqPA/Zr9hF0JH5MjuJ/ObaJf/gMzEta8
h2MaQqldrkq4R9kFX3Zq709MpIwRmijpDEn8qmoxbHtlmrKzibZvTsOtVXYfDm62OWMAt9H7RT63
CxCqskYJcPW/DaA/551GPF7JZc2Qfzcai+BiikQIyOniQgPb1BojKob+iE7/hVrSFe35ZZ6eX/cJ
CDVOcVP/4DYK1LI2g9uu5LXzzW70DHy+By4G4gfrCmVMcQon3cpCcg5tbGzBHa9geT82s/q8jYsI
d6swSiM/7amNzJSkI0jRcaInWyvl1wuQKDF2ucJR6dNymvlY19aBWRGyQ3nj03+6w5ld0OVAPCV0
RWAiFksUTxfxQyufyssEKNmLof3EEi5HSO7yhnazlH/T/1x8Xvpbxt7TNhafLoSjMsI+j6XHL9xh
gZCZvF19EIBsoH5Z9/ywKgsUrZCyKlor75gu75YcS9IBebiLDxqt4AFJLKqMS1Bof+AW5l74ipzu
JPVZTHOCpiiFSa2o2T68VtFxIPMUEyIx9c2tGSP+XIKVEGM/M9TCkIod25rSsLoE1SW7/untR/Is
vtpUUcbJwIQCrUKumwH1zHICiFDgq51k5bElj2hoXUiS9UuyG14kbmz1k9gCXbHXqqrLFbGFUR/K
zVuwww+5KznkrYe5AKiQWmn8CiJ5VFqTRPxnEIO5JEOhcBHH5wiXy4Wmzup4YpkrTI9zXFPSbFj4
353kReEaMFhtuAxgxKEZ9P/wgqkXFZ0mNlamoX0niR8I4rXLGeEWVgRhileXYUwBCwW/IYqXzNX5
y1kD5LEd1HaheqbZ6Fr6PfANG4PZsiPIY0Xjje2ZMujuL260Q/eF4Eb6Zi1nxM9L2YLdPoZAsP4B
/PigEsuDFcLFrN7jCL2XJtv1u7hjoW+WLes756FWxtDGBNAQAS37R/90jNjuaZTRI54+R76+u6cg
LsMwQIYpPL689X8IzGzc4Aixl6YZqKbi8xVEANNrG1RMYxHPWl8T19PJ9YomYh4uzyErcIWC2j4w
unzi0s2yAWpnhhTeXoI0r9xPN8dYToETAd1JYYT3lLbIor4C6bZwd23QXYm3nhcD1lWaseODWBPW
pumQhYNEUJ7x8J9LimiFj2+3admPWPNyu97xn+DEiTUnstjFRG3I+u1kM1AgT7sM1M4W8aZYK3Zh
QZcsDJBI1IdWTdHcZrmjT/c8rScNPJKfbkwcW4EESzNCIMv5HoDSpleU84NwG1LgMQnzmnrsFRQi
FIrxzvWfIWVGg3nVmZwC5tWG6X6VenC7ln7qUzgLnvh6pshtSoRSu0QMhZKyVWGMwtlao03z7bFq
bLliq+7ibTJsT+TDrYPzNxsvWcsWxI26WyWCTXLJY6f0IZRFp+zAEhFZklvD6J3D6jMcVmLVrtp4
COyKRzm7OvXWum8fkw63VMiz2dhsfbDYh6KRa6YihlRiaUObCtlOu3LksZHJsZwSIhnVdX76Ymnx
kznputYYCX8TsmyA0gagouJbgqXOiBbAqMf5fzsdJrm3mPu7tZFXmDGod91wIpiG6tmFdRoirnbp
OGO2KGKYtY3S8UC/CK/vvQ+nFNimbfxP4SURKWxpLUy4aAwwIRhuhBjaehkmlFGll1hH3U+wW7l7
OxVku3oLmacm+rLDjIG/oqkQgX0fSi6CNHj0e8Ea7MRp46T28C5PwHrkvbB8C9LTYX7qPVid8PPB
nrBg3wdgn+WMjIARPIr9ZXSvteCRvV+hKXZtXz6MTWjpQNa1923Pe54yyClApONihtiLklMIDw7L
Gcm0wJ4UoRYTNgw5bWH1K6SejqupWtqIPHRwAw+wJIrKYeQri96By97ory9PxyKTHNKKbVJQ0O0K
NMiBwWTOm11NUUai6a2TI6w/bVjf8KzNz6CNHa/A43ZJgjQQFJBxf5VBFq1YmADcr3gZr3pDXgup
sxdGCd4aymxBXP+W6QDohRd4rXS80NJruBgra4fbrmpQUwRrEv924hKb2CzIz2f9AjwROwbKkR/3
RqTVIg5hEeKS6RAd3AaH0EorrkyFFi1yPnDFLJVqFDS9GVBzvUy41JWe7Hghs2Zp4NJgpOif2sJ+
ZIXIfTme/ujZdo/taYa3rR4cY2U8Axu4pN0iYg0hstFyuPiDz5LxBZpH02drMfRwv9wqC93Tuqhr
YRZgDGg/W4jW0QG1n6vjjmLR/Z8Cg/ax3re09lfx7IkXiSKW6RTYCyyp5V5r/gRT2RyO+filpuz9
W6jdRcqNYruIYIUDvCRcGAMjZ9d6meQ9uXC8iEiMiSUdBuEtuYyvodzpjnDyqhh/hCO/pqrdyYXx
bwPLkCONEbJffE48r/zJabwoDMD5ynDuU6Tcw2LMWrT44JmEPBx0OTKJnHcEOZ09sg9KnZQhdHFV
1QFIREsKWl03zOypyyo1oPFCD/97o3r+rKybCz+GQF96MceV0pZYAMni3c1eDbvodPAIRm7JTRtT
vyvVbT9zi5dlYTTvQVkO6rMRni5j5BcjGl2EFYE4zgqAlPAsJfib8bDnCGwxv5NjeTn5GLPEFbqp
gChZOOnQgY534s7F5iaP/+qD1eMgnafT3ofbSha879NwK4IBu6lOPsi8yNxcsfRPxO21UHNvvgvj
GOGniCS2m/PCN0w7N+CzypM9IKrYbFozkq6NrwwaC6TGZq89vgFZXIqgz5kik6dYFDcQZPWCDfxK
i8qDHzzecBC0rGkYD7JcurigPA4xrhzt3bQDCAewIxYJb4cBGhm8HWPHl7vSdpK/WFpYyFa/wmzW
Kby8wDalyN5MYWxA/LOVn4xtWcFCI7ryE+YWcnFpFCTTOi1J50BR8ONdh6q7TleBz+qyfJUnuOQe
K9rbfm2yWGkuhgKqlKfcmMm1Sk/tqDss3wfOgAouf+TsihhrZLTURDYB9O+R6hcl47Uj86/JKL2Y
6DhYGi46vPcgB+MuRWxkWhH+jPzxBV2vfvVUTkgmUtwL8TKMRYfrFkKNueQBIq9/B2hxkjJmsgUI
apOxZHnrl22I9iohWt8ROeOe14NIbYt94Q8IcFUXQaLmMVGtTt/8myPTfqwMt5srTaK+6COcYMKp
ldLmQyQZyqN8OYn9UmO/f7usBbdEJOmNf2R9S1b6aiP8UGHLCNvEF9UCHLoWHVgrA7+Uw79MVEL2
t6kJUpiHiA+/YyDY8O5Xi2B+sERRL4e0wpcomfnLkah6cxvvjFSp6nNKgub4A0mq4cug5F7gu/n9
0uIIZGKRKCyRYIjy/42+aPvyzyT3Li/rYKl2eMfQH+0mREccvvOwNqleF+AfMUD1zEJofmV2cpuo
ufOPpYX1rJ+81+5qYxVxLMR24idwdfRj5EbzCvDHeTaze0+CyzGjZuXY3Y/oVrXRhJOuWiXorSet
PXxz+CeQ894cuTu3yVJpvC9ZfwcWqtOcQAo2ok07nSwg4pQ8KQ0Cm2GEfDwKKmufwqAWeyESN0Tw
j3M15jiqC+D9KmDSsGhcp6sLC4zrWlIfmrKouXocAu6MZX5/Ss3UAvuIFqRM3Ob1+RCHb3RTu3I3
6FOa5oh4rjdMwFpTNh3mqRwAn9vMOENXcvyxNxEPfgUJW8/douWX7x0Uf7uxnHv6t5RLL/1woyEu
yszrJcEySTpHecjFMy4xeyXjT1NuN1wkMW05Gv/pRqQfKaXj9A+IKKWkffov/5OyoXobu8JDje87
DvoNZ9REQhXF1xFwsDWrKgV7b5ybumSeOKwki1NEoBcWZZ0KBQfPlUGfnG0mbH0ocJwE31jraLwb
AQYPyKyKU/5dTE5qYNwfR09gf1kWViE72dBn+sB05IoikUeBpwQm+vHQe4PbCpzZbTqLjZB8Iq4j
N6ywXVTJ0Vl9WtyhfSngNk8ZmCOsG1N3meubb8tIMXxu16qZfSPQFRrtx+QtQit2/+PVN0SgLlG3
4/ApmGimVOy2rdeprHFlhGLKjmQM8aSJTQj0uFb4aPva7zuH57xw/FD19VWsp+g3HcEWhiVA1g2D
qASzKWYlh3kbwSCXDPq9QkLibYfYSYx2PJXsbXnP0llEvK4nvCZhUkey18TJ4MXzMXonDjMQKwQu
Xm8/V3LwwX69qKQpBe2fuGNGYB260FUFzykvTlo0VfYtR6nAq7z1wFcl681nqG0J+aBsbH9Glinl
w2ykCoG4vBvA/8mYTMPE/dUNRH3GJRyh5yalAV+hJ94orUqBzJxP1LDjN3dRT49UQp3onlQ1F1ET
iNzP109ePGgeFtHj9Jm817obpTy6o71ZO30zt7NNWByXLCaAT1O049e4zu16ElZSdrIESC2UvW02
KaJXy1P6aHXb98XET1kB8EgxT17KXAkUi4aq2EHBNijxxkL5gndYlq+4K5GoQX95hpI1Uq6QZv6f
76cgPd2r7DoREmt+WzMCXz9tJkBDN1oOWKQfcJa7j/8kdyyaPVtUZxTqHNA2utnXY3JO/n0kMp9L
5zQjSlpdJBpFuTsbZkbxTxQ8k1oQPe3z8TJIXI+A/Yr3c8iRbNzudH3IzblK9tt85Lgh5O15RGK/
ROHymb6AfmxsQ2kZrXp5HJNCcTQfw9JfgDmSX0tUM5Nu7xRvwXf1I6hcFmYbR82TgA7Z1/ait8DW
XJGgWb7NqvOxZTS5wWJ1TySYPBOviPDLmDp4jRNhVAEvLu9sZhiZrd6NLTvAe8Af99BO1Xrcc3XX
cLZnQE8C2zCxe4fUua12aEduAZ064ifGoZ2+XQZt73jc9niaxTjCUF/LAywfp8GQtu1UtuPUA4sd
FjuKp95Zb8DifOHuDq5CLfdiVVtvPYwkEW94ApzUKkWmi35jdLqqfiSkZOVYOV6ONfRgO0AOdF+8
DVjKvNx1q+HhmFDLhIni4HoVcEiT+MdM7GZXsVATQcs7Q1IjKy/CBapl8vE9X/r38rukv/4sleKL
VTXBN5EkxXmp6k284bdezxpmZE+ZqNlRj7A/+76ysb2VG8am1OglZ+80J3VuOPg30YeWlUXrlcK6
SDEVQTEZwAyQ/1fufndBDg06VPH/bEvsreq2LO4L17p06ooLCuPI7TygO6nq2bF7KtS3wMfxicdc
OkkG+wUvJjqJAfnfZ+TczKfV1TmxmzNhefmAE0+8f4VwTAwsDRvOB2owZ9rjicpm3xNikvy+luMP
X42RYnUCXY5qybIab7/YXKyJ5uPS+TUWhwnZZzDExSEKLj8j/6WgFAp25ASu8DCnuJsx+p91qTuT
Gk0fYpiZ7hU+ZeSLfcwsCjNnqffMYsao0+q9CSMaV4H/o6muGi92OHn5tdAP5jUXtdrhTXsS+hHx
jvJH69fmepikHc/W4f0/0DbzLf0JYf+KRrbbHTm3U4SkVuVb4rc4t2jupeiN8Z2/FrZWV+MFK5s6
SNOBiVWsLedeE34hlMGcln2I6uArwqs1qO76BYphKmIZan2U71NoAFeTebUsg72mvZHkiOpFLadS
OM9rA0C9tHQcKOBTrUtXFJmC1VxDi4NeJBjcb/u10ZWwYuKNUc5bk3b3mCyzEccooH2BROiKXhXj
qMICY8cgigekILQrYR4A7SORzjtV56Td/rdMRZO84p2/L9Oa8Sc1IJKes1jiOUYx3zpFV4g8RgXM
UeE1V9AmpOTEkqaC1K1ZaywsKlhOEo9DcfalV7r+wN/74O6cPZfj3ZC0RVdXMwfRrXOiyHk9t+y9
N3mhr4GgHfbAudAvReOsEk12tM4K0/mDCP4DAYb8okmj8uu99VAHwT9abPm03gSpje39cOrYgkY0
oJoohcmqjhuma3Y4aSOgrz0a/FZUkCuSg7zmLnscJle+IhXPYwx98tp8dsFrke35gSnWo7/tP/Ma
xQM4OIsIAMJ0V1/7JbUaBCvY+bvut+6MzNrIzhtmO/Ec7/j6oikcMznIFM7N70ZA1Qfyz3cquJet
L83+FG0wkGdQ/59ohewrS3iu8uhta10AfSw3l/eIKeDTcKuAdbxwVseZEwlmYWWcZ4SvGyjDbXVQ
Kaa7Fz2Nrv6D/cQcN0sFYJL7uYd6wj1L9JO+zBW7pkbtwZSf/zwudDgeBse1ZCzVGnfyKYwQBc7C
WksrlnPKhP9TmBnz4ndu/A3meMrH6QG/lmxI9Bedy/bXum06GDDdm9tqM146ugkr3vrPRF3vknQ4
UCBtDHeG5fKKerr7Wycr+9LpH+TNlz1S8Pyla5xtOWyNEgQX2lnZmAC1OyF5XFZiVMPvHHfs6I1r
FEfb5I0I5I87VUrh/wInLrFcJJJDvSm1WLoV83lWoEWie/sh0MKrflEbbsIoyegCtFWjir26AjTv
OZfFCpDke3CDstNXdjJxLxQX7iOqQwnvUjV9yXe1X5H2iC3T4aUijOtmlSoYSGUxTl2XVcdMYyHS
jLlZTw6ZRBZbmhCjO7vY4nlzEqbmwiZjUcIPjIV3pAQFijC51IzFOuiUMjeZhKZJGdtN638issMk
hs56h5HIym/Rbm0SnER2JManQoP+DW37ltoDn71MJkfKc+UK5kY4qwvOAqepUSUK2DHbda511TcB
eulK7K9lwjBsoVJkO7UBPtyneKMuQeFw9su4QN9V8rZ7vkdMpiGCTCU7jhLfg2grXnGD2ZzIUPd5
MiuQG1/ZkjqmIeOKY/g50NN4CFYYmsmN/TV+GQ5uLhInG2MD3dFKCsphD8ieqNq4zX/3BagjVJXq
51+ymepKA796gDQ9A3Y1C+fYXmJlEj2pegGfstvj92Jk9cNuOJYdYAVaBAxATazsnx7cFvfhNqln
k6LW1tHY2BM7CEZexQimI7GPv3yTZUZz0Fqq1s/HZXlToGPnuawGzN3FljNvEEgE6cjW/njGUzWE
Kk33pXjib/CUB86s8XXR1zHkUYXeVj19Vq1s8Zj04EtwITDrI8UQPa2wKj0Uc+5IZaOuLmOgVWCE
cqbTislLsepqm+tKnpag1WmkFeSVOEaHJzTcgFj4Q5P0/bB9Zylh/oLpVrClB7YjqqjJ0NjbK/a6
m59MykhvwgY3AG+9CTtCpum7QluGo70teOU68p4sJMwSH/r9umLt4Hqz65dBAiO4olA3H/oIALnl
4atr9S8PJMw30ayKGp846iYL/gRzttSU9hL7XLhJCRBXPJFVvJXAWdafbNJEqKsc4CLQgpzBb0Vo
rOSKUfI0cKL9MNwm36D2qusDbLrgc1VNTwBc1bomZnPgG67/dAhepbibqtQjVbp7LU408rZE+pvm
liVM7wJVWP/QEr0bkrUWg/UG/ZMoVLIlCnAYgogrTgH7ufxamp/MZeaR2bGKFy07+u2eJmK4B7/l
bhG7WKTEZ0b+TIW48K/T/etr434D27/5vT+kB5UOooYejf/DCCF9hLGXHjrIrYzqUx7SHrAuNrTB
07GkZe4gUYRABnRpvsYCymvhGMjdiYs08jmHSgKCnqgC48kOW3WCeYrNd/7bOrJtSU0+zgvxmIY7
xeDO7DJKPXaUG7K2kNhF4r5OdHBw1uwVFnZ0UWKV/Lruoe9VqR7I0EiJwOyoMlSffmxfxZhr7ORW
423453CF4dFQ3gYvtXF8S//Zgw1Tqql22XxScHdx27rAv6JjOapZhZCcOL3vHTZovGMuBHR5ngGp
0m49O/Od2HJT10n9SA8N3PdGz1hZbxxZCu+rvKG6xo8FcZwBXWM+C9E6/r+BKAEexgecoQqGzUd4
GA9IXrYKvOX36Dw5pjPtX1XXE5g5XtZb49OG1x3JFDRBDf17xVfH4R1vKNw96MWZDlltIwTKsU4q
zXx1H5Kd42elWFC+9tdGaBLW0ZneRCyxppZ6e89icihikE1qan2GOvN+6QF0Jb2eLdrjKIO/UQCA
SfQsWNJsOwctm5P+D+mMwZWTk4MC3EtUkaxg8ukjYpKmuGFZ/3XhJnk3Btrq+YiAYOHUpu/M4ajA
JUwFVpZpYe3J0MhlKw0DYmXCVYiQGE2HOov+W2vwp7dpR6SyQ3+Rj6lDLPD73eb2rpMgb/Rd2y7y
8jxo9xWvkAkzkw1uEk1M7PG2YeLil++hCe1N59UNSDWyvBhUmRZWM7ikbLHA5S0fwSfoJb/QD591
wE7iWi3BgitM2ZYymOf6DTJz/Xin57s7xHz4u27F6cFiyCLGDzX9pkOwJVQbghLLTdE+i6rMQ/Ce
PV0fr0+zUUbiZuIE7+9saJO0MkK237mPsvdJzQR9mxRZCrh5Pvr+7gwFigWVQza3FXxLjCnjgICx
LIpxHvybUqk7penaDKigJuJ31S816Wzp0ChNs2iwdp5QZ6f5CgN97zMNWh998f7Ceu6IJpywP9HR
vjU9VjKKcUPHWLL+R9yKYxwIbjcpoCxbC3sIn8GuNVrq3/m1/uhfZfD9Vy4u4qAPqGsp+QlNR8D9
VH6y4+w4x/xruLQlsQa8v1RjmEHp+r49drkSLn//8KerjV3o6DxAr9FOWlvVGmChLQHCSHtiokeP
oBxXDtn7fpMMT3BbhtX+JEAG6Q/Kb/jj15AIj9NtokpOxEz2vc2nyc0HjMEFgvYAgiIu358YgyNJ
fYj45ccpNs6FOLYbfJf4LzDBCsyYohiO85nnnw4pc56lIR2twQIpWefK+tgMCPJ6MFge9QYu9hKx
E6zT4+20YLjtAEQfMbOZsp3PuPWSaHFY+8w1OO5/wo9q7bYOCfkL1lZ/BNx8sGy91+ReT93He9XY
SlXGSdUypAbOgHbbokfWruYhMtAYkI0QvSdMT4A5ohKJBvSecpEQ+pc44tbgIWWXVHCT9FFqlTp/
Qgs2pY2doP69SipDbdFf89h9Ny1b7kxCwgbSXZ9St84v+jkU31W3nrQHD7TdJ9lvkvm01mZkTbYo
NH1OramPG4Am1nf2jtNDq2YRGeDbc/aBn2HvsR9ysZ2szbdF7Geo+3ifgjOl7Dgeas7/goHil2RS
F/uBXpjaNBw9LBFx0mnQP8K4UI729gBG/pN31nL5S/TaTmxP+skA8rtfxTEYV+S6dnbUVh5WbD4e
uR8qBYPb0ZgOrQ+s6jZDKFejKZ0vjFaefAdbTJZkELIEKRx+2GGyQWBVXYpnBopesg46akiDVsmx
H9aJdCPnYBoiNL9noU/N3LVJIcLbnH/G9ySjNE+2F3tMzgQqJH9RXQl6MCgh9RHTn9JZoARmNkQb
5gxMne7MVp7MszLhDmNbqrBTJogBCPbB57ICmDWZ5UgB72c5ABO1SCzZlouGA/x2haN3KykRokGm
lCBzxIDZO4hztudhI1yIvRKt0A9b87s3f023qVuRMd0SUgZ257/V3FJpcdMGujHV5N+vpzD+rUOT
Ah5gkGUcoguxogV1dxzh+5g/hR+EZPnQItVKHFQMRXbJKouizMn0SphfDwRewc+HMN1rdQPudlVN
wRNWL8cxt7O4jJGCM3YtpNt6Bbi2M2jFescnJH1rKeLGEB0Y8SG+F/HZ7xcZa47HQ+OY/vgTmCiE
5VtkP3Qsm5cPRuhTW2yqMoixO/3dD6EC1/brke6gsJO56AW4hVgGIOGUH3ZXs3jM6IGwSgv02o4z
46bs1ITJD3kVwY/fm5rNRFjdQ+8oM8sxuv69TKHsejAGGTU1XVGWhmODKu9RuAdmGxSp6EOQrrkU
144xAj8wxvsoKlv+OKsYJww8Nf7joE8AizUAagOWUgzHrtTrjfga07Remtp3Oh9J5DWCmPrpTChl
to74dkpslLT4tEUkkVLq8GycjXnGJd7CEDZQcSj6nFQcZdzu56LxJNw9ALMaq6PnvKG09QNUP2NP
YIRWsKB1/86JIIEoFHSKNckMFqo/VMs2ESQ6hanw7j2kTU23txhKQoEck5uzw7s0YSKrcMgFunWK
GE4yWZ8zxBTBeBgvcVa+z0/yoqMPM/A1VDMP8dtQoS3FX7fd2q5snJzQDuEyyfRcRODbpHVK7xP3
tynV/v6A7VO1uyK6uLYtgxPAMhcv5ws3jeOxr5iaD7XGT6NQms+7tBFte7v1v4OFPrMXA2RqIWsh
84Yf6w+vcFhYxntbXUQE5/NNfHOuOFhUwRmtDETJh85VXkLTy8KQF7utwXtOuicdu2lRqMwCBVSQ
5TXsSlJwDsQ010l23ot0TmRuerR9YtTGn00WctnDW6i0P2THIcTzmdtO2FMRp+Y68PYeiPhmHje9
M/cWKOxM3AwZSddgpWqWBfTubZZ6G8VjLV9XKn1P/kU0YNV07ub/sRJLW3Ms3/VqJ3jwGqkewOET
J5JWeUJ3ttF1PzHTGOHxonQ4SQQHL3k6kzxnegFjH06r9F7xeLQCvGCAAseWmlS9e5nPYIVG3Xye
s6TxzAOqQTLun+40t+W/J7Ll2k9IJ2gt0YG7flaRHl6IcJWCr8Vj4Bo09+mdLlBN0SkzfczYqKh/
+y1bQo9gjey2RgNvR1TJ+DeThZJw6TajA/ExQepgsr3lVvnQ8m0nydNa5H/TXDnNknalczjmartR
S0WbVKuDh0MR4iybDR8QW9VTfQj77UP9MMK1KmXpV/5482i2Bek5Eha/bLIFeM7yNaOObAbcbrS0
mqsy6i1+mVuIUgHbpCVVMBplJ2nnEUK6GdvET0QYzVZxY4zbWClxXmQ9WI7ldbyCyhIll9hdiEDb
Ks/A+h75FFzX7uIGH0iBbfaKPSpioTU2B+Q6U/o4BJJhQpcWBlxjQajCubdkhiR7Cu++IUTiZvPk
/IcY5h8fa6SFHK/UF5gBlBD+OV0/I1lqxgw1olcbc9v+e9UpXrwULHiV/0Z6q/Vx8LY5+zvPUHIp
H5akcGA+qTX1j+VUK+RpkYs8PN57nopYI8frZjenNgUviC9ssbeT3MpRJfMUbXZX7W9BVQW8BSDw
Wv2P10+BiYMrB55HbjeoWrg1MCLvu0+RfGMeSPDlTVJCpcPg6D1y+gOMZ/ooEaQjsV7lcX8bXspe
zUsIpLj7rYOKy3bdg1XnuD/YhuYXrSfV+A8NBv7Q/pyoH1bNJpkJ2fVMfgzbdMoU04LvtfEexaOQ
Ry1aUY2zA2o2g9N6fWjnE0fZBj7PZHWPWQVHNcsfGozcXm9BXg+tHQ+YjKJoaRmGYxO88q5Vl660
jkXRC7H47XwMwPtk1G5CJYgKpBmWHE8d2j3ubUABqJy2WXgL6QtpC66dbg1ONmI5OFAXh3N0/rQb
OCWcIAasiDc0yoJePv6woyNzZRioxXtHtjdGt1DQODIuN/D3uC6EngOuSrNGVmM7Sjt/Q0BH9hqO
9OjFInR4hU3qmiQZDRCq6DYPbfdT0mqAbtjeEcwfmcvKn8G0BKk5+2+PMlzcPxCfJLQlBL7uQP+E
rFhU4iKb1mfadyMUX22Pu/G52/0dDJzq6pYyZ4ZGNI38j18gVX/yR390KA/BrPtiin+/VB5veMLs
r6KQHvCxnXEHGRk33a7vmg3GbtjX7FYCZK8H/TID6A7laioS3HFIGaqhBxb2oIaT/CXIkPth3IJJ
NH0GkmRZP3t0KmzLEhnzcONQ1yV2tpjmcI2L7RyYJBlej8gynOvmgFVfCqHlGlWnMKYpb5Fwhqr4
/lfLDStLyUjmRR4zq4ZdsEyFIz93OkWcLzKph8ZZQEsLfIlogu6FgrRhr8PSocZmzLBB5XpNC8Qv
E1H2WV+kbz0ux4OrsF139JsdJqqZY0t6SA0GJUMF1rlqdvkoWBYzRF28uuhjQpprrdqJHnypPx6d
ZlrbxUaO8BQawfa6AW2h1xzPZs5DjzR16zrVY3J4FyXcpDXA8BGlFMEd19xlIptsASNBNPa8YSS7
3WJZfGrksoPABNASWUP3lK9XomUE7//zyk5+mTxhYxt3v83M4KshEp1ajOHM+xYTK6QqcmP7Z35x
XNGjs5I09BjqJswrHzQPTnfaneKuvM0RE8kw5zpNUr4c/vlW9rHH2usHHyFeMtxH4MhjK586WBcE
mFgdZbLz/Ao46NPu9EmulSxd+Gd3WTWKd/vmd6tC0sMRF9ClfUD4D55etGvZhdT95Zz5KF194LJI
CWcZPwlS6mB84mejKr3QZwxZfieHSyKuM3jbh0hsI07jcujuy8O1EwIxRFzzYTYzmDOP+VAggfVz
OMDYk3sMG8sSvPr+Hgc9hSzqnpMLFGdFvhfBfyym/1oRpsB0hN+XgDo3EdJwDRBnNqwE3F+TK8QI
cZNM14qIS6JPeyRqsDhOwKPJ9VovBe/YKOQSbpyh0oXRKda9X18kYQUTT2/wThgMv8SqjrD+dL1Q
NaKqxbFRezzTS9RCkc+elBNANVI+ExrW/rdoN6iFweSzeAsa28tJYfGmF3cF6IaFrlEIzzUmrml/
l6wf11P9j8Zc5KcjLQX1uxTQX7LPGHmMnd40M3x+PBbIJDrfBv/Qai7IYzyJtk1uKEfB3UXkzXtZ
NvNy7v+wccIFelVbSO531W3Cx6K6juwpWPK3J4GSXgCx52t+t/wuwqZh0qww6moS2pJlLFvhlm12
O9XvbdGph/k/dqgs/WVMpE9NOdIQjRmWBBuy0LiKGcpSnxeDJlvZj5eX7UkiLU1DW78KtCOr3VQv
8PX7uGvcxcLZkfcF/PbxW8BWm92kX8ZGtfNa4TwmXBApq24WwWyhYEFmOq4uu2SAXR+Rd5BFYCKe
GMH7j0zFqoFcZdb5iuvmLYs3F+ZP8nPrbvcKOGRvAs5rY2ROGnc/FtWhdr+iQgmD9x6MXL1FixLN
JgMuYe75yj0CNJ4cDWVBZlSDiL8Q3LSjLGP19+ltmR8hgQh6hg+Mt41cxdOBFLGa7lNSltXEI/J7
Og0tYcOw9RDAtaaG1kWDmOawu4mNk7H+chpdBr3C41pY02SAArqC9VF8mPp2G/WCzqNOWx0BbTaV
dj35nkGdBx7A4nnjTZArV9X9Cr4QXWdZXjuRpYwZGUtJTibTAsbPqiG4wmK3WV5A1pPlcu+k5IfH
V28L4Pp1nJTdnTiUqQmcZBaKECfsYFJI2xnQVGrh3+9S3iM5eYFDp6MNE7zO0TswhuJydeOCMZL1
Uah1K0WflDHXBh/3RFUaYMFUwfPPjhU1il3PpLip9tNpjk5aFQNT+j5MdT032qfcGwqj7PjlSQFZ
4bX5rz1VmHcXZ1AK3GXtG4OvMuPGiIXMQlwU6baK0p8+6yqiJxtt93IfJ1TFHqXM4uSBtcW6erPV
az+zpx9Z1tH+2g/INNO4jfRRgTe0wUmwEsQqh16W42Ec8uaqzGRfse+LLDq7NuIyea0fwr//pRQz
vCLMEXM2ej9PI+Y94S9IHLRw4TVQuRMzgIgrqFjkDVViezT7zlJgQQFCFX353pWK0fRiuryINqPr
cJOw3sgIM5DkfwNa/imdZqO3FGw88OQRa/5Rnysk9cIheZ06CB8qrQh2FenEypIVR6P5d5OUanTq
T1+KtxVuMqrfkYOlAJDchhfTG9/5zDkJ8WPF2W02SNJeqic4i58Mw3Rp7L3lVWSNp38fuglNaSNt
lxjIqG7Mzq6s9vwCXpd9sBDPmMfqQc/0cNXkt5JzTKJhnSZ6hEKM8vrhmTSzAxEQbQwq+mJ5xc+O
dDCdcNhfVrySv1DwnSkhGP6IpYHbdR4PMnkgC1TvfKSEltplgzeFR4X1JOXJMpfiBC3vOB14DyOs
s1Dz/FWlYFyrynfA0II6BKfjvPsB8eyxocZONyiba2wrT11CqRBiRTU6dx2hRfJLPWwm+HbVfsMU
x6rp19KmkJ0cMWJH4RHWKdQN0aW12BmNBT/vWlwk9jCKGICrZeF7s2YWP5x82Jn401YnV/kFr8FH
24r0qOjWIySFeoGTzDvEeIZTy8NvHu/ojIQJRvawMtQBud2x8UNIX3WRjKMFNdeKrA2kYW2AtxDb
qA8WVTaO+Dd9t7aqZ1kmwhjNMDzFFJ75iGIaXR3afLmmCwtRlU2jkZdzN6C8G381BHnXeWPniy9+
kODaen3x2etCH6rQT6RsJrJD2DaMZbE8xxwILxLON2CRlHmnbnvUgc8NCC7VkEYaBsGs/fiDKLAB
pSAbTdtVN7c/QKC8q7AqFZkwSNcLb+va6Wnm53gJHIvlSbRmJncTr7b5n/UKPqmUkSDWKRE809MD
1xviFvOcIxRy3xp0QkS9BnRNioPHmfnpujk+hfX/Rylbm49BWaQTgjyao95jT1vH5kAKqLz0sryi
HMlGKH+6gBsUID7exSF1gEFdQVUHA3HAU2g6f+yYcOroAyA79NJVjHK0Xbzmko/vBhuuXPMD2BqH
nMCJQtM+XUoK/JcxMz3CwZDSBfUQFOJ1Dd+jR5Upph0Tk92ucAZxLFDTmNXKmNqJfNxovoBV0ZFT
RDDRxe4yZf1HRCb1qu0+gV32LBM5ZgT/jrTR0fYOFLKD5IavTMKgdZlPGTbPv67//j/STDNx37Gu
uhMsTS7ODS4yjv1dxhGVNSGE19rT1Ef0JgJvDsCmlAqX2YTIXRXfTZH8F61HZ2sP4ptjOLBQDLcW
Q/WWHB9B+JcxzNwyDfzQMEEB9W/LtjNXLdTsnAvKXlFy9AoQSF49TEQZU7ZKYyzebBNA/fbihnyQ
TXzK4AlVC4OyRLUjDh7KAXvVt4qBhZOMyDXHgA0nCzPgL48XPPAjsbOrfb2aRaU5sbCCHBhI8z0k
qLUwl2YUni2R6Zs8DQBedX/Y92Om2Pq6cDICVrJeyQkkbatatMfLaUILnm5qE0BAhJvzxyA6dRP4
QzvF6Jkj35ArycPPhcVxyfRjhyPED7y9wkhJik+wbsVE6aBLFlUozZjdWrH1/mhSN4Kt2JhspWFw
v0dZByIUcc2qxwDzyTtEefQabYql/LNgmaPLR/gXo69CKltKEvMFc9X37efU2Tlr7pGHGKJpUONU
eBoLyXIhH9qV5J0YKSgcFh/Ux4hzQTTFkrXu5HO+ie9W+STUfui+uduhCP4K+QWRW8jdrC/zWKuX
CJwV8/u8WjyV6tliOI31quclIWmSvm1tXPcf2SDhLX5fe6RaAAviBtbtAuw23t7LylMr/S+lPqhM
9nvxPNEBLH8h114vkZXn2aVKPiLYSRIZTNvftmu4t+UY2n5KXO0hbS7kQvdukK1RFpaV6mE/zVlp
0/ml8BLHoVW4rVNYSDCKhDKSSJ29JIb0X3YoWBZvBdJot+N+ImPX5gi94/Malvjsz+Jg2HRRG/9D
x1knhNa/QfFntVImR4UD1Nh8/8oVqay9vkavcWAJorn7p92bUh8lUzMgzHZc/ENJNxsO73BubsNE
rK0Ar0q0tR4oRDpdAc/sn07z/libCz4SvSoamSVFidTSkWvv3HdyuepAtQHRz+u8teSuMWwZ+2jJ
VZsJiz0UN+/YBzFvQZ+J+PwU5V7f8T4q1K3ec70jzjjtQEm5CBeT2puPjTnwHOGLRNJ+UfmOzJ18
E2TghxcUuQ9lURRZ7o3qOuDPx8H0Rizwm+mLTpNcPf+AG0aJYtJVEccoCHrqY8M5LNjzvduRritC
mqsFUsAM5/3ifG/a1Ulso5hTlY7cwVFqqgO9hdwqBDD/Cs0xKqkrUPj++LbaIN0Fz5N1APTkk0aw
iql8DCS1CWowPTYecbwsMNJpUESXofo85R6Vi6LLBPXFsTPdqYRotYJFEZPjK3QSYkwEmcGaLPoz
oV0KILEuOvG7380vmL2SCABvHuj5bUcG6ccnG9Xh2jyCPJOPvjU8V/IjvvFrnrBx9FCcNZ7g7Z7n
JSATYW2acjunAwQM63ULZAu1PrtYzaHzoojKdKMYZW4+nIX3kaOh0eMSsbG4mWQNGgzuo0kHX8Uz
FhCTzHVwa6lfDGjzJFNURxAYsi68mKfv6HtW/WVpG44eN0/7CX6jSAZ+4VMyM0K/yUeNxrC114hc
uYDfk134VqJig+AGMd4EaGuaiVkRp8Azk+RRjgUwxDmanxcM4N9ekBUZr89tZIDX+NtFrfDfi9NM
0GnV/LUP56Ikl4+mCW5kzHqMQF96V6hPJJV3UH16wQ0rsdWtI/XAfAkKEZTEy7ZU0DhJCKZgAeLq
uFr5Q/tVTtzsYLWLClxFu2m5Lfvpdus5AP81j0+SxN/XVPHNIKJDaN2gZNbLT9QiLjz5NZIvCpw+
tT2YeGFYFhxnERp0WQo8bkhcUvLmfdgIBFw7nl0n6DirjeWx3dMpfXd6l7CBCHjpA5IHmIOP9sPT
x/EKL5D1lEB6GFoiMTwnDtJq7z3QliR11QdUakxhUILtiuT8Upty1pSQoz2XUkcZc1Mssv3vTxcC
7XBsBbRyGsptKl1LJJNOCPtMwH1yTWcDlhwnS8S+Aqvh4HWOqXlawKytWZ3dQSIf+39WbAep5MKG
wmRKvfIJGzS6mKir1c3fk5IegMmbgo6nzBU0VrBGLXXseq/j9wEq9ZNNv2K1g4gTTCnc/34vf3Ka
VMHU9g+ZW58+IGREWAZc3UjDpgiBurecibr/mQFE6rQxvRLcEo7dEMZLLf89KEuFNCp0CebxtEDw
/lj82+YxbmghquueKYCaI1iR+97TRjBlm7ybmrFZ5HHYgOsPmNNZ5sxdapzGluPyO7sgNuHCl0aH
BRqcr8H+Tj/V5LcKyrMxAUnUNVlZqTl6E/dP55LS3eaSZNhnLV1MxRBoOZ6upSwGOwEFRMBb5DnF
O9uUCH4GrFpA8AwVNs0fLOPoJU1ybOhm//bb6qDve7Vv6DxvGefzglAWnTzUH0w2TAOZuT6pvKbv
Nepkdz4GjrePfn1GWnBeCr4vzugguoUVHJGRdyUcP5g3J0H5qsucKF9/INqY17lmnxq1X9W3+ceS
PuIRAq/7//SCr+0d/mrcNOMiGx5Oe417sJE50wKUGOulaIUWAonJUClJ6tjIapEKHZFeRSmvFW99
0InJxMYkt0oLvy12T5eCJ+2LX/LcJPCedXJqQ2y4u7cFPSVomVBI30NAKSTp7JlDu+1Ls7RgQJZ4
taOMQyl6ASXij1mljYB9yLm4R+hvtB7ajrfedcF0Ivdnse01HXElNVP03xJARFycFH5bYqAyI7r3
jskJE7rg/LwbGcjzMbgcbS43GBzWmiljWyNHY/IcnKMpQiuvTcEdtLmrjTEIrGl5UrLeiwPs/xhV
Dsv4cnJ/tXg6zSx6Nn9KhjeY1b13C2zKuul0GqlEP8sS1n16PToi2beBKHisM2st/dZ9jpeqd0sM
/ipdTqVPZy8BUic2l5l8g5hBZqe2VO/4LBcU8VCXmU7q5AZLmFOR2d/tq2VJ6ZTX7mNmwJcSzEKF
Zml2kxRKClhwYQ+XF/rowCYPur69cXqgGIxZ96VaKZsmxlfLIXaveC7+ZKZLbqUXDm0D7KPaXVLf
FGkXKpg6oeuDaP3JmP/jLq43jG+drEfGdY1B1OYx4g5/mqU5El8RdTrgjZp7nUpwGpQklh7MW8QA
ez2/TwniZICHEMrIuZUf3dpplEkzJ+gErev8hCycjbgttNHHdVTTGcvpHPsRC/EjntDs8vKl1DLW
AeCqF00f4Vm6ITYf5nj88AJjiHAIUbl606iA1W82tMO1v33FVrQ2Lzne+KkNG6Y4+1G61sqPx24J
kUJHBhAaqZx+dO9pts4Ic2HonkdkkLeR4Ufo1l+xDNMrg3gNK5v4UcruMHmvfHCycq3iep9QC1i+
7lHAgQc+/PzNGOXnAtazYMNSrHW+s8QScCQbGOkZDAtlSQN9PQSy3PzIwbpo5pGjFH7HCiIYsvOi
8GlqeZny1BuhWLHiywDkZcAUaskBLCVd+1uUKH8KcRd+eqkEeP4Bk4ha6Sm0Zr0Eppmji+a4P6Tw
3PLJhE8P1vv/SmlpYda99ua2syfCwmvnwrXbuJV3hBA67ECqwYy8oz2LAAXlVoa5Kc3Os5EpnyeC
US0UvfHYP4JwgKxs2lX81HOHFSf4lh+1OW8OG3oJnGoN2uPXzyVgjleeOh1hkcVYkOkZkrDvCOq+
L+bNc/xWVOrFJ0QRt8DQIHJziaMJjso/FL59D1dVXJaq8FyY/7CjN3xDfnKkskZXs+wXAT2sAop7
5nDJoWUJcQETslJJH7iIEl/zcyRVoiG/8ZTmSUhAN/SjljCIB9d9/sGbnaB9BNSbceBgTT5EKNNM
1innAD1kFd0pTICkeJpv8QrxZFP2Hd40xyTt7PwSBQ0/MlMLKLoiwNUSQHoS7wPlirYXtgGCxa1e
1jUN93ESkwkNznnbxx5zzN5kaBaPzZOQ/ls09vnJLXzoCYEsOrEJmnXHWVK6aOhEsVcaMzZcCA3U
ZvKItpjclC6KP53Xf1kaID4vyjIL5+2N4Ua88qJNggt/gYt7CRPLpUS6nfG3kdpLPESoSOHbGP2J
Hz4LWWw2NTTegiKrUvDSerQesFuVrRMG1PLuHjaNEGsJ7vwCIVAe2zBciRnlQ3bF/cp/L4d7108i
9IaOwOo4CNyMriUQc46vVlWYee0a5fthTJW+Cg/KYViqWTdDZIdfrb1NhiMxJ+zjqNd5jdE0VweL
sOGbpoW9IbIZJVc+9F8xAbfrikMJkmWU45hMxq2jpn8NCu+kph+XfCP/wKmbf3vLKszSTgfLfdc+
S5rYNWTK0zKVz47xeM6RirQIylYDOyH8b37ktokUaXy1naE+woH8S7+PJ7mVFY9Jqv+l/2+OMp0p
wKCKOKefXJyPy2SCW3B61el9xjUvnztVA0fh/PCaHKPOVIVolob2qo9ZfDhBC2JJa6B1UA+es/QX
EXBXo/hPGd3uhrn7b6Ww1rGA011m4vWSHrjZ1KV/wqrbJlSJHcL2LvcaZj4+H9Q/6xrmRgnGg9SH
6uTDpgpT7B0K5KMm0H3zOKSjMhUNeGtqkzhAZM+wjC85vitArfYfAjg9UjTFzZybQhdm/ySVpkj+
2gBQz7M6eNnKDUjdEKgm3BezYzF8XY0oc6VzML7XOcPtBu4CifX8ernaw8729TpIntKSqY41PRcu
xoslu1PW+MDoNectkWXuJHvMMEDJUGAJKXtkeiYchnoRxrIi/75KXCMpVhfYeXsvQIX7lOxqgj6Q
jZN1GxqID/JXnCpHM3UI0bAnN1kFDnSiPW4sKKx+GCmNE2vScufPXEiHV1ixrAOr17mgDbUGwBlq
TrBwRym/ZaZXD/a7K3BM03Ws5kSZsz0ttmtnvjPEyI2sXzAN3lPcY674gSKqsHsmJz4bsEP+sqt/
EX8Ko+xkHuWpIiC13EZ+mruXeXcirlwqXcufF9Y4+u07Dk2JCyM8OEyBRHxg4Ru3I7zHnmByxBek
gsWP7kqCkaq+ELnSAH6BTlfTDgeijMcd+Xl3yyYZQjgq9hWGTreW2gXDk3YRfzRIic0MobhHJODo
wpIARetW2Gf2g2hb1BMXA6UVtSuH1/2azf2FZYGZ96lq9KRx3SG/7lHV7kJGdx5jrbscoEZ1SuqY
086/NeFBIL/uQdYVHubxjuEwr25z5cbQH95xgtxnSEmKqmbbvYQoiBuEmp7598UC8PfPEMSNs4TY
P0kkHgVVVpBgTHGC8PdzA4I4SPCWV487C1iNZo0kMWT0004B5Ihe8HBOGr/3WbegZBqyFUPG63KI
OpnUE0iqNYcQtkjDFUtApRA2GnvwvO6vds+V70StMIDf704ArWB/FEUM7CT7eYT8U3MDg5q+NX7v
4av1AoJfHgCnMDwgwZcTrZ4GVTkYuzb7YrfBq6I14zFklDKtDfXSgKi7FNgiaXy0C/gOaj4LfDFH
oQBFS5YonJswPt87K9Fc/Nn9G8EybLgJ8VUC+XxnutMgoO1te1PKkjC+u6C4sX+rOg2fFv4094hW
VUUpVsJhqRKj0G+vUDBZ+HWtVSRwrv620V9nXmxiOgk5EDApHAqminLcCVnoVYsTT0TbGryCYkLD
bsAP/5d4gMswD5R5X81DG+g6r4DA1VWcKDT1/MfwzzYdw+zrd4Dbtb2icipsa7HHrhsWEna1AAYd
COi0rCMK0JymfhCcUzTwvbG1qLQuDwr1TgVyZnO5szZKrHi9PSIvyzKoWAAadRHof1gZRRJ78hdb
Ir0h4vH4m4QQl8zt2njeAe/E+EPamo4GT7J9J2djsXoo0N+mKdUKpYsB6hNpSXnGrk4iGlcaRBO2
UUNi9IsW9bZakLutAY7u9Uia/VaBcCLoI6vWdV//XViMFCHm2zmX0SXZvEet5CH5RzphargtlKgv
FqKM6kV6+1s3TGgf9OmthN0vmVIaEnqnmo/DFIduDm6MVfFGdVNLykpb9M7wwD7L1r9OLeP4AnSb
hEvQkUinaS6NkMVMA4h1koW3e1L2i8imTMs4HYcoacaU6nJWYMBR2p1nC7q8YNCDxO6cI96Pk2Xb
9nsvb+rrpWOE5StHrwQMXrVuqVRnj/jycjzaWXV8GWfPE0otIMcSXUql0ypCzreITthWwT0R7mxJ
NKclWRdn6ZZQ+HRGWBGpdiU9HhhzfOs3B2CBeJ7dUeBnTY8WjFtNvddZCIku2q8D0T/pALFZscbS
YpG6vUGnVD0ag1Gf/Vgy5m9aajDsNal2I6hIbbG38Vg/ZKfSjsRCiDzDXBklyxVbXZaq28RPascX
cytyfQZ0+1Igtf3soJKi0OnMATYUm8Qn8pk1GXBXmrAa3CwzW2gzasya8zQ+XFjYaPzVwcBDffrE
zZafzY50RRUkneFEhE7nPWAivmu+mrmocLX4f1uZs1kBi3TuUewxQWQxytcV4OLgyRxoiUCF4U/x
fcmzrmf6GnLNyGaLMIONJzsSxLhH5gaeEfX9/z87MlvojKAfIUgJr5EDv9zAPl9NatwTOyUOmrUc
gyA1bU1qwEsg7J6Zj5MBvE80XJtUFhO4hGdREDDtqK8TJoq2R/znJ1cNRyAWGnEDXTgy5RQVzzCb
1fDHTeDqv4CM4hPHjFSP2wC6ba4Z1oAMbydQ7R7hLSdK/Va6G1MsoMDytSblnNUyC8bD/mo+z+nN
vpuc/mLa6oVyinoBejI1EZE2312wi396Spf92iMGq0cCKA4YHYu/pZKDDJlS8gJybwkXDxOhz5uf
1iGglnLfojIbqJXhwTyfLPEtvqb/95ux7UdrGGGCsfXZoc+p9Tx5E7ih6L+ye6RIJ1tZVWBNznQi
0WUmFEb6PJ6u7L9jmdLVPf7Troz061cBxvUrZN6xxWcqlpCK1rcD/aTSUkjXZWg6O4XnJRXpICwg
9G5I7S6euLeo/a2vOx6Zu2msrc0XmTtKjCyWBCIMS1WgzB/cuBlYAMrlp3wyqzSROjKHr1i2wHkB
Z8tj8lFN4SROZIXLFRhGLRbHGDbabVKiBppekNEnAXdgzVKyNtdetzRJl5z8ri4dEksNGmJyZLoB
PqAOSK7AZfVHbtwHxT9U45NApMvX7sy8BNL6XDvPgIBYiUX04FH/IHtq2D+BgniCNKf3gKVdzDv/
czmcm0lZL1Dt2UouVcFJ1tZWKMEdOmjblfKwKD/tg7Y9sn0nwja4rd4Ea9S4Pp7vqO8lrIVGZWMR
aa32ZTtaMvDolJ2ZUcOVI+xGc8ItVBudn39vqozqImXRbDWACp8w5hA87ppZgaWR81rdzBXDYpzu
geUCvFZWIE6SuMesX8GwSiyrVPUqJixaN2DgPwG62pnNsPtbJXpwbOtwLIKaqCQm3PG8fDAd0KTA
o8xejULk8UlT0N518b5pOnnzLCi7SyNz/tkYZ1TG3U1GqVk1opqGinYPr9pSKgrG9OVR4Aw5D31c
95T1+jk3PxfvBJcGms0+hOqaSOWItU77cMz1YBrEmFuslYgPq2MpdBc8Kkpu69B8l/7UaDwpEixl
xZDMEzUisuyy8dNU0V/z+Wak3MNRi6OtkTWa3OC85bu0KpgBtTWB5SFCF1Ld2ZCpMuB5Zo6Zt2bJ
HSfKS7qa5Y90i9m++34euUfNSvGMmLwENo6GgMb2O+G0ENP8+ccjY8Y6kIpV2OhLvD0ThSoa6lpb
Gbhq1LtlCzisV7BbNavoRvQI67jEQuUY11RqenWODB07a2F0RNluV/uzcs9hrYjXiHs6OSW7mXiV
NVlE3wqRobDg6XOyXORBWUjhEk1fZGLRBCWQA4pLbl37/68ozw+FrmZnieRBu1xQO7QCUkXdpllS
R42LcNOZBu/QA14/HW8uug7FrX1XimkJxx0WFxxzqLEYDPShpGIVK5oeKrDSOW9HonHMpRQUbIuJ
238DLEZnzyiljOvpZuJ/xvg/BnOQRN1Lt0r7VO6jcaw2Og5e2/n3mWBK45BV0Z4X5Y2QDBQEv8ZI
eZL7pUseAFduFYwB86x+gSy0gLJ7nWevzr8wPYcHv0fP3Prnf09bdRddB/qw3bKKDmS+AQqoBg0N
Dk2iQGstsrzKxf543gNB7P+NBK6wsTf+7hywOCpSRD1YRC69Po7zZRpnYZUY9R4KYncVqUlxYqLp
2uV6SzwxDrdGrZy7AHE4T9bsPs9BnImdjSKmcT/HqiJ0JQ+wMEKVOZRhXLIO3j6BPr2i1hWwVihR
qH14B82gmRcHvr8eQiIsmwNFeZuSHOat49S1uGTmCOx5IvIWmo1hqjyTlGKfL38zUkgN9CQKjuxr
rHLOtV7QIR3LrQTUsRTzHn/OA42OMsqvT9NUwIDbcSyiFfodUM6LIgvC9cgVUQv609ffFZeCqCj0
UFDUG6K9pwVs//FIiK00CnKcRieeszkdsDPxlVFttVN9G4JPwB8PH396XWhkbOIR4C8D4jesayum
tIbJEsWdMCdh2RokDN1QSoX6hCfq9BAm0coNN8is4X5S3F0M/kh2M8B7qKJMccsGgkPE/UVj7Q6J
erYP02DJKDKqZ+rFlkveOEZmHzZVs7/vznsePpjUy53aA4CRsGePx+hnhzY7nrvt/CTDdRplsMXy
l7kQQ5mU7TX+UlIglRfq0o+U5IdYE0tMZPt0H8ia6uNnDNCG+DZFkpa/hHytHb9bMzqalYtYk8EC
Ilu3frJhRT78KnlMBt/cIMgtMjtsutnBf7jbqC846yaz4glJQHN6iA6AiEitWr0YSEM7UH+SIgVu
9khFaBnXN9aEH9T3wDjQPCvbuJRZkUjkvM+28+Lh+N15FYZfeyOT8/t1CdKb7lVOuUV8GCvNjuvV
NDhrAUN7fyMJVFvRhy11B4Q0Gh3BFOwhLRfWt5vzvWNN5ZsYiueqyC1HStGUOWO1esWZcCxpap5U
RqO3bYBOEsJi9DhlRlOpTL4hcleHWZ160OxRf/XR+M50W++iD7+7M9CUwhoj/lqPj1K2YhmxGbkZ
28g/pGW7Jm6+gxdO10APdjhrAmmfFz8QPQYxhSJMwUSdSI1kyxZrX+Jvy7vaM5P5jR/RyDF51jAv
Yq9fwjLyA5W6oKlZalu8orplme2i0Q/VQ9Ev0CJUCcEgwMVQadAwAHgfOXiFOEtrUCKHfcOdqJ/f
vmHAmTWaN4SJSXaUuTZkxXqwK76Cc5XBPG6Q2HMOSp2AKbiGonbSmpzci5cK0lh6eppcQzb8EasR
ooDcXyAuH5pc8rnpNIiBizUU9GU1Gnu1+/l83IxuLFv5Yklt6IeLfNV34veGzm/gQexFWQtndFpH
0+HVQY6p92+fhUUMK2x2t4votWOlzTh5fjg61J7aTmzvBxFXk23VnC9XLVHOc5Su0Jfk5Vcnfw3Z
s72hlIlicIT2R8wZZAh6DmgxoRFkxegRHSNf3bel8ymjua2rieFBu55t4Zlhx5jH1+wHOXIIyaGZ
C3flFhYfmvyAur4JIIg8C+OnqM0mjhDEx5DXFPpajn4NxaGsl4qOsXJpy4ERaqmHU6quyQGHojsj
MBnyuK8NUz85cBl+q9KHR/TwUDBdEBovk39S8e4zEbEjMQMag+Ax9HyZzsICBjSr8/1F4sPEUtor
KtMFZRSoX4f6qcEM9lxOvspUR8vw0V2ZgrW/wR+GXO60GAsKd4RGMhRENGi8avq+mr8Od46YD18Q
MGYGtSlyjKGccgUplwFRgKrqNcU6r2QLY6STOQ7p9aGQetSx8ZeRNok0SNyAfVf/Eq3Pq80JlxIL
0n658i8WZPZJ3XzyCkKQYlNfPS4e2uIrDFr4PKsDrCiBc20kjARNeeNvwlIo0nvSdt5CB0pZKtob
MrtkFagAcrNIJ6Zjepjeif8iY290bTA2Vj6M1KHboXBG3uxu82LCqwFH2Ej8qD5vahIKpzE1ky8V
gr7tswWz95D4+x4V07nnItCJMpfXiycdaqzGb1ocCodSgj5mY32g2pXEEJfOgn0v15Ps1BqsKZ/1
EF84/Y1DfNN7Ha1p51fw4fPN4LpPFc2OZcZ5cM6TzwkpCyJysOJGrx47p3ryQy9IQXLyQ+I2JakI
G5Ut7uWgqEBHYojiKso1C7ZacLEKnbPmRbnXPwvV3kBxje5xAy1pWC1Othw9zTbGTo0QZ4fsnjHK
xajFj5/tnpVXLOxtde1G2gN4m2OyQ4i06dLpPInnkC5xiUnMsO+RGokid5/U+9dKrJ6qMsu62gbM
CncEVOcB1F9djdRAkWsAa3UBYfxojw4EzVY5QLvcyIQA2Y3pZ+IsVTbJfMXCYintbuZGWuQOKM6D
mTLAfsJQMvkjEE/dkHNbNUK8dFr40j7Hf14iL8w3TYQfZ570hPkQ66ZLYMnMDJpKB8/nqWSvcuC7
9O0RZ7f6saQNEiRBTeplcgfCpVg1xJoaeKu9J1bs8pdmatpYAWX/PeU/kTMzIunjlUaKB4ucsiNX
qI3G8+4VUxGJy5Vsbhxq1DfjPhpgrdeEsytRWJaiA7eNH+RhJmoAe9OYNF9JJJy5KcrLZ/xqmGRd
pI7roKA42USLze/biv5d8uFTF4zDPo/woFZuCfOtJIWbBy1C86mFeEg8ZOjxF4bHxkw/MI64wrCy
Y5zHnHnPg/EEh0nIFigNGS2ixTg4kuO8UA6yR8DT/J4Od3h+mFBkngjcQ02FI6NhgkMFgYolLwn1
hxgTOKrOEqF5bAJnFxSRXYyL58kMMb/5CFiY4hWy9AUcFxpF+aNLlAPAvQMfXKPz/+wvLYKh5mfV
oS7kOksmVMZj9pSLCiyCf1OrGyxhumXk4GMIt7hVyP5hQHEO4+L4PdHV6SPrhHbNRJ2WAlknq8hd
tzgJhmerNcDAbXq3FWk0o6p+D0cmMbAgLHkd37FU5KI8Geb39K0FTi2pIzU8fAnhE7I0udvhPsXX
WCkhp6qy9o+ZTtgHLLrc3UA96G5816rGSGTaD2z+O7oXWm+PZpwtPl9NBXfgtki+QOS6X6IWJcxN
kYpXFvXUj8xqXUB9lEgUDRxZ8ofnA5sNN9xm79Z1iX7xOP/sbdRdnUugazp7nbdMPggz3yldPntx
BewtXpzaDFGdds1FtXQzzyKAmeF1EXW0SYxcVXUhzq2db+OoRBXGGufA08Yw6SghedcRXvvhjeOl
OSDhoiYTmVDClYSehv27wfH/O2LZs6dOOLmZvBe/wqXPDmllyMfv+AjK4Pdp3VcNy4dXtgws9FNw
bC2m0RHFQPcrPiOFPoT3h51YpEaJmu7MElnXAbqBnCpZCeTHqivLx0VUbdCseqTXGf7VZ5huN9L4
pqZuRwG8FzS/AUQDYlvDTzxRccwdf7UCcA2VxYLnM+pTn1JVprDBqT+LwQ3WB/JtU++w/rilEtwt
gf2e0ezcZYSoVmz7UNx28zoIguEWAFLpAnMy2biheed4csB+OZy6WeEpG/PKv9MUtrzFtguY++3q
7S0RbIZRF1nxkY0toZy57u6zrn4DRLlkwySEDoV+LZGtxDtnJwny77PoO5P+08CP7MMzZ2pua4Ri
v9p9lFRQjlyq5apH2E73ZWmisrdfNAWQR3+Ggfcdti/GJ3oGD+qVkK/6QrGHKNqFY7oAnnAOV/zE
qWa3ov/zXz5Z3mlq+ImGjBVZIhouDcLRXueuVyz2SLXDjqu4sSgQD1G0gyz3Cf4FlHg9ocDdqodR
SPpYDV7bHQHyX7QvLXVg3DVsyy9DQ3kkPG5JAocDO/SM+oFrVhwrP01/RjnJeg41Se/HEO+L4g6z
cP2S7sORng2iIRnhnl6jlvIfOIv6CIlLgm4f+SJjRxWrjPOqf1W0CR5TdHdtoNT/9B/4XmXf4wQ0
cxxhU7HgIWWfRFKg8KGrAdoXhwf4Pz/9ktn5BaRGcSgy0kfTvSi1M2rK4Gg19+XsfTyuoAG+B3rx
zRaIPfGa2wrkkLk5IytZ0Y9HQyxBp5eNqdU8cfyN4Wtwctajarty5Os1nOW3MxvmQGhnA+HecfwG
vk6k8q2cL6SHWZsTwzwJx71DB0u0neatYLTR64rI/d/bgZEtEhZO9sWR0Wls0DxIxHeLFyd/ymAS
YB8tcz9Jdf/pzJuSv4WS9HFmAmiyppdMOuWlAwaWRzeuVfZ3FMWC9YfvPlC5zkf6wRiKH60+v9b3
OyKaB2aglP0IRxQeFroIKMCqQ2hBEsVQr21fcVTj4bXWYACMfKGqXlmPJcdHubWhtoK8awUanvvu
P8/pSmZZ6NaiGoWMb5OWP7CHLqkCqX/0gZHrwG9ahiPuBtpoB6EDDf5b8pqPCUrvgER/S8QJrQa4
wQwXxZbgxXDnJdsVawYI8+huGOI5PXROlV8Jr95wai/q6eJdG/yHCPjSK70/hVd22hhAki932tCD
/XAW4KNwOOhkHIPkTrwyi5xruWZJmm7g5ffQGlDeOyfhQdX9qJJh3UhXzWlmC9jKYvu52Q7xS/Kk
26I7wPQMYIKfs1vzCkEe7PF5ytBmElgKey69NsslA9ASd4VNJ44S18eERyFmSjgq5T+1mBP5CIBU
k85XBL0fJ/dgtecW3LX8DGcaOgVP4phyjYyiz7g03gV9WsT9BvJ0/x11poM3qrmSUmOOw/V0ylTt
nlSjpCLTvzbvidZ6rgizPNJTEd1ONvyBLA7auCIABjZrHVAwLjjr+ltq+2auynXSjB8nQRMp29DK
P8J/GcfC1Pcobo4jT/HZ5tCF1MupL8DuoODjQswqtNWMMTpWTkRoyuUhUDeqp6FE8ShbhUSJmPv7
vgavM3QThN7obmNBTLT+Rzd7zTSfe1XxzEy8Mn8B/zrshgBVdfTWvF22I3bdIHSa7cl0Tx+wLwA2
azB44O89YXzdFFdSEQa6w240Vyt9wEIyVjbbR9Xf8eN/PoRrbns//XHj9BpEuYjFHXwJef5LC5uo
NflLi5xLGwiBDYATyZCZ5DbzeJ0MHBB3u6Z8xdiduexMzvS80Njkrri83MQVgCY+GCWIG0xjMycS
XH2/Fz2OU+ZZJH1PvkBMyS6nVWRH5IozhJoaKGYmKsUj/cC69QCr4ebVwp+lM5akoArdZsOMFOZO
PFGZIVVR0HIUQmNMzCw8+NbYcwu5mXh3PUtMsHRwMKQsvPsFpd8M8XgPSxVDA5Xc2DRsQuDBsiTW
Y9dIOFg+52pB3sZH0jZFjmiC6DmcgPFerJ574vREB2sxnZDdHNmg7DCiWX1SFFdDhGrLUAWKlwlQ
YERGKJue0sLuLJQ3kqdy15cYWM7pbAFj7xp1IczMgoT+RowC2oxeoEWx03ggHYXQ0vTJE337nayk
tmdorJniohl9ghnj6mAedyEHvrQEuI9s/DKCGscYXarOcTvO/NXh0Akh0z2LLGjeedR62NjOpeMP
G3WtIiXHVuOscwt+puXgrcv3HZIRlytnlq/p6khTuq4UKeWia27t/2T2o0SI/5V3lDZli6Z0TNRt
+3FFLtNlUlurGrU17CJjnRZcgTK7fEryKJ0MS6I9GlYRiKVgrtVLXT+VEEtV/MWeddorS51NTk3w
A02z1qvQyoPOrheUn/iu+y4b0e6TJ9IGbzLJ8ae6ye5cVnQnwB0d3L4cXjIj2aCzoyHfBxHxWPSX
2NU3a4kh5NIkSIgBTAhwgjznuWm0dyH/XrLGZPV21PKr1MD8iZFUU5dJhG7pO+ba4PubQzRQlC7R
lNYVocBh2LhLkNcivBlzjwdR9wmP9KSS5H+qAzdtku9D5VOwQbJRACbb7neNOFErvn0lHp/vfrkE
+gKqD1C33KKXwjUv9j5Y5P9WOj1mXsCbhCOA/61NjTNbZOIC4I1MwavrO/iR4rRrCCojzX4LOxgI
TylI5/28hVlIG3M9cXJVHm7sae7p/pponJ1UbGkdwBncTHwLN+LBGOLiSxRoX2yeokRwFCEO5TS4
KHwtWnXsYXxgzSx9cBgsBrrQZ/W8EuHgm5zvqnxKmhgZsIFMjsdlwRRQp6ngKrscvw+XUB5S7j2f
F2k+jBZrZASj4+aTiT8K3eQXpdE09Cj1r+ObPznaJoppyMMIa1ZNUY7zITKZL7lZUn4RN4titfIf
plxvL88R4662jRX9uUKNNng0Qm8YnfdsAJKjbCMRuHsQKIPiEDhgj9CJGARs/8gC7wGktJk2r2p4
g32bkis8hYm7IANYGmJBEEzVyNv0Z2pX+NutAMDoZBUj3DpVwOx6SxA04r0R4aOTjmIB8CUR+H8S
fPK0PfsWrEEUwTOjax3rfUa3lCpevKv56l50cw32vVtE+MD8dWA23YqOlopdiyGloPyyqADMYCDL
snutTVDiQjWWyzam8D0ANf85Gj4cTyiUq0MCZ+J96Xgd1gsNcKtOdC4VSucW8xVGM21KIJ2F5Tnb
6LFCpSF8ph28pK269j2muUn0HYZiXg1eLfW2jv54GABjShfeRWzeJzvF2d4sz5PQzVPh6+oNTOqO
cc74qE7Hlt4P5mCWmYjodA4MwJ3SLlQr3aaWwGhffNicJQrR7oy1vz3uaLdFDOoIoHhZBcrmLujj
5WvFbZ5FI6D/IiUQt1zignVUlM4QGqh0SFE953WQ4Tn+f4htkg5X5J0Pk+XG49mzPbN4AxnqmbS6
c0jw0N/g3mdPMZ0bRKZ6s6xiZn9IM9HQP+o1GOI9nINPOdhdYaIxxcin2tu0lD1hRhh50p6YqctE
8PCaUiei4tYGRdxTbZPdxOt44iZQfahkkM7lbzbwhkbp3V4XiqzqAH6MySbHNYyFrDnsdC8d8FlM
T+XcgP0K4WC0KDfGujwGhHylxqkiZsgeQDt1CmdhVvWlG+Vy5/O2zErWcIbPBc/rnfhM1cVLijFp
DBxhLXxSnlNg9uGxsMXifdIHOgEydqSQNCSmFSXev74mJqqqIhnXWl/0UW7YmylEjFLWIjgB9smH
juOoMgZhD+tywpCubTRA5Cfyve93lCgAtiLzNAEDqzK26ogCciQl3r3ZwjJdb2wseRApTVOBp+wW
xsIcG3WIXW4Alv3yLlJzGnEySYXd7WhZaPWgUuzRyzu4EialxEv2gdjZ6qLlm3ARYu4EUX0FN5fR
gUgjpyJd308e9Um9+/0DgdUGAWBMP9q+/6/+v11EBGXila+99UkST9wfOSHdoSMDBLPNm1SBG7i9
2KP59pR5ZyNy40NvV75FuWjI4uU6nsQfwn3/1E1fw1A/dGqPaiElVB2MW9xA6cBSIUDLsoscQW0X
8UoK+ffP11R4lpGx0tfRsetfhEJpANIoayz+yCvWPCNmHa3w4ma9fsBiGOi3Tkt7ku1fnhMOEtEL
btvdoOd3xgT3FEZgcy6HwRwP03a1qjWetp/BhSFNewgndi52ceTNfxfZTyH14iRl1dBxz0UQdnXZ
Hv09xvn3hnE5qxMQBdWnmNtoU7gRbmxSmnSpiqMzRhPavPn8B1iIe4VoVMH/w8T/JmAxklEyWcOL
lHZFge1UkEhHWm/JyDamCIWZhj1a4i0O9+rt6BOUqwchQjDbUXSaHO7oC15ZOgI7ysM83grKD6mR
hem4u+LVr4TqXVFEvT/Warhdarj52ruUyenZGrvEiNcMd/nmQpsbNEC+q08HBzR78FD4uW3vPpt9
nteGevhkupo+VpBWy13ZNlnH+q5gntTVbg7F+l5eKLjbW54HNnOhOo+oRe+w6MZc5tn3Apk2PL7k
oysyM5nTZWyqCz3tzW5vG5erV999GqfWKhuXxnn2s4S4qRg8HYIVVRjqSjOD5xCUCJJTk95kmgX8
RMxy0ltivTWPYH/lTLGj+lLhRPOL8E02YceTR0IR2/wyd8WYYLDz00dtuTGufhtdtZQFWTn/4f+H
s90YkCYBaZRXOk2dx6ObK8seqey4UnyzbqV0pYI3AxXFd06qi3r/CyjY3GBiz+NtN+0GLbjbhbqX
iVcfPtFeZfr2XQ3UCtwOx8UlFn7lSpQVS1IuRr06QNiRVuw4FZChe6ZT5Yr8euWD+Nrq5vgE43++
yW+7WsiYrwZjm3Okx0mqU+ViMIzxiGvDS2dsp+RVhNnaxMp2Lmyb+iJX48ylcx1BKYWtljF79oXd
xK1fnlIuLpVjQ+t3SekjfceJ0OsT69RB3mHP3Dha+r8GEMegH1a4AIDWongP/54He/LhIk0QfYcH
LVqPmAaymfwt3R/YLHcwpzCgG6ULE+dTjtAewd8PDHXr5raUERPSQgdeEd/3GaQu0PZR/AaNxSqz
eb09X8mlpsfx6xeBg1Z/ml2TcNpRlfeKyxjlISE4FSDrep+SSnnrv5XqTQEs5Ys1idpGGOKP57Bx
RrhQJrCuPSV3SnkL0m7gUWLSIb2lH0RRUi50/r7l3BfmFweQ1H1tDuKj7LTxjIfnaKsbi6yJvwnD
hQBWSGVwgXWksmDtYhDiwusZKv9hW0k4wZ/I/0IOGHKsaU5OBVIDf2kFb5yyDD+d/61gualHDriI
0qpO5YIbenTyEqZ9I5TulVL3zMhPR6n1xvo9/Nefbi6EAcgW5SPKrZYHbmAzoQrZuG5DeBw5bAYp
lLsmtpOXOOUH4a6OLbiQUN8OivFrevKndDsC0BtY/82FW0YzwOA9ngPIEL+gPjSP5xtYwHRtd3cW
6MVizGzCO3WkXlag+C0Tv011lA8T55cUE4EIvVYOShYV/LRtQM7Dm+X1JNTmkrcqH0F8qjOIg53U
k0x52GZkszbiX1ftuupH+WQGoDe7EW8CP1JB9Fnujp/PRu/sQ/nKViWSm8wpvAilaX0Xjn6DVXeL
63tF+aNwgTebLzeLXjtaoLapprRBBrdP89TMcCQ28gNM8+wI22fMXX7u52TocDIeyaHR15tEGWYp
UOhgrXe5jDM0mlO3CQDiW2vSKrv0Pk/ToD1cBIxBKtzhHI7W3/3yxOWy2jCKjnaTEFev5RuKRNMx
oqjzaotjtov0RPz4/2BGV+yG8DtNVDTaT36ZgO2OJo4aJSYPGCDCIgMt1WqO6LhhOylbNDFpwPoJ
JxfGsJNZDKFjE98FPF5ERzBdlpiKuTLD/aUGMDDnc2+GTFA2G+Nm+jm4ZZ4rDsRKeU7nU9CiPTrB
O/P0OlvZHQo9c736NCjlnP/VdlJGNAy/XC1i3ypJ8McwowCbFgr+N9TR5TchL5G4yawx3RE8e48f
X03Yi64b2KnlpJ5cctGIdVBlAeTnA01Vfx5vxy01cuhAgsR39Lg2CQqxXGOoMcNU6q6+qsdMlWB4
TSku8hof5Nkj9V+uKVHAHM8oOTiAiVyYcvzrxFMuuVluxJGNGzTG7QIYmLdHETv2s94TXV9t5hg/
Dl0uJN9hzDN0OhCpXYf3Y4MMyfJqGFM2bDKmxRjw+xI6GF7Wu+J9sPkvFLrQ2cGQD+jIcy2V77U+
mJphHxsYfJn2wAKNyHP2xP0gCnIejRbDvFcrxAoDzAH2cpj2j0VEyG0uPyPT6mxgA3qJGFNgWCTl
V89QhPibf2dIqj38RDrf0N2vn1DVVSjyvcys1H7DiAL+p/oak6jcJZQDSxPsKbuiP+l+yCsIoPqG
ee93jHsTXVa7knt8YJFfOPzh2drbpPPZPZJwN8EiSTsdQLM29F6iR9C5s+3073UylS65znxDOumy
DBHShkDdkuPDdQfk1QY8EMYJdQljVwSAXbpnZBJCiA6kpdLSTxjk3YTpYs3xEWbR6s5CDEjuIWCk
o1vrDSsgQo16bwrlq4qFjpfuFWvRVkk9Cw7n2JE2/F/7PvtsywB5w9V0xJxov0BSmqvEfWz9rbnX
wt45umKumUN4sEyud8Obqj7MOTcdF8MbClp4ZvtQ3w8cNMA+bXo40Elj1TNDT8Z4ps9+03ksFPeZ
jaV0Bs6Ed440yZQvuU+wJhaLHZ2TrRmh3OTct7uwQGmHzuP7EPVDyTGIjETpz1mcawwsx1QeM9N6
59LMAXISNd3wogIAZWFmOT4bF6+M5CtKgQ14Mmmx4NIAdSVnZIt4dzUHHhI9NmdjqOaQYHhi/qTR
DuzhUVcXVDHJuVs2v30JUJKh29ZzC/AlWBT8yFPzCVP8UgG7EF5592ERKh6IJ9F7lM8fPEITTZgg
yIQOvgwczWaLTGpcyHs3itnKefhORIsZKfVQfZQ4mllHzjdGDPNp9R1vpifTbF9JXPs7oFvqdON7
nlwVy7hHYKjm7aFoRuKgscH3RFewQ3tht+DqWEyDL/Iop8SNuCrMcB9Pz0gHTTqwewm8yud5LH11
9Dpx9LqYSsdAV6mlB+sHQlT9PydI1K3/QiX5mNw0YDt8gQ66wh87ojTRChbuOAGrg+BHhhiycFE/
vXQeSTuNOb4BXg598tUgp48Mywuh2KcfHIAmoIRPNS2cc5ukpdGrRjAqKfVIS35Jamxp3YXyDzsA
q49U4OgaX4n+ppVks43EPeZ0QAnDdudzanZv3/Sm1qYOXLOMNeQwjho5dwjDHaP5qyZEOhe1fge/
+vgVh+Htxx8Lb7Y6a6+D7LmM6Mf78uKHz51xtVCxeEBFqR+K2E85dbddUv6AXVFmoEzVejSYPL4Y
ObQuKPWo2RogbRZQaTXJx1E24+CglOwbq7AoOcaHoMLZsmFHzDfNMEtHdslvzWDKsglUdcnanRQ+
XpSkdA63ugQMbnGdYy+oBOJ83Isi+qbRPBMYEsiLOLeVT0Y9RWNeDlvSfDNCJGzP2HCNNN4ImY7G
hV8F92B/Wr4mFcyDn2cyDb5H6u9ZjlzFZGQGk0G0txqldEUtZH5Q56dGYxjf/VW50lwPOEYEyHz5
tARsi/jMcx/1caGXkcWS4iz33wAkEq80VGwfwpf+V9+aNhJYBO3YvEfy+9+0h7s1iAUbKbHIhqWz
Adac/OrKtO5kmBpHglwJhcuusxYVAW5b916tWS2z4A8U+ggzQJYnfMUhKpUmU9Juip6R5u0+xtYA
fwYl8wEa6TDERxEyBXye7d4zuW+gQ/D9UweP4uWMBu6WB5GOJBn9rWounu+R4HqZNHbqPDXvodqz
lJkZ17dlGXmE4pNu+4Ruc30hL6czKs7UmTfmDBXPfU/dBriz0XHbqVe7cnZns6uP6PnAForUDaMr
80IwniS33fbtciqht73vDKvI/6XE73BHONAcfwO2anFGemhbs8MvEuufrNnHb7MHaTEOFCtPnz2u
Z782KK3HjOIUnQkBYOMcgelDOFLUp7NR+vOxtOTBt6gb51+uT/HLr67m9eGGJA6a6x05R9FG2grK
Tw95qInQ+//b1IjlYGEEsUBHajrSPjRs3Db7ZrtGwHXVfEBAdVSwVEdejwNkTz2TMrWic01NWtOO
+WYF1u7H6Kcayuo7ymY2sjn7+vfx/V52Nt5yK5RWNLQBIZXlTtqub3AnJ2G6OkNW6YQ8INOAZls2
N6sC4zY0btAx47smLqqABaIaEowiQHSUkezJKsdNqNyQUOakEQ/bcr7ehHtNQ2UOBYM9uBgKXoa0
ekOIsyOcHc6XipteReRLapgTAeyw3Cho1QArzTvkuhecH3DiVdYLilYlWcAuWSyrlQoRJKXcdxjL
xjctQdzoNg2xLaBtB6rp6aZlTyUmyQ5JneES7KNLSgO7fmI9Ozi1ZSk1vjWgwpDEVTo4VSh+v1Vp
3oG1RvnwqeaEWPCn+UiZT0lJjRQ1TrJWeesRoXTjXi7rBP4mVT/GqmKkE8qpD8nGwHDBzeIC6Nkj
vxy7wpW0aip6lIDoCizcuLKSgQt3p/K1Ico8zWkon2buSr+aS5n0GyROjSzHL1rIBB3Tlkv2LYIx
9TWc3bpOP8OTNHDesxX5UZp+9rfG8UeX3RFwV7xO/lsWVsvgTGq6PrROMUFPTX5zm/pR5ySpUGWr
NBR0Or2ro0wZzasN1awEl/uZELGPDwqLJak9UW1yDGY03rPtdV4Ef+oV/T92Gy5SzZUgR4UxACJh
rdgvIHKqtvySuzvJlxTEwExh5Qlv9jbRLd+HX9mQLxZRm66pbGOrblMDnMkmAewy4mb/E/R55Aei
p5melqcHCvVC0R4n4MdRNamfFm1NjwMJGSTa+M0FCnpKE4cdi8stHHOoFx5TpUj2SbhUuUlY1aaC
RKVUirvp/wWWwpLQaqWLfryi1P4H6O8Eb8aBP4qVX6cGsDNNcHZLzxkFlUuYVRTvHhDYCti56ZLx
ZQ0ng1yoRT+gBGGtMBGHAU17VQnLgoEC9Yfe7Gdc+Uf/v8ybazac9usM4l3uVmLdY6XZP4IxxQHL
8I9yS4o1SKTmmvpFvFnreKRJNe/wklmFE+TPLKeAmTD0ZNvKP5zsjW1pIyvnPpSp7uRe/P/nqRqT
fvV5RE4YiG971K7CajTNS1cqTM2RRzu3oQuKCQR2ZlL3trztJM7LnSGMZCiDvklOYY+KNMTBKXZi
2EMKhkjfyinVA3G3F2UbWRvOnj+WruwBqXhseAqN19exqYLxGU7QX4VFy6Qaejr5xIP7f474ukQt
xS2ujBb30zq25Ca25u34N49pfmKvibc9EniP9jvhCps42kr8+0CuJVlv4FvGfCg92DOVFqo43v/v
m7NWGDeBaScCJBDYJ3ZzlJP5aD+LQqMyxLP54TcMZR6SC5V+MTcNzAv7AP5O6LC5zw6fXoOaWC3p
1/Ztv/0Gi8xyFYoHhNnPUcalAHk4jCu6Zs1MrBHyyes6rwjSTF6DEsgn6MKz7NrN6KQBgVfduFhq
bvZKysbtqPDA9l1NZ9Cp3OPWaDjp/0iAw0CIou8UftI7nyapkay96CUWwChyzlOX3LLMiZmdRT33
wEztZDVzH/8mxYTDpRIMhAQS0TtbiuoCgNFyxeHQ7IGZ+d9KnF16DYQWNsI8B4KCmxqVvZeO9mim
I9Q0IMjxtge/CK7LVQtFGvHbUu1VMOADd5XaPnc2LKkdHzB9cTvL5rFnuTGZrTZTaoaSyP9iM8H9
f99dB9+65wW0r8Pvlw6yzqEGKZDEMIfkejb9VD2si4DdmDUSByGZdJFY20x6HGZJuYUX0dsyae+u
aqVZwzBKl5uErs4dFxLnoXfFfzSXJEGk3zPWR1jZGQZ61wJlQECS+/A0UKir2Cb3gRQLKgCJKHCW
jYvD1CaaAk57lKqa9RWTQgNUAAdbE5WUQAu6gQiZ5v7mJSlcaEfpBMztn+8Fz7CgRtx7gmVl8opp
TeHGkQxiOs6mpCnvjx8aJ1D5nAzYVqkwE/ZvEmdqDHEAOkWfdzkTbIVsNnDYwqj7mSAW0Nej6Yo5
8dwCzjpIc2v+iaww5QFX2qVRQWniGzfhK5s0u+S87CxUqIdBNY2ONZkQSPQE44sCC1GRc4a81eBs
OqMTuDRNDPirXEXvOf9Mdy3YRo4KJMh4RtFe4lXzEAovIFxQ7qAbQtX8Mb+MCTgnKtbcpopu2r7H
s4tGo9JXyZLS2EjFi/ExFvTPuBbJkUSnZmoYX+tmAekYH7KrHCT3nV6Bv9Lqk108u9tXYdbYrcyZ
mI7Ur35Oz0341UAcYYNw+t72BGblNRKih3QDTizYO/C45ogbeuuNzXnwZIkFW+utaUzsQb1mq1Io
G97BndtamPoQ/5sTGdq+l2Xf7gLU0jaDV/CsP0iPc/J2syYcpWTh5rG4F/9lqrKwKRsNdxJKwrk9
ugXa3tb0XaCHQxVHcu14n70QEKemJ1GHuoLbnP27lGjqCfrbH36tyWgF+S7rNHzoT5D++D+HI+T1
kbLf3UQ4/2EGtLGAZCFu7JPRAIhYHII79ByizESseHU4CdCeRNaVSMUBmP715B9w9O7Q+/O/CkY/
FdOXhswT09sAZ9YY04tpRguHKVs1q42fXtrf+hVpP+zY+74xlgNQ/Ok4E8kztWQRYacXxMM01qzj
Y4+migTXTRoUKuRwjfgwVZnBlkarOyocjJsej9MMARFE4kxfIeP3GKOqDzDfz94rAa6VMEMJFb8F
y06Jn2n1DFErwx6YiejWD2To129Y8wdAW8omHASes1SWC7VtBBUSmwYDnvu0LN8EcDwkv7SLcCSp
aWooCDcr/kwL7qG0I39+9LymBPasHEeJ1BugK2AvUeOYZZcJkHZwYZg2Goam3/ATs8fYPjkHuD3J
PQzERa+AkyNdywUHu9jKsvhJan4mBWEfTI9AAGTNSzfy/XMrMXaYox0VZvvU7vTH5YTX1sQ60bvt
OBcK2LmNpnCzuAbN6P2R3MerhUxK+A7Dfvhz4vR3yNGU/On6Hn03JzI1vMKbmtmxkjNed7eancsK
2yVGFTFKSjIioILKAjIqXwB7/QLdEJnsVo1HGBvTDsebozsQos1D6NeUL1YiHq50tWrYGgWy75rs
7SBNvPicu7lCapE7pIrs+PVUZ1/asxTqg9MUeGliySp/lQOzoRpugLdWT+DPXwg/wxvHsZ7eLBHJ
eBmu2Vs8umr0dI//ByYzXm1mzmX74ctv+bZ1oMjU3aajL9mk8YzXCqKpxWU3symuV8iR+O4kXnKM
syOeILyJeh8YTZlKTv7dTOqR+AESMKdNSA0bQDAcMEuI182vrkcZ3EDfMSBieGEJ1hX1fmXWKkNn
u9fb7+N0KcD6e2Lcs0t+oLvTTgFc52CKwpYmyEekLMoBfgH7OqRL1a+tpQgUrtMZGsITwa5Dl8HR
NqujARgwkTpgTZL7RENxixN3HbRSzHfW4U3kyXE9ZZOmcaT96FTHeXoPSM+Gl6o0qp89Dv00JDHW
nkkcyXSnD9zUR5B6tNAvUWPfqt9Thceb4O4Kr3wGOP7nrR6bYzqv6lkWcyuCBU5BlzRwXfaaAMeJ
1bYVLgNyoJJGx1ixriZAZI8KO/pSCKQ5ELBQhpATy6zl6c4G0sdXG3NCp+OAQD6gxREH/iUjXfuN
rUjDWqOcZlUS6WDvJjtk9PVPDwDTSB1AQ9H1FRiizkyTtT8ZIY1yFtGs5hUTrBr4On3Jbb75+pB8
mghc32NZBdRU4P+8OHN49kK6fy0/OMoPC8PDw+TLLF5Bl1+T3/NeJxtlxFTejZPXpR+ogwUbLqZ5
yRJE2RuEzhDaEAhpYmncDTxhQbLmNK82SdBKh5pdrhdTRky74zPx25lY/Xy1dGo0mp1/tbEujRWD
xs49VG1RUjoRyTKniYNTB3QEd7B1EnsAg77HSVwt7oR9oEf78Dcg9x+BEI2KArJZvTEsMqJfWDeW
x11lci0pI6WGOA43cPlngdo3nS2xcergxjkreHi/col5PPEaNj30YtswYfHpViwMb2nr00FjRYK/
TRpnoCuau/fmnENHkGAiddsfh3l68iI/EUWpI8oVc2jVn6rtrmRaKSGtXpPPZZG8d3cayUEne7Tz
zdG4eLYKZQ7IH7xDiOJx7CoKxEYY1lFE6VYo4ZDVKTGC3rhloaP/tHfAK5HfahFTAwgtuTalW5QU
dkAwot2c9wFl6Y3LfV8CKcS3J2JARRdLaBOZguegRQFz05J6VQhPY0UwRH0juH0zJzxo7c8FGYNM
8MhNn6w1p/Odv3EyCjIkQqMLzOQaNSB6ZOpiKNWt3yTZ9SBytXxMcPR6ZlPHj+aFp2SStm+wIuax
TyAYlxUdLCEZ9LqZGxkdOwUsvVOIzK9ejkOjQ7nwMASTCwnsJcmZGs0xKuUf49XCK8RbKRrNn+Ap
tTsw5kya1uCbgnW1Lm3qoeCbvzqO10LobDWwBFjYQ/8djohaOQ9qDBxBbM4r8cvE9QCuOeMiWS67
kXpHQRa0XqfEeD7bm6OJ5+QS6ZvI6j1trO90N0+rreRlUg8foBm5FOpN1g38gOFxFTZbLYXObkLV
4nNx4JbtjNkTfHRYqpYZZdk84WZm6LuG+k9Ljmm+ExlSwm1h/wKUqrDTa/M2iLFF2+RrK/HD1F/B
0tVbz0Z5imRk7GkZT33oWoRdUNj77MaiAgV1FwTGn1were4lMMeYZBJX1lcHMoU+aDasELfJXMv6
mmIronuzPzpKgvMHGvYDSkhODzJZyoSoWhOCvBNZSPlbyQfdbPVIPpzUtkazd8psYXknw/PxP3bh
lPOIEl76CgUFC9tA+CCmbmvojU5K6DndaJxWFo4DU4/XTXmW55/F0dQ6/2A1YswRNURWh83H5tKT
Vd1UfCFPwyWN4MkZF++mDJxc2fdgBLmctgvDAzTwhPbxf2zsh8mLPGiWY4gIKS4bLEITv2xcAGF+
RVuODOOg4ObzBDojo/1rvuCwKFX/ocBNnZxCnRx3w1M482XljczNFEptIzQCjLLBbLZtYbLYjGHz
IWT9aAZAT4LcScraPYy1zv9o6uWOAOgjZzf8Y6DBFKkHjngHiGTS63MGzlGz+q15MHI5LzfV20zV
yzkMR5Lcz/SzLYB9sBDZ0u+0H+MxZwy6aUKU9JnLXQgNs96rjlWJhmDxy4BAYRfI+SoK2tFBHbni
QOa3ugtKYfROLuZQlSh2/9yqt/vuTWsNWv1dFO0TMxWh5L30nc74rQ71htr7DuzqBdLhuE4oU+I3
vD7dn4iEN9U//BZDgilNFwuewUkmivhql/J1wlT6PC9J+aC78v0OxhzbXoXjzyRByNajtx7WsNXN
UmiUhWxfpQ23WMuBfeOdQE5c7Y4RYtr+OvuIX0aajwm2QKy8shp6hjFmWmurTkVQeddwkQ2EPqyx
ok47THKUiceozJ8qawUZjdWemKIOnBe+nMz7E3W1TYOHEX+mH9je6/mxt0HMBGjTCrWecvVsjxne
LaqBwQuSCk8NZArixj7jX4HnfTQ2SSvl77NG8tYP5LQdpwQUf2BghhTyRFcakL2vPGlkPnvX5GyL
WhygZcG/C2OxLwh3Qtm+f00h23Qj2SwXr1lB4R64T01UHfXO62W4j59LNx2JmTOASIX3WAs0nyMn
5ptXUMfibUtE/5ly1raNT8Y51MHxUBrEO0/t6bF+HoUT2bc2EQxAiBdCxeSP6SjMer3pZF73YMEM
HfCaVgzHebcn1jDX8sEOOmVoiw7VonGFU4obgdY0f4b0j2kgwH5T1onMiUbJ2XrsaU1/bUJobH0l
G3fkMQs7wzziknWSJdD5WDLfkhZFD7vj1snIDKB/V+TgMaEqne42hpHa661Og/onwWu8YnFEJv4I
vQh/mRXAgNJy/adcuMeQjYLti0ZjsFpi90Y70KsWQX+B9cwmH2TeKQ7G7LPhTYwHUePdcf6r1auR
Ti26E1DeiNqU2HVxU2ywhv+YZ0v9JKLIA/wfmN66anDI/xl4U8FDXjgGGpZvEWocg4jJtSXqQkM3
3WCaGNhKrDvw0536GXaeetqiRQLT4ASeXinN8gEnejNewk8WrdzUT2C/EnTt32xD+VYKXxfQW6ih
iUUDXOhw7RznIRHYEGK7ENe9gI9dnaX5E/XoqzUeBnRQ8Wgq9LlpQJtzMYUhWUYRO+mW8rdgsjL9
B/5JkLK/GqNYNJQrIYO/7XWpAVSOXJrr/WMFnDF+DvhuiYQvAQDBBZD6isrLXEeK/HqGN4ji3XtW
BT7QOkpI1CK0NjPB9fUvr9GJ5utdLlCYydPOEuTsdUmb3KJTtJvrZL+h93ZhjbfdhspkMD4ydvnS
RafLsFuZOoth5jZuTRMdgVwEK7jhYpsZ+QUWPupZjJvLdYp14SjAHgviJtm5afSBSEMbZ9WqZ6Js
9iT166JrphJwTZJI/gfMcMtcn1PvFTzEjpnCOoR7FvZ20C79HFOJl+6o/2n0feJLADFeZ3Yysf9x
7S/knRzVEVDWiSobXK/3wyTq25yruKcVQtkCfWo9rSNBof621pUmBrG0ZdskPxMdJJCluevI9ixR
gQ345Oi7BI8h3iStLgaasaklZDtJP6RqbdF6DGTwR4TpwuTbIvyX1A6wYMlaa9riiygTZRhkGu/g
CN51Suv0iFT/g2eNDfKBY4udx/mzo+ddKc/iQZ/JcYKgYRHY3n/9mmqoDZZa5g+cEvW+ADpFPB/5
Uoao+8FDZtSWtzK0Irhx05DZ9sd/pIWLAJl6Ok/GuC9nDcSDIgAyR31M8RKvUfgTllXAT9B62oj2
3F8/ic2QaV017GbquCdQ6If/BbG9TlDTuip9859WOypOJ1cwhxac08sWQ8EtfHbVjfzr3LMphLfO
kghDHpPyHOzXqKLyuY0Bz3WJJ5E+OPkOUllecs/ghJTOT7ZFMG+luY9xB4Yu73y5mQqut+nb/5NV
NrhiAs42Leuo5Sj3bSNYBd0UBfDMT70319UB2sqcJ/ARQtnkeheuK0byhB6WOoMBLgxuhCwLmsPP
tBlf2nCVXAw2Y/bK/dv6R1pSE992Iskq5QFLYCMlHOJe/0jnhBKeY47CkLctx9y1DCOgUyJ4j80W
Sm5QplqM95FSt2f8MNLeIFCzaqZK0LrGGaLOgosa6V0Tnj40g2/bZUetpsPJ2vBL69rlYk3EB661
yn/rBiFgL754fYNsSdyQ75CE+SBazC5S+KVQbWTcsjqPWZco0oTM03wqgVT3d1KX5HigBg3BRAAx
Bq8XgxFt1t0WEsZNqnP2lHSc0f82TKSb0WVbXpFYPbm4uzHqZHEf58AQe5ZEyZCaULlJ1VyD4vlj
N1aH5TaSEAXKYE2DKD8/pRa+0blyICS0dDE5jdOH8qcZWp7ZD/qe/PV8RUVnXop9MvBLbRMB553B
XYgviWQ0iH9QM5dMB3ar0KflPGGa10g2PUXknNvIXgn2cF67tXA9Aa9KX1ymux3xJvAoPwul+gS9
ppGDntlpfWbhkAfF8yM8VHr8LNvmdnvOiLYAudaQC+OCFSy39wkGryZKVmtivo1+Z73cQ2tkm8k5
nh+xnz0ife4U0CSHUFLWrS7Q7OlnFScJwxsAOJuVYckS9zsGanthgpNTox+am91OapV6cVoMsBlP
m9uUG0LXg9pe3DHxH6nv4ew7G0tElkoH4SUSskULN8tjywgGQ9S8EvMs/LBu6Y1PgwMgttHZUOi3
Re0XPKqa2UDOuD1moe2yjOzbx0g7v1gL2DT6RO44mNa540DHTmlelqeTXBUN2d+S7H6O5q2QhYE9
lPGxIdD8YDfPyEJvqALbcjjAL8uMSG3motvOAgZm6+3Ch+4rcF9k8CyZF50sA+TqPYUs6co1XQfz
ngevIFoLOqmaQwUtAguchjrN4FwHv4WiD7J6DAMEHuGZuTn1dAAow1mtmwswEXgxYX8cFfIXPNmo
0nkjU1C2I7Y/p4LA82UOQ6/MMenk+WKFv0zHArM1951MFMmp/mzczmqsgFguKRN7fssIpF4fA1Us
LfZKSFJAHtexDoydw0kioC8dM3CKOuA4339o7md3SUSffTW5qUUWK/n7pHmehXLQsm7E71P2LjlV
fgLyHvlI070a/kKHqcxNKOrqEMYHBRrSb7Gte2u+3Sk6zZQ9MDSDKOwzn3uzuBnB8QPm0kGwZt8o
EMq/5V+ZoPg9IkP2Jfw2fUplTE+uU/accXWrFDZifUjS9J/hW7Nr2YPvcNab1/ubnPhRHQkXM471
7EgWuqWxHNbjNIhpgWGvZIM0ebKqTq6BydEMMIIvjTKfZhlSD1R0GAI0t7oMbo0HVOHOnNO813cw
VvfHOGvmhi+INLVcdIMuizBRe5U8GTetKm7kwYpavHocdnHh/EgBtTFqqnONC+RbkJE/ugs9LHIw
phPM7Z7WeUff7ng8TmA8g2BKuXERCg+CzKkIJLAD+MJ9OhnI1HJXrw10BA/TzZ2Jpmz7S2wV2gwv
vv6GGIYXwgGl+gXcQUkASG8QX60xJKPjVSNLHgXml/Tzxsgq3FUIVhzRggTy7E1Pf9ByJ3/bfCYR
iSHqMiRK5eqY1pMIKjYR/w6E76/QoByHc0CgW/fLJMIfzQx9ohfJnIuf6sm4mvcmuV544ASMORmr
AlaCJPK9QucsAqFxQv0y5vL/sk3gsDNEaPGmycyUzK8EeAhooDgtOf9sxWbhKv53Olefc9mqnH+5
LewDP07K5J7oeoG8m7OnpywUXYxt98O4qG4eROEyObISNazYTZ+pwcrjcXTz1f7O7++I+vn92G/S
MQhesPIAvm599DsQlz9jRGTG8kgStEJiJu5KfssHzom+ymUnovmMUM8GcZeY+4D7Am50o/uZb2WP
zYzhEkiegJ7mI1Dx4aYSHPKBP/fwMmjTdvnXCQVKF6vUl/voKgSPbWFVNDtgu8/AjkqsQdYWE9hg
RVE31r4fmj0i4tejSq5j9ikpqDRIa/Sslzz2x1xLQyAvaZPURcDlrE6EQMONAzGzN1JPwDXAhtAu
LrhpC+4gW32gkwqxUakVLnUGw5Pk+AGu763fI1eZuOkJOKLe0OFtWBdecSSIPmmg3XmcaCKeWpJC
ilfZVaxDaq8jnVcJ6tZw7ZYkBORCWCjotacP0ZS7Otsk18n3zXH2v2ZcBuWiWVZP53ERP2d9LoYE
b1Iw+vtPIYZJgCFJ8U3nqamBIODkSQk7+/oOZkNm7RJM4UpL89NzzLZV/A5dexHUBxYZsFYOwfQH
Ua6xH7CcaaJfG/1GnfvW8gheRba5Tj57Wbiq/JbCoX5nTHzOlINwr1ItqtMy55EFIUFP4PV8p5aF
pmWeI5FoHf4svuXRbNQf/6uv9MghEagXjrhbotJISEpdxJO8WOH9YlwV/YzlT4qJmA3PiY3UcyIb
3pEcFYlGO5P9yMW2rGDXM3FmhneNobXb3k3Ew6EMx7NV14bLw+pIshnE283cyBQSNZw5Bpgk9bMm
vYLb7K1o4DQac4cfK6U8WgGRzz513xFiXcpc3J7Jm9zvb5PJqODOFjjKu15G0CHwv1i9bclCJFG2
tV2cWrs+6M2yqtaZtaeUR7orcuat6DuwaM52QIEFxyHupU+90p1JbxIjrOAEz/txrGfa4iIH5JgC
ZyQCuEDtGfGFupuxOLYWBb+HMqMMEYsNoXoFxhcJM9ZNnFx3F6bg6x3uCrRlcP6GgQnQ9/gA3ulh
PlGe1OT+B+oOdai20xfzSMqRiMyYsr3627wlWxiafb18wz7PYuNvZ5As/UamR4shWA0fofh/clbw
xZXzerQQCUUr6z2Sr0RRdq5aX569qocLGPl77ZU9m4YoI4G+/Du9PGhZ99SmqCqF4xhMHHbT1eM/
Su1zbtiOZfJNdlHmAq00BQtpnZDlfzbeLguskRKlJv0Y5+NtbVfLxaE/ISetyPN5dofm9fxvJW8d
lih/cQ3zch57IxG4GZnNIi17tJV/0HnaW6c/QaUaDjcTzNSezIElAKomNPBXWkiJTYkphMAETMbP
QMJeACYcdoAkoFWnVVQ+ljzxeETkrA/8gQnEU7WWv1QM3BpWlli9tcwxsN/0MMENeuWX30RViyyN
9cHKTBikBrfL1knXvVoaWr/mxvvUrfnxRadEOnm54jtLc/QHJgXfaQsmmvRYOGASS03UMEuKvJYL
/sHDCbzPwZ834h6odFxs2ra1rTciHwN92WKUZU3KZo/zAGIZwk473CJYV/whUmPnUimIhQiVOWSd
u4S/Hg6flrqlnamWS4FR0vG3tD5TdaPhmDx1pier6lbW8pxjZ5Ite4nfQ7/MHE2kXW83oSD8zjii
V8VtNoJiiVvuLTXT0oZ9P1HlM6EvI2CAzyShMrktqZLz4aECjsucZOqmQcdfTPn0A+Czc06ZkeMM
oUMHcU5jHU1o+bn8YT17c8ZjtBjPCH8IbuajezDImjn9yBgLVE0xkJTQkKBQxo/S52CJjZ2qP9OV
bWVqPr8JZpTIk890Zr+XVF/e2Lb6Aoo4GvfXTJzZfjWz44PJ2h9B4TkG1AsKZHQAJ7AaQlznVT4t
Uakez3pmhdHvLmWUNm1aOJZKli2EqdY+YaRcMKm5bZeEZKBXyOxuYvraANxWN7JFY9k+wO003hB+
Bc4bvtmJeDyUY6ylndarhvYRsQphc/dfjBQEn8/maOEDZJA+CFRlBTa3pp9aR1336vrw+SZfHG1n
YUEzbOhIe2AZDMi48n1TC4nHMgS156OVOIeJBbF4gOICiHWEHNh9B6VrS1BQ2P/6bt+JAv4hikzo
z5czG0plyPpjXPxf18KWXzBFq8/fwJ+TipFfVXu0KBQnxMrnjrDPMCI9ms5gAtoW7nYrvXsKCE/L
40Dbrnh17lFVD3M1CVjkQygRJyTb6ZCu/ETjeClVd9+omG1nSNwaviv5lKsk/qcCNXfxUUjTNk9v
93J9ohSTtqhYg0kG1pQK8mHequuiWWTehH9iCj/CfgbiCnZygq6TgapDvyn6Ol+LC31dksLzTOZI
I6GCwl+dZHQvdhONA+bdZ0c05i/aJ+A5Mi1TcVNaLICG4d0KFXLrCKn+ulO6orV5BtnX8wMbbCw0
mhlKmK5wQ2pDa+qXjfJJUkYLirGyFYATGJRExry8YY+I+pPPoPkKIxlzlUMdviJCvUCtzxACDuN0
7UnrvP3O9UL2Mqd5G1C5zt9ZCK+irdv4CWNRrPpmfmoe8emXpI4iTIyvKsQLjAgbMVRx+NTCq4M9
JB8i8QP5I+ecvwUk2KTK7jY5JFRZIf+DRMLgmhvk28vpSurfrjpruvaDN9y/WAq80CGBp1QkKrI6
kDXrY49MrLjcBou75SBWJAyYkpN3X30XXDPGnWhEO+Vk9gkIbrnKU0ZMu99T+L4sx2SwugyVex/e
3/TskSaPPq0RjlVJGSh43Gdqif5jvx3k/FejwlkO4ZYXcoiLdi/PA+yNwwsLHvbkf6ndvuKC14Kh
yny2Qpxj19drnEj/FYLZZPAx1AcUM5d+bH48HbAQ+vF4LXCqfkE2HFyuOMuopGxJKvEHRQlyIbZE
ORroH7AMgM+UWJM5KzphsCvkvPAG6mD6ktCGBe5BkrhM28+2xVQbMnAXRJw44EoFu3gwXTzAC8t+
VldL1enARnTMJfYCvsoF/GEBr7z+rafnRzQdn80FsC4D3ypMOlFNJ0SoEl/YDpbBZHi6e/vyS9gG
8OSjZxs6ibuOh+TUxkIDITERPF1KF8ZiHUBuSNuZ5tkjxc0AYfZzEtDTwP0f7kTiBSoEQ/TapP3g
g3pSml8ZoZvK2UZKETG9prnaIeMZJGW/tR2mMgm6Ws9UNjww4p0ycJ7jm8IDOY6KYnAMt/nguIxs
olNTKMt+isPAnch0x2Aoh4d5I9XRalyrkd/HpUSUuXt12wVVECaofcRqpSuKNfAQpS4irFb72jpJ
35GgI/KjsRa/TR19EzYosknBi8fjFLrbHpDrKb0j9XhdMZxAlxb6kjP0sSzW7mlX2QUh8Neb3r7+
l0M/AO3aVGEkHi7bihCTgmloBqZ18N4vqjN7iYniUuoIsOQ7VSc0BdIO/7GBeLVWus+6jT6vk+cP
LPBZVlXxzvTVtYN0E9vT+G+c1Vo6Ew1R/N0AmFN0bp/gmkJiRbbSRIIEgtjEYZfcw0gaXnx2R3s8
psPUHaBCO9QogOnwGLRmqAb55mih7M2e9zhx/E/ZCUelcis0jAMAR7qi/RX99/JhBhUNqHfA+jeo
ydtHuShyss6teNIe2IUfPBDPVD79D04k1PYRmQgg0QJ1lhHeE8Avv/0XD9F4HvUh0yp8JyIcPm49
hAdfl4vjrbc3o7DRqjRCmzZVa9VERqE6VC1HKe2SnPKkSKDzulg5nmMLR5a3WWTF2nZ5JjB7m/It
Mcnafk6eZ9o4GGTKtl7LgLaIvO2WL1GaKBwJ6nVzpA+b5bBtWeijpDf8w8lX7dbnQt301oWE0aqG
YSwdGXjSfiJY8ASqrr+kSTCqfqjcNKKBvdglT5QnHiqce62Vff2gWwP29dGxIgVvZslUpDPgsxKT
cp2VQHJRQK/g94hXxd7UK5Wqg0w3uaTcvcU7lb9KF9K8KKTJPByrDb+N4hqZdyxih2jrryhKnYNx
VLtK7VGfGXXm0+MS7tEq0LE7lfDx7rTY6zkHKjO8qf+XbasDahxeXF2SajV/Y0XkCrin249xUgZk
3g3IRZdSQRerFWO0ihHEOE0U8+7RnVB3U/IC6YX9WuQy/dlqGKsubrkGC3HV8rn6xUUQZbbsx29e
nWXZIlFSX4n3xPJZeL/3ORKupj2aZGHhVyytwihXCjjfZsnrML+23pec+AarDtcfoX2PAhuK5yL/
KzmyigF6fzbOWjLf3TGYDGoVIEirwUw129+ucUajfN5tF2irgOTHgea9irLLpoZw7lAPsuAmi4/U
kQm9lSVRQj0VogaPCICQH39lFHEc1fXuA0s3T+jJGq9SwotWzJqDHYU7mJj1s6VpF2teslW6sSsY
QbrkA2e80XGmFyFczReqaqO52x6LnjuPrunScpcpn5ACCF7At9wTwoCp0g/aqljQx7JWyqaUwJh7
eowfHUPbPKLeKPmnEivxpyVx4I8rgiPecfoM9SFifuLme7yfl2LO57S3oyz9dgnOLq8WWTbcEOHC
9eFq99lVg5u2kmVU8vyMgN4JByKG3HPIoB+ZhVWycDmR6kWcvIng1QuyoZB8GvlKqlEbO7lQPdPg
VGkagKAyMp08DTCC111I9RZQV8HW6iEgHkCOpMC7QQIxUAsjKid2XDuPjicKTQHgCas9i/X5m+lY
MG0b1+pQzk42lgsWDqnFSe0yyzWC6SYLUO+eshCAXx5V/9poXIobq9ivaded1zRUzoh4CdwE3N8r
vIp1BSVW98jUs3nNwtsnbEcX4TB/Dsh1bY8qakJK9n7024a/Z5gzoNQnOsgtuLHbN04aR4CLnNN2
emtMl1wTNBTbpplNX2Wrt407qxIRrDDzk+Y4ZBPt8LjHUoREOObZuhJVI4z9GPZpIJiIXxiSs4S0
WqFiAqV8GqXNTK0KEA9mOMVV34WLM5vqhvo86o57Q0xFUK9odCDFxetOHSRm/yK+gALlkFcK7nyH
fUCaga46s9WVbZZ3VDrc+YRGpgmYjpyDJldvYzL3/38yYxb0Gm1tvBbNgaNUZx7AHHmTsNNlogiY
d7YLOm7Z67fPaiukOGKQvWmLzCeqASckHeZy2mSpCWtAfSu8sdcda7y5CLbvOkkO0IFPADETDUku
FEJiGsN61h1Iqs4yVlGu3yK4NGiClYR7o5RuJ+V12GJAncWS7zAbBvRpJ1pu7UzR+l2ybyLYA4ZG
X2ctK36bJBg/mJ94VV+4JnaR/zNj+vD/hMXgmrmRAc1m7PvKUQDLkz/O2gO89cGVDButH36aXI2R
7hcK/Hku++7y6L/6T3cEGyqJQ7oCY2p44gS9x40gPhS7tbBmJiXA83BL+ztjsq5D5PfxeppJxbsr
9L+qFm+YNJJp/2MZLk925UtHZCnExvSZobmYsk239E5kXWD1vzqDXvjqhgGvO7MLDnCTazZokKTt
qey2OSWMcJ1OpmdERAlI61EHh6p46af3cW+ukQrDpwvhbXuwBt3RytQHfEWJaigz9KARuKFo+wGK
D4gN3RkdSq76W6PP4qX/fdUTk86KGKzR4f1lI+zxQkzednquLLDNUZEkpy7ry1yxbXRKKt6YNdxm
LTqs/2u1CKpwL/5EilrDi48uAqhla2ufjvHfYjXQwGy4wYDY/saPulhpIh6nNTkir2s09q1ZZv5Y
H5wY6eK8yfXU+XKXa+nF/nhRF4EVcrkwFBmk2KrYFVbXVk4aR7h9DLMSXttlf2QNP6OPspZT2VL6
n4Xld5s2AcEvR0aJ8PwJTTyWd9YYlnCnl2EfjfNAmxW+NHDuFxSG5iV6tdBOQVwHf5/KlvlE3YUn
ylbKaXZukOlPgoWq6l0YHHdzJXdHpX1muU6fNXteQKOPbs3mTMfN1+8Pg2QATSqrYw6su8qOTi6g
XfHG6ZIjU8TGq8R4hTlU6Hy11a/sTWBFaVpdJGPlGWKRvy+05reLZ10dXDTfoibM6B0HpvgpR66z
r0W6E0P3CVfkdPGFSexWcW+/VubtInQ99cKn1EcaOp1vanUgLIGqbXJtdpfp8nesJ3vuJAaf/K20
lEVlqEi4wFJ+N9QQVK/+Hs7pHB0IYcE6S7CMKSm1oZ4AW8dej7rDfoAE/7VB0RC3mqZJg8tPaYkc
RMNQcry0TPXlctkyY0DjW3Arb8krZG04ScL82XncYWb+29wcXnM0klPLlK0lv6juiriuOndbHmwY
yxkmQ0MVF1jfTKGKPHrGq5qRBZdbBDX0s0EgvNI/95YRwEKjkpzuXYxgLYb5TKCSBWCqvwklzGtB
pLJi7dAXTD+dZAZsj1MSJVIsXXi8poMiMnMC6AvkkRV3D/ce9g5HSrmo6QH/ji8BSezDoxiTuCO8
6MBuOmgAmrzXO+apdmT+flyFHOIGPFdLk00ZqvbnkWpZOzo7rKH1aJpFdrAR33i32B9ifPdLCmWQ
sUEdUd6RFNfNyajl1EycKZ1rrbuqdK/53n6W3uEg8K3CQh6d7i5Zudd2eaT3bq06LDUIF0QXYC6u
qqKCKBPaJWYrAQPznwmbglN37cF74VEMtJ8oqycarZuBTAPZVRNEN836OzUjOpdrJPTALoUZVSe0
o09BjVFknqnW3JhX73TrhKzLdsOK3QTrk6wsHB44sxMNDKSekrGVD8o0XLdu20nCVXP9OI4UqvvT
Bhws1+u0kKnWYC9eMVzho0GG0F8XMj+vKWILf4f0a8460bu1nr5K5Iv7I7ZvXzxSh7qiILspt+Pr
nlOh0MFX7HllbRspcyjwn9uW/dZAHfMCv0KHBkCJXgRSGylaKRYPn4mzRx6pxSfGoWQOs5OzGu7r
1QGCbuYSLzcE3fxeN1rOFe8YYO2ttWJIR/JFlKtRrAKvijTLX2An8Eesp8vFRg37OnKoHTdZNXws
pLsgMHgDPV1LFXI+Z6evRliF1ajD8RRoMsOLuiZ1/eLhTPc2wpMuE7u3jlxI+WuoHSgEp324meyt
x277B3H0MJrsiJOjA+5s9mRCatplKITfSfUmW+ETDZlXRF88AdDScM/7Dz+Jno5ZS5lliu3EYDDJ
QuEwyfelfcdmlfTqwFg5padxni8Bp9gEJrx23epnK1EzIRZxUcz82hRwEVpQ+dZHFc8wHhH3tVFv
rOcD7GB7DhmK+fzxm12WOMDwuEjYvyPcruv9jKpznSOgbKHLd8SXZFJxxGuhVaZA/BmHuvk+FJmS
KdDl4Yz+e5Im+/CDQYnIJoEZEoUlHgtS67FmisXvRJpby2p7V5LRId4gE6DVkyShD8/c6KrzRXqy
7zBhRAm53pGILCC13QbjXmH0U7E6epjKDBG7PV6K16a4cNX0kPCt+bmROxJIP1u2dggG1ZbVa0BB
x4VwHAPSNE9WMRrqCNi4s/viOFsPfJo9XaOhlp3QZeRQ7udKmxEzjKE3xpbHJaKJ8j+JEIQTBXsV
g19JoM9k7CUud1KDnoQkWu+tshNFznlYO1lF/yWVbiFifwLc/yJ85TApEKrJHtXyley+AFxcu16n
YYj/ktnCqLmoUgsw+QJ2MO4iSWg634XD+/h47QByFmTd57lh+/UOW9QWmLEvBhTzRngzcn83eNRR
M44EJj7ctNa5DA4TJoAB5qME0LihdhvHhT7JjYL7hIKdeYFJDp9LTWmeKtIjkyEfiNsBqk1LAkeV
ZQKDGSFjQToWJtzPWY6fqBa1ECLmI0soRpCCwsv8Ysw986+ZZRhEAyBIL1VoY6dK1kcujbGcO774
wclvudAjwyixanDpvU15fEcSpM0IH/splrxV35yBkmzdIw5lA68drh3xtMEshaSyGi1/5UqHsz2C
wXJuBmPJ5FiOtceukGeCygyt5wmzcED2CT5IEaVkZQidugazNr/WT7Wgg6DxM8Q8Wn4KhDVR6V1r
s0ftcJeqF8AlohZNZBwzmO4pLFKXJfJS2xKe0/X+p9l63C8TQYefktnsT3y7NOKN6xAI8DLw+bpZ
uPbya67mAmy/meT0EQbwc/bTnC8gcCyqv3I/686T7+f+71a5NWEd7TTiYYbxUIhW2Ob/q5Ffo3oW
8/6v8l8d/t7Li6L1eZQ2YuDOIDewXIj6N2q0kuF8aeKhThcG6yYP0tVZ3QFeldKx9cSMGTBMxgSN
leHQZ383kTHz2YLckA0l3JjDy0WmVYfz/Cl+FOqOUzmQgCIz+zzfjoRyXX9MHle0NIVni/Yzc3Qo
v13hrX0y/GgPNkp3ndY1mWg7ijPp6BMs3vxIbeA+V+jEiWNW+zICPu6CBbd8L0k47PZFf/9QFREk
z5yJLbxm87Z78abzb/AjIy8k92QePOqnh8PlPN152OXW+e2pL4M42sAKcpPzdt7AKd/LqZtsTZtE
5J9HarwLKKQG8LKEIUmsOGeyGkPtPYb4BfbSBNqXVekxfitvpSAm/gR6h2a9KI+rlyyljyssxO5J
nMGLlXV02nESJY+vye6dKxS+ZY9ugW9fUMCNDuYr/lB9zEmSlMAWFddglBuzvK9ktWTOGq4j4hDz
du/rxcCfFXWYfRlBAFl7n5/SlDWlonieyxNMkf8M8i1vcUnEdQlgh70mgmHLTAfUSnth2DPNfu9p
LttsM8QluiFGSlRq7p1IkI1+W4aDT4qhPG1m0234ANsxcP0Vkvsp7y+StAn3alyJJGRa6XfwjMSZ
DFfsLmzz0PiQvqfM7/8R1C4hyC3EpeIL2WPX9V/dFeKQWCx5jDfh2yXwD2fJJ854lRxSGF7zceeJ
wcTlllNnPJE+IASisqlBnGazrEnfLbdqaf0YJawfb8+8opeJbZFZ72szpP1Z8ebq/5HXtP1YkZJv
6Q38+OBKhHlbnTU91QemAFpi85n0u6DBcVXJHdY7IwL3zojK07DRS/FTHsEIaybz6xKxmzwE0w5d
SyE4OquwuiVDGG+4No/U+inrQYtH2aHT6JUNobyZlpH16vB5PdHxGwkXrUesp5OQA4gND3qEMuAL
36LNNdEGIetcEN36pSWulUFCXPlQHP3GJY6uhJlHRpCeIPEbVR5ZQVbyVAwDuOOxeqJcB8FZk0Df
SEJZVwrCmlGTdyhSjpx7KhW2whNG+ukHJZDIm2ixYkwAZZOfE+UpVJsbx+lfGRhi7Xft3VJBXdSI
nDabVYnzqYjxlF2QOrfX9MHhGmiRsFzn5HE2cF87bSYSb39Zfrn5bnkBVQB2aQNvkaXBD17bj/VN
qrBDrrWFhPn4pwxDAU6pDXeAILIQ6m7/nKR/aggEDCND+bHGMo+mq6MQexbJdr8kTgVjkFuQTpuQ
Pf0VpEsqqeo3iz3R94QJ+Y6iWQOWq/LDr1Swm6lKe8pf4ecvZXzdSiGVnTz4T1wzxZcnxq+oo3qy
sHVi/hRm6RlsJ8DzHn6rI4UxKQgC7ZASEOrWm48dP52fjDdemsLtO3YyqbAQ0Y2IBPijhYvYHWUb
9bwe/xYq0bH9woR76/P/g8MMX6opMlWbMAvd5CUrX6YNAjZ3OwgVvwUKfnLjn+qIGim4Us4M3TAq
pVl+Bjph7FYTBkLJ2zlwctyEHJiOHMhjS6t/HuGSGl4CBFoRpJ33RnHVPbpcaEbMG7hOs9d1tbEa
DE9IYfcNEgaZ5zg1UflUEevwSnFwCa/U4JQmKKxg8DHdbmUMUwEx6Kc+0hQ7HzgOBpxWFfoTzqt9
w0HPQnkpUEVFjbBfJKWgeI1UzUvYmHfVSV0NDfTIOmuaBpk9v1aYpjIOXglYQDJc9+48axyR3KFl
p+Oq7PIBjIoefLvvzdVLp6hyD/pdkJx0x23FLzsMrcwR5ACyK8muUKZQoTa0HOs9OULNL8e46P7q
Occ0ikr+8u3ABBfA/cvLcbKxitfX61O3tO6J/6hOE4s7qmn6qx3hgbslDT3KAG6HLZXc0jOPS/Gx
OkVf0bfZ0enwWagzcwVnFU0+vEn9bq57oXPnUcXyhlgSCGP0Gorvq/EbwdtsWSAsC32STJzDId4T
Dh+eMRan5tiYGtWVkNQGcJsEgg+J+rkYQqtNWS0L8ShICLSBflqXu2ovuERZd7lDiRIE0vl+RNZ9
mXyjX1Yn3LoOe3cJiQT9GCtJTk2yR669Ib5ES9mnkNjBnY2hXlxkUEVnMgCpDJ9PD/qlLox9l+4z
Bvpp7o+vja5WZSaM4/gj1cJGx6nInDKGDuK8XrVq65mYRQM0sM59LegTPwXAKirhnqU3rH9oNsGJ
NH7IbrKaObl3kk81KL6xNKicetid1WViGZMB4hVJl7iaQHF6jw5Qn8SicGfR7oXBMRb4GDMJuKb8
9JgkWpoBjQ9Crjax2bNVEfcEjMh4s70hgpTPyix7d5+pjolZT2qobB5gqAeezrOzEK/mVUvpCibl
ZHDbJ7oD8jYwy7IRgpoZP2ia/cIhC4dDv6eLfnurJB+q8ffo8deFQ4fTi0fvv8IkXtcOVO9ukTub
NGvLsiwn6KASBiPbd8YrmqhheAjoknDm6cJrV9dnrGH88xb+TjUlXaZlZ3iDVONS0Vv/dts/EReH
bYWc0laImmtKwM5JC1h7PketyvNT85/PWuLN8fZ3UVAGqEkx8XUuFLQcxu3lcMKCzBlDbTOwfX96
ShTEp/dQedXja2NV+s5E9jSiO4PRCo38Z3Ut1E4dC2UcPS04zZBG4WVgnuEGq5PLC71uKD7vFerI
n5IPv3Z2b1T/ixxrjXQmID6PMXTDQCAmlkg78UIGehzE3fxWqGn7K7NJIyDi2iPR9tRFGCA8AXyM
AjvGjGgm4nQ+7doegw6yVvY1pJLwBo5UZWLMlQ/p0irBOv9dP5tfAsuKnwcZsxkBNZ1vp3GDgllx
p64t4QfukxnOfyrtxwEJcKpzcIbc8aaHZudntQmLXZ5RXuzVtZmL8UIuR7VPJkWgAVu04R1zvjAv
ZBFGElMJ/BwsFqz9E60Z2pKOekeB47tSJNwujo33jhZZKjl5ASAeMvumYtMePSLqhhqCc205V44L
T5HCmtwg1zdCkL4kfPKKB2zJ4Elp69aZmOflu/xl7x3MoZb9eQmfxuzDhOvxkwo8DwNWFFIM0hi8
tnbQu9l8Jfy3NE797QOhfWK55FjuxSZwiF06oE05VjayWtdrQPNGlrwhrM3cOt+i4nfl8pqUezAk
e0CkQa8c787xRTjY/E1fQJD8vPfNbAX7aawVTui+KY8/spTKcru0gdg+vzGfaE/xyXehYUwJck9r
Itrfx0TtB+5SMD4fKGSQ7zLlYyCLg4sn+TrIvC48zAeFeQvtBbHK+k9ONeociANk78vAGI3wOxwT
mCVlPd9YLYXLwCFqfsqpCzxxDzQYlRSGMI2Bf9eUeP8uVo+dSjheIdwu77JfnJvl91PjKZvHeXeo
pUtitGSIG+jgqWbTYFtGAdUYVGmpla2ZDomLM1vv64QcfDxof+/dAdTnn+W2je9xLhV74QUmIub7
uPYetjGg5K4JvyqFu//a7ovAk1LhmWGpuKqnZPu89xg5dpiNSiTAzQaH4bx2SSQGR/CFHwENZkfc
x0wv9+xgd2egDCpovCVkA/21dhRBMs8jV40hpfHymDF+FxH+ozV+KJPYKCIK6bBx+6U4vtxCYdST
MTm1fCD/2u4d1agiVneOzF9wVqT9G6SEuX4EgJeouhp9pNV4m/0pPZweo2LmQY+T66JcwnrLSXbD
0KD18MaURBpJlEhByqUhPFQpqWLSuHedq2eYyWAj8YY2hCu6yilbOWgDSkCvTBPsZ9F3RWszK9n1
646yMZ76D65PUkC3czpvmAVUnNQ3RMSt47hREtuWRpW6vRhw9O3VChn3fhEV/J3UwfskS4MrNGpW
zTEWzaoK0mpE8GyWYcfF/sMjQq+yDNSePwF+vdTTYrYU6aKTO4LAsmOQrMmkf95ZrLgwRM2jvNPA
qicks6JSrOwBaf8d0ma4Zpl1Mh21WR5oE4Ic0pIqXJGLVjWHpm+iSuJR5rLbctMKbabXJeVa182n
v3TEwg5pG+KeDZ2e9Zz/q4hCD3wl4U3N2DQP+Sdh987AjOIP1fmOBeHWeCq3PndA+ECkcZl7jDV9
AppkeJtwQQu+KTWJNvXnso247/q3TbKllmORN+P5yyxVcecRsiQu/JqLRUB9ti6yRKa1/v4J9z/R
mNH4X59Isxbye95HSfG9kbdh4H2+d2TIhJBbHinO7IvIq/JHArFUVC+6LloeC5wFqAiwj4RQQ+WV
XQmMM3LpwPYLBtCi2YbIPv/7c/+8DN77s3HqqLUJzoUR0GTGE6JwmQeeweRhyCBHTMSyveQ0L0W8
cgBpmPBMyM2MGcGH8ASiyv9g3ETGsIT/lBlykpJDCpBfh5BHi+qcnUBODBAo1W5exCnAW8YRTFXD
TA7W90rEeCLmuCTlQAmR+rKZvGYFXv+U4e6Wm7X3CC3y/qcR4ThHTDb4tlmxulOkYqFzzla+nutk
HCjrSw/p9fD9biTA5Q451HQ4NYFMwX/6tlK3r9ehCBxM6cko20ENJ1nXMlbKMUWTT2wAp4U8eXIq
EaH5ZPhsaeCIOMpgsLLxUs5bs3dsghu6adnDtOah9G+FuHKq9DHP7bI95JUlNf9fGJyviewUeifY
sizIzJGzntlnRuGNVSm6imoKs6ZVRCGMbwRV7j5612t0Rg2a3CdU612uof32PKkJQH3bGks26eOX
GcV/bF57sj98G550zIBCfc+db8zPm6uPyLHdNxCriY3Nt+RntPRTPJz1CEMlK6dw2niuNTtuKqua
9iNn1y6HZBWKce98S32LrenTt7JL9jWzvd9U9EGNvx2eDYjA0knRUv2Evi9PjcxtB/pQKISkoxv2
Nb4+fJy1CnxQmGmDdwVqxcVMfSS/BdnGl4UO1vece2TivTDmbae+kXEZDL4CHqaBrvPWGerta2LZ
dKNDvU5beVWkJA2wc+89ORcRwe6bWapV0XwDSXBc7D/pH6zx1mkTPm9q21XxrCNthlom3P+KG6QD
uNIdtZ20ToJJPLwCmmtNEbTy13acmie57Y8++fcAhjm0BdW6FTK6+XNAAeiEk9R2wzwp7pooIvfU
nUHyKSymDRM61sM4GMeQoB3p1JzBKx7yXE7a2f34EPcZJLwBtt9x66c7WTFMuRMJoqQ5cwjNlGRT
X/DN2L48onzXy+c0lueSeMd+0RpfnmNSWyfaFDng7gazQU3mMzTPf48UNRRI1Wa4kait8N1UIq8c
Qe2gKHV2OYPOd2350YuBh3YyeQzPmHjfaNgquuiE4Y1fBRRvro1ThzRbmJyHAFWaU53b5aUeO05X
PR9VgXPO95eZzOPWrNYMHgIi14He0PWiaLlpzGnBrl5/JlLGzsYZHbLzqc1waBFPN81E4ghGePcu
k71j/xCMJWlmk4AQT5b2GbF7BgdCOpiuS5MGGTkIHv7CMq3PDpq5sZ/MGhkwZp1XZYNf8mhYj5YB
QiqIFBmXwQCCxmwx6vATeADRv0TdzMObdBkfZwtDQaXnYWzIvNLTCa8kyz1CdKUyBBZny4rpQVMq
PyrYfApbkLro/QxhMAh/tdu6T1cR18Bqa2f1LkFIdwa04gJNwXEnzrkZluGvrJUQ6m4d0iiggteR
6/4+FRFGVMvJvDeWOmW/ZidG3TUVzMdLc0BDV34inZqJ6AcKM7z2BvGpU7toO+8y/8/BJZyzMzuH
903oVYoRNReSekHi+QiccnRNasCSEOmRY+FkUGDG5beBIa672/OMZMGfScaxfTNGIB3lbh+1bqF5
CI0eunlA4ZU5Mmg28aSDGGIE/gvCCQI7vnz6o2hRbFVrOIip43xW+jdasM4O+Buun+syC7XMu0Ov
L2F5hkYCL/dWH8Mld50Hv3ghustQJq+gcCUbRd5e+neIjTjC/OH0xNSyQkXGsN7GYv9FdTGNPBaX
FiT+AHFeEDFFST3RrVjyJHGKYHEwIqQcFLh6If6K0qpInyWxehWX4j22A9gaSaLeBgel7m7ZDiIn
BqsRFAw54jd4bTJNnNwyajL8h2DRP2WBq+dF2ESU+HbGAxIv18upOmcUqPFi7Ab+tlvi+4cW8aQH
uCZE0vgL4y4DydbDnecAWra9XCIDuiCJWZ9OPN+3bmvt7sHpD2Q6IABy5vfJGciV7M2nQQfMBe1K
/Nzv56KC2C3MkmTZuhWWw6J2BpclB2GlgxDY7NfsB6rlz9xEXB+UY5gmathvRiEtbrmq50JertnE
Oq53yP+zF7GQBEM9ZYnSs8x63zH1OYuNObJEpEaeeucum1U2zw3y9BXyoM3npL4RH5+tOaAGSU5Z
MsRWW/dxwMka6UpSNB10yMU2SK6TEdGC13R5pvXvpvu4ORMq1uE61ZSHHqnbRX2lN2CshODcWpHx
26cK3gnNaCoLczl1luqWFmNuJrUP7PVfUgmkIxbYB4eG3x7bEWQq8vNbTsQDjCW/RWfpAH+Y0oYO
Vkp1EWHO3Fk4pkSpyUiK+bfLkpYU04Hv1tA6ggAbr712GKBx5UIOpySEZXe3BXyZ60QG2b/f5tAW
9tMea0540mnu9f2gByI6ZBZuE5Z3JjuKBDpWZTcWyhkqG1d1gXuw7bx9wyYdTEyC9gGTQrg/1KKj
bPFzzFeyfcm/iZty79Zb2mc2rSGFgWPWqQNREtfthtek33267JIKm6kdm1EzV7gVA9/6k2PF87lA
A8KWN+fKv6MP8YGsWEYJAkCz3j6ATmWE0X2gxmS2LBrGDT4d5nibwaky9R6h4+do/u8iW0RQTk8Y
poGNN15laKLjebZkS3lRXENPEtN+4fdT/ujJeh5ZBCPkP9OMiYRYddkzh9+ajzXmz3egWR06WitX
gz+ahnGXXUCP+hqQgMapuMtIgE2UvEC5HRzPBMmpYCwpcVbCnXf7mNXt7clAerDnIT1Iubt3axZb
3bUpBP3EH/wYMnwnk4OB0zprsGjgV/eyQHCpn9ZobkDDuFTGMiskrHrFUssme6kId0PZDKXVEbVJ
qFFja3UkonxXYUXxBSmev9wKGrIOv+ceV+i0qOl58RvUf3Rna3TquQdsWQC3lb139VOmcX8Y8iyf
idlHHo17t8zfE9xCX2iwZ++JMGNzExCO8NYoBJtYdMExtiRFUFJmBQ1kkcRg+oaVN/dTIupCwXRj
4qagR5jAssdpVUEcZBBCXKSeK0frDN5coD0U4MM1Pf1IWBX1DSmnJrCpl8d3Z2pWo4tEVib3gZb8
EcVQeDzwqFKETUSSPh9wdh4aIY7qn+qcHbmR3Nog7Seo2gn08lakXCJPRjkrH5fuSsdTPGjnRzlo
pgSIL36lgwxFfRh+S+o/Jl4nOY06jJCylqQ3gAwuP23J49zNP+U+a5yrJNstkB2z6/mYYLcF8W35
0v2CbVxBgLW4nFa5qLnZRQ0WIQ8tvPXgivGJVz0F2b3iIRRkMdJJlhfklTPwbswxG+VWILP8lCAW
3jGMFL2SBnCCz26hu6KM6rfbyJxTh42+HJ0zPj/RaRJUTeD39aZZe1/8WP/Eyim6tKRX3b6YyBpz
qEi7pKCh+QbXukE7lWzuMDJUaP2xIFsccfU3jqlRbqaFjj5MLu3VUb4FQiGCXqVcIk9/pqCW9EGe
OLd4BMaG1wUWLzqRJQVsQhSbDXnp4ytoBrFV6jnBxY7D03GgkaHgbwqua8SoOfRSurDzS2AJNi6g
t1jflifIMoeIZy2HSIth/hUDtsHcMJxVGHlSSNdu5TNN61WdTCvPoXDeqVb4lD1zuX5FNVzu9Xs0
zyXiojKWKOFWws8XygslZvfKlcLHgePZuRR+LGMzmQspCDKP252T7sRrbKwsrq/vJoXOdv8CPg6H
m+MUwdZFX0teZhuVkBnHuyvKYhn7Gaa8ulAAZOUvwG1n1mi9ARCbtAKR9C4yG8yt++pBQ59KrxmG
wbb0AuY+eIz0HSziU8NLXD/XVHXZEp/3iCGdvFKECuAadW6icKITWCAY3GFIjWugXvyt3hATOZw5
jt7/0g6nLJUvMBYTuzvrWAYPaQ7urHi3VAINLvuGYSCITeWd6+HGNF1jCuagiedrP5a2sJNopr/g
+QOsEoL76LqJBv5HCLDXvZ+HnKC7P5xI7pccIRR6CwbfRcv8GDXntU/x/D6hm65UkWEiizJ31Wrk
WCARcU84WFox0+t5kpqTVXZ7ConhEdcCNIphABndefQt34gcR6wWOl1G5CqDEAGmZUsfi+NfU2Ol
o+O8cFmMMk9yH3cDukwse7beysa0k6ZlqGJbvmiP/rM4NHfz+RSqIbGk49w2Td1zATAUyblm0S8m
qPHP7F6R3BYqqcxjzXSEHjkMu6ITSWnqSZ83NNapj+OIiOnyFovvPkPlUWnVyUgg2XP8Hj/YHTxv
Wn6SX19lcfd7IDvNuIGV7d2hyAHKUAM9UUiUwKthGG6IWSvRz/o3XZHAwfWL3uwEeSIZKVgZ/43u
spVnWJUTuc7sLbVfyVY+U4gwvQn+8Gk3LOxfzPUubPntav0whSz/FAVGBEAJwfGmUjgad7eZVkQq
YkoFsY5SpW/V8o0jrzVsUCgGkYUsFExJ7/wYYzbfdXXK86VvpuGCQM+Ui2aR7WDWtv7wb/5IhAUA
aa1TBdrJf+f9bTSvKcec+ldNdIHP01QyyKeGYnxPjiEt6W46QToM/FMyCOqLbwnEA9k1jg7NOs+s
RQF55Jy3dBdu6NfZa4hHAEuCGA1ZeldXSumz4Zcv3oPGaxx0IPr1IsJr2V+vHFXOLai4tRwfrC90
mL3WULmCSpo6v4ZN44Dm6cFM95fmJOfix67lvNLOmCkL/QqPZCMn2Nzc6venHSDdi2/HC5qfo/RI
vHkGiN1lpf2G/yDQ3DqC/WFn5USDGhQCrlEBPB0+KPtvWyCa9id7bpjIDYBDdz9EZNjk2MQUjV9m
W5KqmqNVUjz2KlRJvP/hrQnd6XjLyl3Msotclc5uSXfR0v2hn0yJK3usikPnvbJ48n6FDmpgEOyz
X4yPWcPhccQyCyGaAnOTvzlbQpXFR2xFV5hZBHqHQW43xzN28jrZdRYAZTpZ7nluRaTNir7w8hzi
iMAW+zyX1Myqvf3+T1CosnpyvMvZicdWDsGLhXtRLzY9CIR2QWMo13g2fyOtzaQLHXCZt74xRrkt
bULJ8JZ8LT7/CNfZS402ipHwSYemhBrQwk8fUYNQckZjUcMtZX2n94f8n3FnKeIeTiOx6rk+U8AW
XLI9Ogj7Tz2subjoxhXZGTtsjDqJK433Lts1zX7cvv5WNvd4FHRdRj0m0ZyoIo5WD2a9o1xu5gUE
P0EdYXEkutU4k8Y3KDOgkUt/9DMCKOYpBs1cI3v/ka7LLdsidJUzzmiPj5qmPMLjLptSXEaG9Q35
kE4j0K3ajRj2B2qeUVzdPpIgl2PbFXcO+jKne3UIDWo16jCY750ApwOklUqqmcJ7Qi0zxSeVuG6T
IESXUw5oTSkw/oVeWQTl5t7aROgvjM7lP8AYNpjzcVzFR0exsWQy7e0BDrXObg7OsJECXkFwFqhv
r5b2eumKXb4If44vq3UdbNyip+QkS0sAQbNN2E9XsYxlCxGy+tCXeSYb9rBeImaGoFA2xXPVqXuX
v9CnW4x0OMzIgwKgLHSBtx0TMv+hd56r0+HKmPQ0fYgqvmqA3cyCV5tjgtLIsTyO1CE81kaTIJLp
9a9lAvwFBcQFWNMKXKcmDfSmMd3Ird4i9iYjGbDLZ/hbiG0iPjovyGjQpc4GQjMyqpHlZOsugjRH
Lx5zOV0rqx2O9Fky9/CO9ITyF8t0fBE/0UkMc7o273fLQUvwwtWi33Uj5sovyPAIL+OiL1iJ2f8w
sZZZnfVYZglW09dDYttPeVbAxRy/FhWb/Ar59AUcZ2UJSL+6glDoB1tNm+KxiPJ7Q2FWSaJFdW0+
8gnSZ6iPHdeD0wcYPwboDkJnNO0CgYAayXyLVPwUreMa4oeA6ZXjmenY7JiuNeUfC/LB0XlBUSqr
Aj+TjAXUV84jRinU+feBGxthOI+7ZA4NXPvBp9hovE8zLiGFo4I+hyuA6dYXJKpvREJeh0511F9y
q05nsFlENEgKi5X7LVrzLTMNyXyQWxsM4B++XSlRK/RxeJQ5IOLuBW3mH8fgWA9FS3EbSHdBJMZi
FgcJilSOCXMBPqAxNlRIbACVf+DW3IGl4co2fCOV6vcxd+1an00A+vL4PitpeHAMms5QOxIdubSr
IP77zPeWlEgODZul+QTyfzoEMEkwbgGcyyB1bM1rCC2Dm4zxP3hrOroC33v50cKnC5uJ4RvlosnO
DLtj1gey6FKFsIdxv+6nXE66NxlwuZCOpfwfaNuu00RoByF7IKpjliOxGASYwhA/Mq/hsmnE6C4h
nQmAXvkqOQtSSB5FUN/cCbgqbDQ3wFKpumRzxkrtq/Nqi1Kh+3wzwvdG3mmKigCnDBf58mIX5jkF
e+rlK3Ab3gfIVcfjAH9tANEUUJ/QaN2f3EwgEKGTBDY5gv6Rsv5X3KH7RBGQlRO415G6Cxbe8kwI
0uSmdD25XT64mCrFVLQ35rCN+NX5xSYUaBhVnIVwQqze2GKkQ2V31EQzKmLIXLdC6qFwdRSN0TJF
Ym0dyTKZEq6UIWf8mawNRj3Mz9r1TtWd/m8OsLYAq6wx+kb3gD2QSX3ZwPd3LOBLV9WwRur3qk/Y
mJJJysqK2doJpJbBp4Tqq+Pj/YXg9dzKe2BBEI4XKjUxudvXJQWTsn4Au2pEAptjYLYt20k9smHm
B1lx1sUbB0J4iNu4S4wEwLsSPoyv3vMzbmHzqPgrMt27koa+Zc2fceuroj9+3P+XKy/GBUDcjGG4
WI2j6Mitw2quQntp+6YKElYYTC0QTaqzmohpNLuiAi7Oh6S6G8h/9b/7oGy/bNv8oosz9WEmp+Hh
8kBNHUHq0QrlymdYalqDC/hiNzAC2zxCuIyHPjFOabVxrpz9yyZ/jboRA/KiwXKZobtR2/adWO3z
Mqe9FLho0mDPnzvqrtuhnxUIiRHH0ruf8H/pKkC9RqMvtXHEhsgOGRWXxiF800+p/7xnnc9ZO02Q
DbusUz69OkDFplM7TFCQ+3nXbmDFhXxMqDXxXLozqtKxLH9FqDcq+jwOpyah7OVchpby3j7+cu8U
XLllbwJhM+WXcN/1qHexdUfevXymoZIZObKcLDmWMCOi3IC7cgv+S0AqVU355ZbmJYvdh3+XKw+f
Q8uAVBHpxqBM0wXrvMgwbJQ/ULwZ/Jg0iGt4h/S0Dl/etJ4BjNUYoO6DeVerTtO3k3iBEQUBGa02
QrMr2Ou03Xc2iXGi3OLr/ERj/NLTSp/R8DEz1KunN4uQ08sy7uLxLB7bIChKt2bIOsO1WgJq5DsE
HuZzqUe2BM3k3aQki1nMp6KwB2YssuXIpcl9Bh50yjXKBrdAu1CzzVrhHsOWaMFfsv3xIp9SdrDy
i7crFtQXncKaHMCk4SR4q6WrNqd9k+IPcBvevQ6+sL+jV/ta6GVd9hlYCG/Rng7oOCNPgGKNBW+E
2IEXEiFJDQnQbl9ueI4uFtvCICG+nz8yjaoFOroNzatoEOmtT5zQYTmQ8W8u055M9lNyPwamelP8
LKhlFJgvLmVFh/RwLgn5ODBkZwR3RqR3IoH09jyKgyOMTOU1cpdv0BiNwdW5srmJ3gRwwcqP26G4
FHWr+NGqasIZcUdd2wFZrUCzjTooW9IUR5kV4qsgegvpwaOthFz2/dX97y1Yb5GeSCMAnwv0oq0z
V75wuJlT9kISUVF0bXwmJysDt3jGiTO1OqPvuXy9qxoINbtl/CFGf+16UY38f5fMAYBkG7XII6kL
47Znz6kY7HQheIY2b2RYTFwCuqMhQvFOU2LhQTnW1/8JGYrHMiI7o+G8j3VQbq9S7nCaur78IDSD
TdNpJm/8DlWqrHNSGU/dVyqXADZk/DsXbq+BHCZ4i3zNpDYTCqRfXQAQetGY2/Ffmq0DFZYz8cv6
R9it0KOqj+vYgv8DvcGGRSyzXY76B7n+n0r3Kd5r5W+MNLkuRSbq4N6b6YNcRLpNZoq3C8NS7pib
EVK8jt3IfYCIVEEmIW4Pri8nm2OtrFNN744xHiNkKnQQD507NlZK1Wb/ccYwxEDjXvcYzjfS17yK
X3jh491qDCLClQ4StuV5cWBl2iURecZVifvfP5yS+o4Zku0v8tHSJ1V6e+cpKM6fOhDYbYW/6Myv
ZXzmVMcA4/D2KW2jW6ldge/DupeISLYKIcaTQ2bnoVQic/WpI+JLERjlCw+EC1HWgmqAPnf5SGWH
AWPHtjn/YUhm8sYsa6deuiuTLlmaTQ9BFAyXUDX3d4Ze/r2Fb9bLbdDnOOMxYaHodZ72XBluIg1n
6b6b7j9hKDMyOg2Gq4DWBtj10UtEE7KDJxTHkC/M7b9Qr80YYgngMm2yFpWG7Htxf7ZymO+01XxB
I8Pbauw/ix4NX1Lv/46n4L7n4z5zazwX0SwG8UZFsx9Z+spM9tVGjYCXhIzf+Mqxzs0c2LFR2MyU
czQVpVQhuNPPMKH8v3uxqizqypXD7Dj8HulsHeqHKZ2sdAVkYtylJTh48Fygs609ZPldqhw4QxyT
JvwCVltxiNpIMF+Yrhm3acoGnZgo7WWUSkysVuLw+8fxz61QrparRow7GlBTPEdTRtk1lAJtSxZH
1LWiEhrBWNxVsqi9Crk7baTlZz5W1yI2vFDBUomSRjq40IAjLWR6kUmLgFiFkOyZN2BN7WiX/oAm
vSEAAaF7MGjUhZJNV12GcwdifqeqVYj1FIHqrGnPof9diSRPOqI11bw/bwtzunp2yytvac3Jhnd9
+LiZKzZUKxSEDFrPYHHAJ+lkHrGLLi2T/EfIDd9jqbzr1gj5J1502uEPiYv0HmVplNDpxszDGuHl
y31aETEOy8wHBlOaj3wDIDVYU4y/V4Y3Z70ko+T1qdPk2TsKInBdEvy1i1gfv/MX6ntWRHxtV0Nq
EuatbNw/F4XMJYxsmB9EKH2wOvwUD965TEJxg8cK6F9wA10mUyuCjOTuOerXIZrH8XakH/3r6hCK
SpnxFsFdRLvNqtHL0EAsj6ti1jYYzhgvhEOiiOf9IplnDq/DSfZOfGyyxSJy786F0zhh0664ExHx
LWJagzcPrD7zYXa1KGOluHGcGb1Dws9dPQe8lx+VM7sDy0eCkCBSIG0Kua2P2DlEgbHAeHOQZqFa
2niJ80OfwbjoEx13EV8705UXd7YTfxSXarkfkINRacxF89IPgFoUlTrRIomrcwDWq2M5tm3R/sMr
akfcksBxW5ix7OLDg8LNVZanJp3lWfXU4vGkUwPLGlMgBVW3L+2EFaCieyO4WCXUPSp6lPvo5dWF
g2vvJSLSJhZW0Ko6jPwz6iVdSNfioX7Lblib1VMEC5ZUxP1usakeYZ1DTRZHXz7cnjdehE1JejuT
4IDC8rNrKu5rA9Ofk/1dydlziinRspQ9W5+vFYPODqsZdehWKF6AywZgdyDnAvFr3uS40/YqLsSA
5eVBQcskBGPXnMm5It8TEkoikx4j3s8ikCHpdODZSzB/EeAqcub30lAMKH5Kw+IIrk7vPyR37maT
tZKWPcp5s7zqfqqtlE8Xc76Rsey6kiQppmHDATFp/PkRT9qbKYo0J0ucJRr3Q8QhwKA/nr9ByM2l
MiyK/CNQ2ojMDeuwRJWxmQEuwxMxc9OMIx5OEx/1txxTKI7arpyHnUbx5sfdQc3TWZaSJIF/EyUc
CKveMu9X+xlHWhkaWC9hhEqdZvdR4Zouls/YxPBiU5jzZ0S6wCduyirj/1s7JQZk2bJn6jq8FfFH
/oqgDfLoFeCgc83JOORzT0V9onoJ6l+xT0hbFeIM02j5u9gnk6hl0koVlXeM6fgA36neCrkzKOmp
vIhYAJPjDIuy45obszQo+bf40WgBj2JfSTya/iyIqDCY3/Np4rtUZavKMXJt9Pyl5GOU8ZP8Vud2
uNk8WFXEn/N4yl5Xg8BwFGh6x9kCanzDb33TThPQBUkXROLPoZXXnPQsyRukGbSaHjfbyID/YE44
bu8cx7MtAxFvWY/MUBRM+2aKfEuLfTvbSdmUMWNNpl2vPUj7eZTUK7FfwmlSge/fA1CARaU/UuuU
s86jTGIzcmTOE1ukivU5OMKZs+DBRP5/zTMy1zUYyPp1wjAtgKi+HzC8UFu/nSPPzwCFLGiJsnVK
a21M3k5NexpxcNhsLJAM5pp+BxeQ7IMyTHU3zkpSuECEDntzJsC9HhiMRCEcyeuCnGzwGOtp9k5Y
q0XSofQafdbta9CYSPv69cnYPgGgzuZwivLqNCrwuNpTbGwoxIPjXUGwO62wcoEBcH59D7W8DvMU
4ZaVn8he5MU9toPBZKX0P2wxrjjBvNqxwTzzSrIeMiSRyh7pCbTDD5YiX0i3bBluNWlQGSM2Nv0l
PPPiXiSrU8QmaTFo0dgtli0XamYi95LzMgMIk0UMjz8FZHVAKl17674yNdHCZGBChMF4+KA39JuO
9XrezgLSWMF6mgUlhNvprgc4PwA4Gtj5w10MLJpDR+nS37wDF0OIRrJLt5HffrX0FvGMmwqA1did
ZV933Z8hc8fmO68UZWQMkNVik9cMFeyxmjPuIX/PB3yVTKSZrOtibSVZgnXr7rlXf5n1G/5kZPdc
2s064SOgAoRGCzZSlKMHE9caY/Ij+X0VucrssqzwRpu/No2lWsfPwxXSPAqS/MHDNFaY5nfAfC7K
gUf/Necbv38hD2i2xDQs4jr3oCVqGrfu3fK5mz+rw0PXk2PbdUiIBOrmTrwJ33lwQa2IOm8abA15
vmZwE1VjaXXnDQTLFZFqBNemlhk63/cndldk4WWl0DKkmB3HYPz3KoXq1nNo3zCcwY9lCc24K13D
M79ZbuMZ9w0ufmVmru8uLu/ZFcM81nlLQ+9FdYo8DDa2zJkZ5JCk1tx56kSac+kpdOIbiqz00v0F
JccX6w7aFSfynrfb0u7Dzs51f8h18ORYYaW/lsg1/kp/xpzZ7/qEhXH0Y9kVYpoPZnCzd54+mS6S
MJOYDQXiP6hQum2XDI0qYikcPXqQrDlPjE1onrATux1lN/W7AsOuvVUOb1VGMf2NSwi4OxUijUqq
3CWkjEIA/iHQ9ywBPpIMjOaIc0USIxmh5gilozpRmh0QJzP80Jyt+lQnmBPiU+IRl+BDi6+c2n/5
/X9mzjAyJbcYC91Ne2K5CwDjJu259rIVHeKJaGCdeje5zOzEM+vwmat0BWPtRob/FcyD8cvSYzKX
yI+JblvHr/MGIuKgPAAWUuvnZOMiCD54WhLJSOS9bce3HUGAygU1LTkcdUKsTjRPpa/Zs4UkohvD
A04f5avAa8Vs3Kx8+pd7BcC7Utx/K5jE3jCWHaH2p8p94on1zafBOw041qf8RO/pYQBVKMChtEzi
y+jWhEFNWDVHCL9CFef+TF3PnTf3JTNXkNUGfpUdkYXahFU/BaUxqDIscaBbYSUKfNS413JvYN05
ny6oadlBNhiyDB+7a1V/9NeqtpICDLcxKXLM2mer78YsB7znGut7bqas96LslPbXZS9G25Sh0mW1
llIvI+vzXtm8v9O5LgoaxngHDcqinFD5nfI8QVjfirOGV+AjsFQAOa/N2fINBBUWakqsfCB1UlYS
2Cw65q5wNuLsRPaG2RtLlFSxgZ9kZSOj5ncNki+5UTw9Y+H+Mn/JxqCTJI6crLHoBY8ap9+83IXj
KkiDLwdr01AmiT9a+ZOHlCfijmP7WKLlZ2+0DiocKvwNXuaVgShUiabYWHsD4t1I+eXksMAPLfPa
3U5zWQwq2BA7yygwe76dWMhfFvP/Wkcv9P/un089k/P0tvbBuvh568zXiYJYTpPA593Tg1DnbezP
u0NqV0+UWhtfo+94qUV6QD2zQu3uSjaJUZvmd5iVX9ciEvQDH4cpYKSG2Crrv0JSNXs5z2ylzndL
4d7wPzhy7VCFQFetnYzewEBmNfjC4GSx2zMIEurEPbwRKVJasNQwlZXYC8+x465lIp/w2yS7xsvT
T2ITlRBG7LjVptp4jtUvGtbGQiLAtQvtaV3b896by0lXJrJuxPTnTv4WZ1lOKnMtRPWg3ITOOhY8
gLjw1s0nZsB4KBjRnaXBhffLl7pmnbDDx3rHwOliTFYEPcsR9laUfFhPHzVlRrCb6P2vjEMZMy1Y
+G4e3kvuEF1lIxI0BzHPJbUcPPd+YS7F1O8NLNMSY8eQ+w29Pt47W1BmJJQPIxG23SGbCQ84FrQt
/Wy/tOwKA3tSCk6mHOL5ESo70eUrkVckDDqZYiDsiY0p/UxZMWxFMdz735ssNbkGF89R0F1FQzdS
CAND9wYzXDXWTV0jBA3g6t4KsWRoW1flwVxQELlGzDL5K6alfRitxxBoTGVfJqedN+HrpcEJOiLP
fJlgV3AblHPjxUIB0U0D2AX/8ItLDLmMHPVEh6EUR3+lYItQjXcN6KGtKkceo18b3pVu2iOzrYI1
1kwRo380xfIZjm66Tv1WdVSR2VP/ALHd7/kiq1jGZUNKnlRNGKjyTPSH8fQ+jRjDyT4DIlQIvoIB
0u9YozPs0wXKYJ0k9DUHv6u9B2garOz9V8sgX1zloqFNjiAg1s8ytWLrexXOXAKnSNzYywJi3maw
xpntJJ6oiQIiHhha+1xShTh+gHs+Y6ImPHx1CCdtpQENbquqp/MtwifupQlO9UABG+1hbuZbvy6b
YL2eRUEk8mngJ/sv8qqOVWIyh6BaYGYVG2DPkv7CDJxJRfH3ccNcM9Afp+dcWxlYreK63E95mshL
VZ6ayPXGvONiQTOzRsLcJSUSo0us/F9EiVkVEkPgOGGlBHyFiJsxuz36bLX2T6xY5jQJWNLcWe0D
kWld6cLG6PRlPY6c8EOss9D3xDTim1vOgrWCPMPn8rX/sPLMGebqqIXYTu+B8xfVbJPN4Mx5VqBE
uML0upSVhs+rGpqWdtnej8EckIGykVKQvhvbsDHc8k5GUcdRs6ptFJk+xNr1fCagVizBx4wbmcwa
eD2tZx1r6k2WolsB1Essrr4cJWGvIhuoJswZ+tvKuIsj6cMoql7Y4M7e4Guna+rUTie78GaOcqy2
rMFWN6Xm//bWJu9S85dZ7gMJoCqs7nUn6lcUzZboRxpZqeg1bkGAbm3HTPSxfPjqHRGR/GG99Bj8
G9pKxXnppZC24GC/V6b3HPWVB4E+9jDBhbWjCykvm6vQGsN48zVebOtaTqH8fG15DbzmSCijDsSX
zGlBfWq3nrnE7kyC5Srvx3cJoBScfjLYmkMY5voD7WC5WPaLitqEXmCKe9bb8WsmqTZxvefgBNxZ
34F/+Vfqf6IkIEcIN2l3/FkzNq84RlDHQjkoYdwuuzw5fDHE49gB3NYpLd3IHwFBO8XSAcAF/tcl
YyJhGo/y2gJEIkecyAb/BcMv9foFhyeBJKuu2Qss6/AiKuKTHzRTij5v1ESC23XpagqtScqppY0U
N1+0RV1M2L9BN5OUUjv+u0aIYmIqQtOHhu7aXXvFK7NyE3QjIdMBy6Bv/ADuUvhz+nGFGrjN19y5
u2P8wi/smNUOYqdaf+3WX4uYAinqF+BZbb5K5xq41DpRvUkoDNydqXlI8Fj4Bj3l4MwW4NoYz1xN
NXxRVcURrgYV9lVuVxClFYWy5h5BzfQZdezydBNMUV7woo3C0/Z0M2BqEmdkMmkAfhjXrN8fGqv3
w/ODSNnw4GFMghnXjJTGLEs8fvkYr+ba8r0wdozeg24ig6wsB9F1eAHEBWvHiuK8zHnj6g/ihXSK
TL5jqCRU6A2jikKCRfMGny1M2h5lqiDFkPyUng8TD7zqsQpNjTcyduo5Yc3p1BSoMRYFJMdPF9M/
OKwS27U4A5B6n4ZAd3lqwGkkBINspHQwGkYY9K60gQ+zYAo3r4SnQ+0bez4vsocH6eEEv3JfE2fd
0lE07etO4botYPh97glpFsCJNeQrO4So416+Yff1DN6U3b9z4YXsSVrVgHfRsUuudl5udwVAeroy
vBNPUG8/Wi3/54UOCuTM7UCti4exerisuZI2x9GU9r/J9jkvE3IsJK8kPax0ZwVs8ZUFkzdUHEmp
V/AJyvQC5eDlgxN232wG8GD9d7tG6Xqcct3jHXQ6UbScR9ipF5rEDtmnFPpLUSZeQfh3F8xmzT2B
Bzo3anjN/EWklY0Dk8/YDdOPqlNhlpSjt+Ua09TLOeGXC6dUob3I8Ci6iV+Nw7y3nrFdXUxM2Fwj
eeE45qfUSTzAKPoAr3lSjLqq3o96c5gZ5jGTrBA/SD0GWm/cMqZxu+ekNf6FVooCJtbR4Aw8no6p
r7oZhSu2CcAMjtnuOWqBBbR1sul4leiRn2WvRnmb6fCk/QlmiKwG3VAB/k+aW5E7FQG5xzyTtOVL
uU/4PojmKOM4LugQGgIbIKNw6k+N7FrWB4WlsqrzT6OHjS39mw1b2elSq+QntfCbgJ4gRBePvtKl
AGdBpTu/5hCdttzkLrQfd8cHa4MQZCbnxP0DWvGUKvEJ7wJPkGYDdARvpd95s5rG9AHejlooYyb1
ZBK069UMLU+QSyImlwmSGkw8Mes+qGq97BAFiJ+8GH+1aX37hh45bkV2poR5EW94/7j0WrD7qzf2
tUF7REdGGX0SOv4qv363c5OvKeaINnBZwpynZJB25Y763IX0OQ4dMwlgu4OnLz+jjWT8YVZlCSKm
dvbSQjlYZa6vKZHoXkR+7gHcvx8LLT9Gp6qaERivV5f9A8kKQRCnNg3jtJHXpF8n1G9SoE5hmejS
4BibT/7WAzvvVYuJZOuq1jyAH9AokPF4ZWpdQJbMNmOrtg4/jWj2E81ouA6bezkkhGQGzBL1i0Pw
AfTCUtLBNMrX2Vd/EvZnSDZGUgjOqHzIDlI9FrtRc29bIUxaDNufnLPVvKFBUUXLXTQsKjy0tmJ7
5/3Q2GlCvqujneB7LhGiJO1/5snYwyO7GqzmvWmpn89ltliyE/8lNeE6aMphxjp5i6AZH+rkUyJM
INKbGKzVsGVGVdTRADLAH2F2FBPM+R/TWfLU+hvRDoCdleTOzbALTCz/VLb3/fS6r3Jx94jF4wJt
LupO0RLOO3epu/pLCJB5IlH8ve2gH6HLQNSCRcrYTGWAQN9z1Xb36pj7WUmiazMyf/zA9pqNiMfL
mAqBZlXJohXEnKXZRNDLuVh8B6CtAxUn/Dxku+4+unnispPM45QtXxrOgPTc8RhYQdCS6uLyf8Z+
YPWSuA3nCdmB3DekSEjeleAqkk1q2QBTsh0FtDU5PsMvEfgLP9itq0Psh1RTOU6w9VDX7P/Y7D6P
pyj/+IJH48AaC1UhKBm7LOC4hVdwsdQFi1dj8NQxdZemlKjg9k69mOM5NEuqqy1cHHJNfCsnID+P
lH55/CYCitaHlUQcwIYlLlSVs9HlZvhb23CRK5zkQ+suHQCRsDwH3B/lJnrDpEgVyJ3H+tyVxVLh
xaid2sCxH3SXAibuYYf1312AL8EjvuTEcJSZDZ/28yT8jWIlae2ymwCOXuBNBzf5TWCJtu39emRZ
PpRABLDcZEOyLdFtMsjnxIC66pC7fiNG/ZWNlec8Av9nBLQMVvmEXY8QKwTiZCINevRCOKyMz97n
QAxWronicVX+RHe1TWNEECDfVOecGuvzHN6OcA7EBIg/HLFGZDEp/bySY6vSgHUUEY+JDXB8Gd6r
4/8ToW6MiK8MSDF4qKKKt5BilCnz9AKnmyjdwiCpk1aMsQsNXYE1eEjiduZ/x8WB/DGZJ4Nu486a
PCM88cmGAMe0oxVNv2an3dMCkR1PPV+4PLNhPhXsAsztK8ipS6e9RAoQ1vdBs3o+Zhr2GMZRdTbz
PcuzBJbkU7wvDRuhS42dEcJ8kO+6DHHkcRdAoH3c7kGQ2fAD5zuontZEultXyQDP+y+JOXltD4hb
l2m8dTzIs8/jc0fr45WziwQc6QdiB9QqRUnc/Z2cRYTG/wpjLS0cFjCR38dJ1BcpYJfL/efspOrF
OV1g0LYsUtMQNaNTuaR9kzYXV1pJxJlurrBM3YTi3y/x5iW2MCPv22ZXAu09ATMVWXP0MMmuv1UP
zwnA00PxzVQscYO9k60ge9UfvY2ldCDA5d7rUYs4PBvcHEnpyyCtKKmX3Z/8XcvAEzkd+vZ1p2gg
NjUHQWJuhX5tHdmcy4cF1vS1THiH70wh7diONPSvMDL6k6UKBRqnaopmTHzKVSj3kG7xXV/8oYTG
SNx3/KrN6X7VbxxBSvTvqc4mhjrbNKpjUCOUbwB/3LeRz+bNJ9YrUxNdVHOJGi4TCiPIRWr44c5p
5EC54aJsxls+IyR0doy7fLm75krrXI3h3ztBwm/vxdmxZOHYqSqBodk16uy+KToQUl3kM8zW6+9u
wm12rKtuqjSK/uKmLjhT8YSf/PcBDiPaKUe4HjEpMfExILxOCiPOqDLG4hpH2Rg6hpqt8fFfstSS
2451c6MoJsLKqOo4bgp7iXKgP/MrAobwCuKejSBTHqP4ip8XGWQ6fu4aNniS5RLEqSQ9Qeow1spd
zYELvB0yGeOGo5uUBK8gIFaI0/4GAYCpvzVVR06ctTMlbGhBQN5HVMUK8MCQJlCh0oU5ZtivCiwN
NkaYilOL5LvuEkMuOYrRts0Mtc3OOUIIl/GJ05mTyKD6HaYknGcMxkZXNED7R5NhSqh/pTenKpDj
C6yhXbQMwRYbwal6wJgQZ03EgJ52JpxVK914RAXUH8xK2kEWYjDm+c+8m/0D0hkYEuTGRnIaR6HJ
z3SDQSdaXB43nFG155esHdaQ/UIx7FjB+9rtUCPyukYmgLBXOUQ3RvMlO/g55zMz0huGAEbguH3A
UmUT8tdkFld0dEJBLZjuQl2JqqUSI1ofeernem7/fD4ye7xRBofjfm6l0Kjutj3Gz4ceg/NWXeIo
EFUjQVD0OIXAeQ/BsEEVO0xkZ5dzdJmJ09FnQV9Ot9ik6D9nV1+vEo/+wOJPyXWDHnBRWnZELci4
SnemfVTyD6VqvFqcmi9sgraJVdY2UAeufK0NaUbH3c3BN3qQKDg7+Q1Q1fjXTWj9PrCWPlcfU0c3
+guGjttSndxiM8KF7/2sU9RhdNaZwj97YGXR8Rr7qCGJFAL7J1xrBurirOmsCmj6pEKkl+G8iiFx
9+kdDPjdA8Vyikb2Uwg56mQjhn/DD5eHsMX6k2a3GJGItg8WCbT6b4ZoaoFZOWBllGcCflPsYU4G
fb28nrt8QPluylzar/mPlt2k9a+B5WUeMZsk++vXgZ7+hnIVwpNva0sdwFhCQasJJ1rluctEPoZw
cmnMFIFhp7oOliHhXh/x40KzKlFRdknMD+uEx5J46vGpqvfh7jZp26CZ82PxjEof8AAr5hJ47zW2
Md21XoFW87YwpPZiFN/RyifR1XP2FXUn2srIFZ0jh9DnjVeyyW4GGZ5eRJ4v+Tgz52nxpnPbtPXT
1kxGAXOZeBaHvSyOuW8pjWNKwWxrzuCOKjB+r7+mA8P/tMEiUBfi+3e8h+KaKDmfnKykasnkxLH/
ifaUZ/YXsUrpun8CTXYjyQFtdZLG2rSNZTeu/zeoyiBeL4BuCOxO6MrEDXyySghe7ZtH/OzTd1Je
NwcvR7c1tiML6xhWyhoy8cRy89UyHCTSfsrfIsjMBjemj1xHXtQGX2B3F3oqI6WcHqvdS2WH1Cyw
WQKKAnLfB6BP42sAnJ/FBw/nN3LCoHM66ihACqkRTrkTh12cL8R9hnwRcO6rIQqe2uxCSxmMx+Bp
1tY52nnQxrJdCD4bPaqygmJbZRoAoLf8+6oMzjwm6BjcX7IGoCo1/sxgAse/edTC7TKCZLuYGmMj
NbFJ3aEYR9NUUImZPfkej480yp3ZtR87F8MYNHj8TyRjL9Hq6Ym5hmH7nemrjuRa+lbFwPK/YARb
ppNpoDl5ek4CFFW5pa8fEkeKDiBLJDOTLOO8CdafiT6UC+5C6PEvyCuK+QFRNXc+28en3sY/AS1t
Z9s687S4kmsqzoImTC2/HnHsYpAd1M4MiAcsSs0wTYgZmppir8XM+Q0rTCuGN+IDutolNtksiM+b
8aoEPOeIQMqKQyWtPufxN8f6C3kmBoWFZ3PcSamm5V9frLOMAYZgzqQWnnVFQlfXnAx61qfWUY6a
1VCQTwDMRd4tCseYqW/4Hkwz0qhV7ps5pM5aFf4gh6ZEfG18cI396cHGp/3lY3iQXV/dubR68X7F
g4HA4et/MJNggYun1lAIRRhyPaxll0hWRO8k/rvM+0yak+n4X5aF4MCLDafwf87tCKL4Gbzcf+EA
xojH5+BAb7f29Es9X4YNwCgTEjy6OLnSHCKrnida8LPHW2l+6VLDTzpGyOnx4hnFoM/JTCofmpcl
LtK3+ZuSDnBxt8TVPmaU8HmEtZAbwYZRwCZE+klY+mzdNHFLernRyrgNTx10I2NeLtroRg4gTvXw
Ana7GuF/sqNsLZSQYktRgmMWPhT8GUaQjliZAqcwIFNJ7ZpVjun/YAzXAt0czAOe4iH5sn9HdptG
/lakBGKr9L6lVGR/NdYFkfcRJseRYHTFNXBUrc1nuWhlm02r+LHbeW79TfarxNCwmG04iabOridF
pMoq6vGpUmHO2HKcaBspFbfdHAq8WiA7G9AWMi6YX8WW1NsF6BSTCNvIaYIpbY3Iknf5RkPc94ru
bmEeShE49Tr80V90rTnA+e/v7OJFQg2D2VPF1yTj4GRrGZs/mOR5uglkGOQBm1SPdZbD8TTAZZyb
zUO/ltCKf9l7SGZNudBJOXS9KePTK4QP242HOlzNl9zQEr4btTm3/Kr1Eu9Fkh73P6s8FQi8U63B
8dy+mPPKCXZlE+u0Sl/KkAyz6d/kQnhs3nnJbsAhQuFdr8SL2FyzRw/Sbap7Vq4p6v3zkoSJLzhR
uDgVaXiW7PoGdWrHBg1FX6m4mDVRUFp2Faoso2A0mw6AOz0pjH5/qi/cz7aiAvv6tbCB0x28yUjA
xVCME6zqwLAwIiaTE898tmUnbHNnyQexUS0aStmqFUxb7XgRcSY1RnfrdzsWqlxIw9KclR2dTLDJ
5azhiJOGrZTuW0rxmXSUf9M7fgh8DwYFCVi42vP4m8NxbTN+joWLEmYzJTE4OGqZENKtE1F7+JI/
jd21NSQWTvvTxzbiHXqfrdAzy3FJG6ZoqpxsUOy/fw6dbLCfpfs920ps5WYHnO35aPSkCNpPYJg3
4EiFZM8GCwRNHv41C8izdnsSOKT4lkAfrS1iDCcQTGXqpjynPivNxColYPcs5/t8EXyZpf/+GVTJ
F6RJRGD7ZQakY4cgo7GNqTrUFM2k2QAPwOthb1+uKR2Wl4xvxtAV4GeoP+DUI9GI/Wm4swfno3qt
8cgl6sB6bbhILztwlwfMLqRkhFz+/QlhDY8yFCN0QgccFjv7lMTIPDNwWBywpCGGNIccsa5YYvAK
TwZtPT99NlkwPQSZrfqGC0y7pfEcPAszS83u7XoCPdTO5rG7ddjUHO5NC1PSAYMiSQQ5jAhTlcsF
IIu/YwfIA5GaetVdiu9V8oi2TZ0ceE4jTEuzrmY5ShsnAEbu4aBf5//mm9dR698o5Gv5z0y75oiQ
owi5IXIiuU9v39ysTQbWZsBPIRTvwuZkZceeB3u2KT9arutphJd40HHT0Bsculzjk7kxRx6kh7Rg
c9YmoaoaV53uBRRsabHGSDSqHEMN+9LRC5R5JA2CIdCduv/+xc5Na4VzQhPL7QrS8dFvkOWpMtNi
XiQJuxNO5YcyBVfOVGbl2H0YhuqvTferZ0nmlN7xl1H7SyU0qs5eCr6JhwFsykT/dfRzTgoZyv5S
k+k6T6PRk2RKF+xRqA9SFt3ieUKBG+DuTPS/V7B9lhlkEu2TzEyqzSpz21yjOPkkiykAMVQUUFi7
eFMAQvc15mF1RPzyOgDHcIMe5ajugr2z60G6upvF0fCOQcr6ys7hEf+njlgXGyUzWfyMqLfQvA4X
JZ+bUw2bqHbC+7HEjTrEmfQk2osClmcCmrME9opVI3vpwan04pZ/FbpqJoycN2j1j7epRoncPSYn
Z3ULDGleyDnKC8267gukHfVOERmyFBfFRa8GKW6pOEBu0tQ97Zc8wkXS1ibR/18oNFF29c8ZcHV6
WN1hEd21tb8J6yut+IVhbPNWqhhO0KYh2m6XUPxomGMY47DMGNXN3p+yGg2aWJ6WFOjLXinqrYQp
0E6T8xhfNnmc7ia70OgGk3RVsIKvZwVV5i9bn0xKD4TKkGle6GclF9MxbBkrP3w0toPQs9LAfJzk
oxF0Kn1cwDPEA1rdZv+zLdX34gxldIrqufTM89N3z4ui7b8L4qCeI433IDW86Y/3Ea2XTLoHkU/L
Qhq/wMzUL8a9Y2+DDz69Q7P3QJL5GVv0kbRXjLPJdzL+T4BIGgwumXLH5Arw/TlQ68HYwlY+xhM8
HyNmaiDC/IpJFFJ3gcJ5azfaZbQfeupZdJxMHR/nY2Qw5aP+sCLKFx/Mf4qr79waxQLO/6qv9KBl
THyJK8F+ibVAaA+tPegDA7fVRW+FKmJ5KFK5D35f0TyM4888SXkyy6x1wo7uJMDpbjIK0P8L8Bba
p3fZS+eefOGr/v/ngwNEmr0E8TTb1ZI3GVJxdbODmBJrFatkEjGaIl9B2REZgmQ1ASFyFSsieWyg
nxjBnzebKmCtaDpz12qjYzMYaTR/pMG8tOI0v7qZfNf/2MX+cg5s8O9K3VtPZc/166goHafQOoHs
HX98avyBzEf7JSF/0fEkLUq0UqqPslpRZ3d8l8LhuOQ6oC6KQLAYYCx1CVGM/+J5GcztUNfFslZT
ASS62vXlHzE28REZ0NrUUS72iAQuzDt5IP/C9Gn7eanokyEkvQRRwD/MZ+Z2cKhwEqMPB3eY4CDW
pS7jMziywMSCNu5yK7Tx0mK0qg5fvwLTby3LLb11SLowUmOuRG1AFneqABSZaMZQjwhMAosTAV/g
JF3IHRnrYxc3jmH6vOrf5iIBQuzzezN9PZD93oKgbvjGSPZ6Zzza3uD7koleyi3UOahAF3LQEiWn
DzIEMevtKbZqpVtWl15NqO2H2R26Fo2Ya+Pq6gN3KPRM/+Jc5OMTy93mbw1MzEtJWZVTX7KMSmm3
1U5bLwMKx9die51f6iXn/Z6uGPrhVkXwpJkArmVV3eq7z4vn9OSI3YueYTG8mshO4Sru4v6L4mbP
QBUGeF11ZjVh1w18u26CHTCsTlLWNdqtOJpHvIy0vjTAX2uvLhhTmAKR0Pay2yluuexbuFCaAuZc
544n0aA5MyypLznPCirkKONx3GkKa8/NSQPT/JF1aqD5ufJ7nzKfyjtFhC1i2hSxchvEe8wV2uRc
gB4ZNjfE/Fv/2FgHDTXWZQVanaXIWMsGWh3tFCBDEQm5aU5gAchfYrUHDX4UfwZzVGTkzw/1dl68
ap8EdpezQ5Z5hOyKw/UPQHD1eXQsZrRumU3rSMRHAbyc47KYMFzDV23C/1k05fYNbktUs/Vsfv5+
UL5QKJ3cLXCSlSleIQQaFJk/TXj+2diyNN9GrMb5HFEgv6ZNEwvfGBj8Jyj15C8wl1qPbz0rpAC7
r3YubELVM0dC65vSFnm5Z9krqokU3d/69aB42fOa7E3B/wlLivW2pP3IUFRPAc8XJTAbFmv7i7SC
uxWLKa0BHU1UDQuAs+/3h4V1oxSKsDJFXtaNAHAQ9RSyYDdoZK92xDgi5lIFgoMZ8bGODloySTht
ecYJ/wyl348XC1y+L8ykGtOtLBANJDFbPmOZTraRgWrjBqtZr06/MnGJDeX/TxR8W55zgBNM/Qci
aTB1+FT6rOKujuYd9ROKLA3wt/4FAFFxVdgW03GbJ8FxOVJ7+TbZfgKSW+DNim1DmzOH/kNwuMbP
5a/RA5HmcnrIIXgBkpWiO/vUPo+J4M/4HhDhreV3SiPie4bDzflhRj6d/mPpyEd5adRwVfGgXPKI
O3CNj2+XGEzVTDuLRwk7TSrA5AHtJ6BBQ+lx2d7ZH84/cTjWRXjWJnsY+vkYWnabfpSu6jAR1yRb
cGBKjhqc5tzJwtEcY2TZZE7LAlNVIUe8Eyve5xzPHbByxSS9SlT9xT+MAFfU8hjP2pEnwXYmlkwZ
uwIqDFdLIa6kmziS6tU+sDUtbJfTjWcfjBCEX9lXk2phSiCnGpjwu/c4ihWYxG2OVYD1LS2zTpDV
K3McmziIf+5sBJntXbtWj1W2SaPu572NYtBOxPkABZmXMgQ0tJS3emGE3CS1jAXoCHSrQOtMJOCy
YhDb0AfF65nVNyD6ucj+wxcNr4abNYZQhmVOF1Kq3moelpFivVnqgpAq+qXJODfnOY0320su6XdU
DldbpBos623S4Ht+vvlqZSiFKehWobsNpHtGkxoYjUTWCwgIVMngI9qJQFe5nOoFgbaZQmdXxLS0
rmB0zFUVW7bB4IcSGz1RvWLwutnos6G+fD1Rcalnw6fzRFZD877HjX7b84nYYWhhKq07GHsAt3Qf
X7w+Fft3LGXd+6W2gTeOHPbv18bsBEG/yIaGggwbCF0SM5uuHBdnXE7aGf2JEcCtsAFw0vLFFroY
jw6DLwpqTYfdAgul0qQXTlJPJzo/lKeAfYJTeQgXlQDS/li2v0m/H8djJtRxRWGVnPUxykn/buZo
jN7gSPHcnaa8t7Gl+HyREbsCWfqVwtHxzMu1VF2X4VIvUiMlFv01S6YieDjR7eYTZvq5BYOnYZhN
lZRxwaALnmeEoJ2UIhfXCmBdZIXbDkpnTAMhvYIrbqn3oTJgow+IqVT2SnZ5CUVndNF3wJkZQNmh
rI2U1JEL334ssif7nqzskD8u0N/Tb47CaNb6bJVbC3sVe7cCF5tv5OfH2zMtDQ9RLca8PUtmo/nv
N9jvdR1LvfIzJjuLaHZQq8qFPimDS28tFQENF1uOVme2WDdrXH+5GtAwhmbRbvwYAoTrePk5vh/M
g450xN78UcfPOV2WjmGlsgOf+1xd/dUtWyiympTD6SWeaXg4KlAbsQzHEnHgX/Da3O/uA768/EcF
/vl5sPpL7TAiUbsdSw4bk11Mv4GLj0UV0pXzYve2JJx8FfXiMVVOzYcc4LSnSAnzHlfNq86Bix1F
5BQJQjWMBiSk0hsFh6jUBCzhHEgS/vv/WBX1vyAyFbNouUTnQRkhk2zYv+u7fvSNU0pm+PSztx76
I49HBS2Xf15kl7GM8YswK8KLIVXMMe8nMxB0H1mEsouHBHe6ndFxiJI7s4kayTAzB2ZmzX0G9Q71
D9/R09cBesaz9pL6V39wEphsiA0ijzSdfAvlZcfpN04Zf1WWs2UIDt86PktP+9FMUn4oiCEWcywb
OYnLrWUVv5gJo+zENeKRHGhSV+V4KLqeSlRy1IsBVkG4cy7Gwqo1uEkb43IXiYvg51mqD6bxe4zQ
G4Jz80oam2q4Rjs67B6nb7oFA7qywJxwueXQD5/9gJIuTIhe+37jJdm1sR9k8o/nJ6Z4emQ023Io
x+VG9etnT6NkUKQc1egXM19Dwqsu74KYFUCiDGz44RWcqM/O/8hSaK3FyEmBzIQQcebMMnQYm/ho
H7m/LzhVyVr3Dxyy7uBBmuh2yR6I38qucVWftv328bHY8SqRi79kKT9RfQYebavP2+VbtjpP7MFt
s+/I9D2KJiRLb/tb91tbLOaQqzveh9mAME8kIZ48txdVQcraKpv4tHLYmUpi2HajKp9VAvB01I1F
i07owr4In7QYzkWN996fH7TIq6rzyBOajnU+I2rrqHdfnviobANhSghxJ5ov8f8HvV5mjhSHZO+/
n3AmI/wCEHIhgjzFKWMtvSOC9+VbkTPUy7GpZ6Hc6QmznKfPrj/XezIaDTOhYJsHFP9n7NmLw13E
DIuckRp0xYv+R0YelmQhhHv+tEfKqWpZs3AdKaDKGKqHdbHnlEDBnQKsOYj4bwpCvvJXwfpzgjA5
QsBjlM+f3N2t2+M2GPbjlUoJp2VX40HjcOrHgk14+v34nXF2Y0qRe1foYttCxpBwAL5JXyiRzxC6
n5eQKA2VHiN/UVHQTNeFfsVl1FToGNBl7VKaYwoAsejpFit4Lvl1JY9OU6l3gb5CDvemoUhe2UkK
qVdvdI/HFpnNEG0lbkcFiiZutIkhsejVbbKKibh1w4jsaZPvH9AafxMaZtZQ7yuhqGr3pYyxaPK9
lDIJP5i/4QijT8ueT0GFxZR5fTXL9Smyl1rsRTCDzbgNFYvjue1TikkFbuSDW3Tgm+dr1RDv5WNn
KMQAOLW8XOs2XFx1h+xy2gd3V1xS26cwmLF+2dzGI7yul1SK/5WJBCNyQ//jlSj//3HKgB2SdR3y
dGAWHLeuAun6bSZoqTXBEQ6a+MF3wZt63mSsVX9NgDhMZB5fVvGJT1yiS7VaYn96TA9+UmQ2Pvt9
cxuRUibM4u4vlLWCV8BpQq4BvsAI+vxyeNKXixK7yBnr/ERmxYmDvaZPtC3SdP+MPVmnzzg0BGsI
qkOw9FtY7AUJgGRtqIzhOh7X/rsIkdpaXQj9oPsqsyYhLceJl/HvbYR3lU3AwlcyKZSshSMmoson
lY73lQ3qv7rVamOVGqrNb5Q+9M9mKylF8SdRxKva1OOL7M7pv93nTiUuIsZX2lgvPB4NjNG20RLx
vd8g1x3PEIQukn73V/Vt24ox6Zd279GD2jzmQ3E7kpYj6eOMbae2tTQTMJ3IH7oSJqCDAPeLQ5Af
ZDfSevnBrMSb0i4ynmPXQQ2+sLFN+3lxGbe8mM5s1SS2xWJ1UQtJATRQuh8hdZvFw/Tdt8OhTJzu
mm8PSMGtaSkQGhjCWOipfy1Ty9Vq4lBlNF5UVE/G7VS3hgPihPfhxn+l8QzFoghEhbd13R7VYALy
XBLAUqCLzohmCNn6C2HAbLKPRBaS0jKZiM1Go/D8+Q+emh2LqT4T/GVfZlCRR3QXKzsXPqCRG+/G
4kzj53cTlj2Jon8OpQzluxEXWGozO0Mp7OxX5dgbyK6wEfVP5cc2vrf709btGCYjhs22FsA8wA1C
eGGd1kGN36CFUPgr2YvV8bQSP0bhVls1f1yHB4I3Xir1EkMpvPSE/3Uj7YQaClHaicPKBNs/UV31
FqiZuL0dkTsKZOiV9+v+85DYyWqBz9eKvOeg59sXWFmMGxzzQWV1KarMZLZdE58M4CjMwWQmY65o
dISb3UfhuUKVX2bIvNpy9UvabzJnnBegnDo2GlUAcMzXocO46w7OB4PIbeYmUeeZf3gurtT3H0vD
RvUwTvZgTREBLhbIBrs4JowLVzxPgl0grB7s/FgHUMPmEzFMFCU20W787Z341s9PdU/AvuK++82p
Q+KhAyTWzgs3cY20jvweHMlXKYeoXG/AOTHyJx020Mt+SSYyD1vSO7Em7HW4ktqHlSvC+KmsHD5Q
yY47MYbnnKiVq1jrGRXHqlY8snYdJ0YK57A4l+ghBum2gMwnjwsLQs7iZaBqu5n6omacOD0exT6n
LxiBFaxBwX9lQXdBM1Hta5wZVm6FmVAmHPUeso47MXhse6xvECncepvNotU4n6Jv6lXrQ5g4wMBU
bQ3vXAmmagUcToEhmS3OFWmCgJ7WLB+iqiAw8bnnY5GGfs6sW6029kXPLfg97AwLwW6vJhZJnKtp
x6Y6jVwyZSOM/2BWYQgglvSTry6Uh/d2c0YXU1idGxcpsmyHqA5zO3d9nc3/OQRMmvVHZWH3UZVN
bPWgpf2RccLSRL+8h0WxDwdYmjf1cFVaxl3fjG1XaF3b9lT2RbJFxJeCYYwO9A5ZCeck4kxLG8g5
iVKwjiZUtDWw2m6MTjYfof0sbQDfAYS8olpr8n35YEcQ5hsBLKPyYV+H+SeqTpWlD7WPPicvRI/2
dNEPlUYlip9YxQklPw7ACbXKElwcowY2fYfXHj6ivsZt/cD79uxIWZaRpZYGIVXrGB9WEI/pquEl
U5KSeLmtqs2lKQj8Gu7ptJS31mhkazfxDupoGzl9NWKApeF4wzxxRay2mP86mAEjyPmUP2llgz9A
ayypiIf2MLTvV226rmmx9hTYlhI+69xcTzGLNUX7hwstCED4v4eaMpzbKZ6gQMixVhLAPHNtGswt
pXJKDhpKXbaW7+iOtCPCfnG3t3wnm16A+hUo9EwrWmdVhZZIENrqhKDoZz3rGffCPJnrx2LW/b8k
P5mOJf/Ja6DfN7yeldh3HotvAPi08U2Nwpc1HPtZIX9JAZBH/h0C5/4Ej4nOD4pVPJRYeE8PEGvu
pj/iYet5+EuCAoDwWrj6ubFceocgFuB/WGsVXIhUZQRT+BtISzMsWu6s/CarOhqs80zvw+cYi9YQ
TbsGQH5n+JJyWZc0Y6AhWnG9v/D+aKpHhCmscDzVqWnfhWjlOCVWrL18KGH6lXB7zGI07YN03FNn
glfr06a1+n2A2ifQcMhfegrrwy0rz7fx7F4SbQVJApX9jQlv4d7CMGLNrS9lgZjurRMmYyRE3N8J
rOJDyHTeskgkiw+4Pj3eZ81/OYq9CE7N/W6Ynl6Fp/n+sCoZww6CUaC+bAQIaF3SrmQ29A4fQejG
gR9QQslWIwHG9dhl9G22nGsRbRC4JNZwhF9lgDu24vS1wOhej2A23JF6Hsm95O8HfJpy40j8z5K2
3YJ5i2VH3nnQydJ7kM1/+S8Pb3TVzyw1PkypzSy28AkovB9t52hP+72Es8PrvqRt8+IWeH0Sfygq
1Sdd9GZKWZjVIl3bB9GMILHLq/j6diVbruNfVwLx33hY5JWWNxPP+ZdqEwfAlICyV6sqFIR5GMru
uBaD/43QHc8R7qPPTEOKgQniXO83Y/XsUSlCeCBFX3CdVrGqwELKVLdBJJAaqVVfjhavdY+H0vf3
eqDjmNAyFxzeo2sQ8/GIZ+bIKymBI95xY74UHOdNhCxT7fzZG+Cxg4+CJqLtg/3Z5Faq70a/vTYK
ypGpbfG78XKADHeOSvukbSWlkL3PUZ7nOrQPDHl18yxJVhDTlv/KLFDpTD1d3CnHlkXERIwnjehV
6Tti2sevYhpGB0i+XXMj1YQ2SBfJl1Qg/3cWSTROKqQ0t7A0gUeAq6z7fyF+UPrEQ928fBwF7qMi
J7SiLoM9vnpJiEJSwB/nNWsCjJTdgFb9vYNCopiY/0pMiLZdjtkm+qfp17jsCM7N53iFZAhLyqer
hz1EPMX1S+fz1YCnBoAnzA7kigPziLbh9qQXsWj8lscnNazpgGT4NK7fo1U66mRPz+hejqWLs461
Mu9DFJnY8EZ1A/lBJudA66wDWd4zBqXHx8D6MBfya926MHR0MIv/5qQ8VwaruLfaeZ27TdSrFBTH
EXUQUN324U0++OqhD4dExh9kAsXRwmbS+pVap5zmLpJ7NvWWD+gvOTn5e/Eyc4LIEQ8F5hDmYg2B
hDUYDR2mBNzBGf9qvukDqm5X4jrfuPvTWnkghIaT9j0NN/fTuhyC2eOA9qCcfUBfKM7hTZckRBb2
5mjgRBVnh4wPrnIJH/PabXIE+NR9O/DuikOXf8vuIidRPwkJzkwppDegwM87ODzM9AWdmI2MN4D2
AoT0Dg45tAN1FEUV3SvGHlm3FS2776cY6BWugjuGypCI7AJ6Coh4WyX1q+Lh1QDkOWf4hH9RbNz7
gzaCkaoYSVFZp3RVzGIGTG4/FmGZgLS5amWdKCU4gvZa6S3qSa0yozrM9AflYr0/3iX10ztDwInO
8V59D0ADPbjjdL+VPKLW5M7wSjX8qyE9UDaq0IHXIaZrtDNbcNiuPbCEt5qrkYmq7/NEMoJYXIoS
qa7/kwNxnjEq66g4KgWID8JC2tzxG3UZx8juxjXe39qSG9mWDy66m05BFPm+FguqTxS+3XDFRWj5
j+bEdweT6IrsjIVgQye92RRY4ZGG3cVDsvE66JU1cS4CzLLJh8/uBzpH2f6QDdLrunblt666TYQ9
KCWcfnf9bNaHb7Fd96x78W80ReTJXham+iN+gNm0jI0+QK/izRokCaU3rJtN0Hq1YvkOH4MrkW8w
rmPVNMAk3KizBA8AkqmHggUXeGqVeeAC1G6KIAeEL2oS9U9ahTEAEN9X1WssbeF9Lgmf6hVszX02
o07gemBVaMaBMhV3c8z9Cbj38HNFy3HgmNocTVTzEB37BSUXVaeq92QHrfhh1szZCBKuzO7tcn8o
LpWJG1/RFfZla1UTw2KL0CGPy9MCvcS2aeGt9rdoh/+jR8+e4BJKOL1TgeEtkCuwevJuNRrAm2Oa
gPB1lopjnCOvw+iqLD/EIGn2HVfwzTrjLcs7Nz+5Tzyk79qRXW8yMHLO+lOeoy2ItC89lUhKMIEO
g+wTN4kRJsfjMBRINDKW0B/TNplBO7SyeSIGrsL4plSBVT5Tc89KNYrW3tSfOg+gO9YdqG9bogft
Vf0xx5jR70dKduAqmezZHxYz9obJ4IWVmetUUIqTfFwVDWuLDmx4EXDRxCnm/YmffiK+HYVTJ8bn
x2LHlztP7arJ8ecMkb1DPaDXreJt4qYwDsBlnUHkeHHQRayHQFPK4gln8u0aLAXjdsitDPku9q2j
4V8ZWB4I7ESnK+P4KbBfBw1EKQs5d/bGrZMfjBSmMZuTDhBN8Q6i3NifS8e1PdGAHOg2E7cE2XJc
ePDQY3i/9RAR/tDnj3z+xGPV7uZz+L8wTdWmleCkSUdfZh9THG+cR+wpV1wzLPOvHIAGUGVI9rmC
umF9XPgEBgKq9gHSrT4sGrs5r6WaPeCqDkiMO7FdGLdJgkLyYIsc+lBYQNwdTuiaCMMsh96+pPRt
AuLxCj5FjUBV4FPyPNLXCnMKWiti+XVfrqRj+QAFzjDZPWGExcyykz7WmyM4lVQt66VUuMpcI6oP
D01rHSXMTzUJyewI2hzdebg9hoelepdaEZ29lK7Y4xEOTMoxXQMq41HODYEbbC9PrkoyLb/wAFkm
eSGta+LA8SDCXgT4Npt3vY9XVcRnJFnRt5WeTLKlvbVf9cpX5WHknyj7sXPZkWf+5g9vomsU8zJ5
hAkJSPKEJGa5GZCo6MWMm+ugDA753C34efHzxXGb5shC3NBdvxkPTRZ/jjkIEIQ88fu76hZtOrDi
Sp/bzpZI/wqJME7S3/hM7qxwLdx61yJPRf+PtZOPqjs+8eydMkeLk3/Hnu3QqWuSy5nNrZfKhgm3
Bu/EMJ2uYBqIdrWOTz7lBGibCNOSwlp+7dYQRWF2WB9aFpt8n8Z2lz4JLBLlIxmrPh3BnEleRHLx
18NK7TL4d4HD+3NMO+1zbw7eXlTGA8BuItm9hg5wfCcEXqkkvPj3oi8JeSlNd+/VfNwcK/SZaGRd
z7XvCGW1Ysto6mJsA0QpJ9OoYVso1Lhnvm6dF5a297JkgYipI3lgxrPkoRq6kndf+zU87PQquUaZ
+QsAXUoWc45FbETBpn6IV8K2gj+q7HwViH0h6NjS1KWYRRZQWBewdeh/op/brb6yqpjyBwBsPWNl
8D08UkxpihvFFrnrDyD/tYWeF3Ad8z4ju1fcJAArXeVvB++KSVlE9MwKNSjFpu8rRlPXArPfvu1M
S6KduQ2ncCzGVKt3pH38w5IUSubBlzLyw4Q+9Cn3ZW/evfppc1DGKjcft7Z4Si4j7k12cZKH3AfD
vFZCMsR4l59Rj5rBRh6ZZSh7luVHsvKmvB0BNq7fkMLqFt5NPhx4+qWo7+acAnXFmoR+beRdwUai
gCAYT8NRzgv/MYUYMCys6CTKksxKK1vHvF3EepxOPONf7M6qNvDI1zOQJILuD8NNWbMVj1ukt/jv
XdB2XjsvFz7qxXfGx5xL0ZsE4zdizB8dnLnjcxORDpGUWqaU4xASVQhp/abrkuVHF2CC7tbdLXgY
uK9zoZH29nHnH/AJXvykbZATxu1xOetMlKm0aybaESkySiFbllDKUpn9pbirAcjvB1oAgz7lNghX
jJ7UaPyFOBImVcDath341g4DqKePmGnBAmiZveIXzNCMs7nu8RUKap1FnImEpGiaAkzPE+Rz995i
S8s9qSVOHFkCq4iGXVh1B1ulvkSdPT0KWaVS4roJiEidWMlunp3OTdf/L0Ns2WiUCzbAvzQgDKA3
Xb+FSzwexO745AWZRl4A8oiM0jUQFeoYR1xrtl3eLm5ND/MzDJxMFtUK88HC2iptiF5yP5qPu4Zv
SwJUVx5QAl4jOgyDkxjb5+LjFViGNhgk1gLQqCyrRViWO/bbq/e4ov55yYp+9FgrbhZIB/R4wLAB
UdQsbhiaQNpcbi9iKozQMrzgOi5u0OnTWleHsMicix33Dodv3p4zPFdf4urQymP69O6SlUnv9cxu
JNy15rCIWfjiKkX2aUfH4fm1XdGyp62pL72sE2yF39NOsAS3G5FLV/T8WLEW0Vbhu0nuj0LxAi0e
EwJygpLZzPWFKV2BT9I2nhC4WvPQ8zVzyIDVww0AAaw1MG6UH5m++zqGTjEFfO9sWMzlpFGwR2z/
8spxTLqtw981t6VMvLH6j0TJ19BIyaGJlEHuk1AsnwFh/OQdUYVfK+FWzQ169EgPY8iJEpACQCG+
YHMaOyHr6qsPlvrDnqppT3qVa3BChQmjGZBQyd96afUxbTRc4rm/Idvr6AHyy0m9Voh9iXlLbkKv
AHi201yPAUwcKVOorp0CuuzFbosyoeB5uAZTA15QSwWBxh+1cM6TWrzx6eDhzmYPonBFAKrVifSy
KmufE9UWVHPL0dU/KJu0PgYtfSSetYXWyVR4kE3l6xmP0TX232zaEncpJPlqevs6LeGcHeynT4yj
IouRUm+Q6cekbtXxAZ+wsCTocN4xGy//1l3Hb/E/8R92dVHBYanbed26MdHSfvUfeMwMnvOPhjCo
jqrYuiVQauAwanKynSvP+LSdtzTV9OA8sc/G77x4X3CJNymNEpw6JpegNDWsXz3wJ2CXNYXxzn58
OAqsb8yJZ5CwxBu2uDp5LKoLhxY5pa/w75CzO/upJcCvI49cl9y8MVvtgFQFcfX23V05y7VJ5eDa
wWWAxx2rkkaxPE0lKLOGjy0UY7rNYbO/8JwtdWZbXjzj42+YK53xHvwf2HRty8OrMOFgBp2Y/gmd
zQgYJrL8uoLSZjryp8T+0qKN9uEc0LX3Xmv35nJ5ya/L6CbmbU3/K9t8+IXcc7/0eDg3G+/BicDn
vdfnk+uyArfYWaQ5NnROd3bhEy3xYt/U0zpaVvx+c8kobGbWq5MMQsYjvLuNsHbaoZXRY3n0v2oI
0c6uwbkf34Tt0GA+R5Bq/lMRrEzM1kF2paj0HIbOdWIOInaXOzTnkXl1c9EzmMtOcqPZBIVIzYwC
GTkrx+8060p8l3Y4vAekVE2wcTCln41EJY2tKiP/OXw+51EwiVsdGvhtO5XzEmK8glZcUpKxJjyY
CCf6bvBfVWE5XB7GnDPbOJUARw85yklUEqKd7rhoYyoQDjsOQBEsZgTOMLBn9E5Mjyxk1Bpt9IVz
zU5YAJ/fBRyLiyND1NTM+mfCkP3+wZzFcIiq8Ifu7cYKy/AwmnI9VSfbECq/uGKpxBlvgJoV5EHL
ihgNmd2xjHIAcNl6iQfIr37Q9gam5M5FacaSI9byphHmRYBlx6EqWC1F89tWcjvr305KJzsvw7Ko
5LtVtkbGbX2Fw0x8I9ZRJDwZ1sc4ynhiu0RZrV0zMMMgT7OV0m0OBXBgNhA5Ahg11wStwRE/SM3I
VLhaI5K7WTruLQPtJrWM/c61uGYOkjrz5uDatk4d8dhEoOc39lQNjuMQRIBrA0CUmofTMT/osaaq
iSTlYiy3NVl0cIxSPrrV1bU1YjDc36W0vji8FDHvAcumijhYB+VlAqs6LWL5exzcDNqRZ/1TqKpx
ASc6mrlHHwKg1eNTnM+yxiHzdgeywxq/iauUV+82KvIvVd4ITfAERomC2ac0Cj/eAU/I8S3GFqzc
xw9UX0d+Z/UfFZFHYFEMT4tE4/PIh1K1QMrzdzO9btUaoJpFITh09td7I9gib2ELRTd4UDZKIgL5
ijMFtnPKkwnnT/fxMYzpi7k9+awpYfNpNHa3l743bR1VhQJMA+EK1Uc78jG3W60az9fefIGQQhj8
CDUVtLwvxlUY6JmI2OC/97JInqAtGcAxB41DASW5SwHKIKcBl7DCzIvGKXKPDSWGcbsP0/u4RlQt
4a8CshInrO9WrCWLtAGMYLNaEGmQ3i+Uhw/a/cnlB9LZJbCTA/3zmA3QkdHiHDG5ZNiAar9RO5+M
Su4KfIXhZL9V67HJkTKesSCYPNzK//1oZ9t7DqZVG13t2Ww+WsjFLe/6CLOLrN+A7nZMSYaS7xUj
0MKWUdUD2Kua/5Ip740rN8K8TXXD0/Ed92FTnzP2J2Qb0QxWzG4gizo1+5GATnyQbA7J6nib0ri/
Z5G4oce5eBnARbV++SClO48cvnX8VDSpYOm7TZuvOuv7K38lIf130MsDInhsxWKV3wrj+okb714r
qRyBPj/2VvSLZ7Uxsd0W/+kvfEIBUoL2dwDUd+AXoiwAodDPnKRo4Z12F5MYcyrEcH3SeunWJfkC
c4lPPuSdC1Pm99DEuhJoWE4i+cx426QsS0vwCCTr2I9uEDp298VMEYslfeLRVYNRlG1/0qbPfe4t
LfCyerdJ8RNAoRpbhv1Up2/hZY5JDa4PHSIin+5kVGZ4G2gx4KHGNfEjWxFrEeQzV7FD6ZQFOPgz
jmDVg2i546JDppzZqSMte+M7IyYvRUUlgqQX+8IP1g6/rSdernz1HZDFkVR+rx/syJ7R5JgJu4br
rN+IRn00wx/MCJHEY7R+GprhJArdQmZVKwqkBlPWuju5RhLfIyJ9btCIzjLeJ4kP5/XQxOmmlmRf
RJ8DYSXjndzveUiWOTI0PvV919HfXQ05XP1Z750iMnEnyvIiP0JQQo2yk0FlxCuST6+IdXP4UQKo
ZElcymgEs2EcrY3n/zUg2zIuNp//GVysDvhXJf0+hsEcL93E1ludr6QDEoyxbZBiRzu8ucCKVjns
GPakEm5OzBtFieTTwC1MvPlbq2blDX++uiW8u3kSuiSVBBm7YEHD3/ccO9ZIcxnKlFoNvocB8PSQ
Dd0G0l+QA0ZL2KKCG34+GYEOW4PtVlK697xykaLiK/1zKeJRvtGv5EOQrX25OOezhVR2P/Tdw9Cb
aanYgV3xi4v9AO94shIu0VHNG+M6c3/kYLLPUDcQY2uOLQwpOXTSJ92W8awFEHAqQlZ7RsoG+w9h
VV6X3/cs0lILuh9uUGfXVwWTpDn+CLyuPPDBAvMaMy3ZNqZbb5mJ/FawQ9hkTgCVh60ebCdn1VfT
O8GXzh0i174Kq0mM/BIOMz9M1qxcz3LR5QF5soPirI50AUqlts4aGJUrrerRA5ZiWy4jFd+J33w5
0TZbd2KE1+HOy93EmTe+BbjBwbu4oCoHah/RmUukC/4CwCYBc/nTTzeRL2ImHPLLyd02ZIVIxojN
Ml1u/Y9oSPV+bsSHldpzsZf0+7BabAmd7ORFfotgfgL0HEmLJpHZMX/cGnpvobfEK1k2MxF8D7Wv
mNhSw0/vg9RWLi0ZRJfXF4zI7nMuzmKW2uCOXOFu9PeFhJknAPyaaK8pJmJvnUoJEKZUXtl1tIuS
aceCX5x1LtmnsVvCwL3XDleINrOyKT5DuMSGgq+zB+PV+i31Zz91vpRVT4q0QSaBf924Guynyinj
HZU4gQjWzoVpJQKOjWFIf94TQ4pgDhiE9Juwfit/rlswsqLCS/wz7zq3lWmfc1DKaUTaxijnIn0i
a74+Rl+N8FrQMZAvouLPaURacbhYdcmGgwJbpFhisr5E8QA2rdje3AUIX5kimRr0FpNVcqZwfumY
OgM26PANXEM2kQ4Qvh1+rsT5IdOCBVxlRpxnTzUAhIhwXmCdRvQtS+qJ843HR/vMSTEAiTRTUiIj
6Mb30QGic2qlFA53TE7mgW1JhRqkFkJAc4Eeg8zSnfkptv1VF1rCNS1ZofVBhT6hPsIRx8LqL+g+
6fbY56eHXQL7LjmlefCgCTzDb49NKsORbH7zUvTgRoBq7jAStTBLUJvhHu90suOzpXb/VIFvlU6s
oHrnVlSurvcRPFtKLV+rfsPtXuLVo6Rb+CAvhz19zX8yhfciGhfxHoNcUHpVQOoUI7xfSetAIrcw
OaWyMMaR4LCZx1FMwPYIT/o0G+FadSZTOcnwHi3B24+fTVM4VQJ8DQdSCJdBS8gKd/Sac20PP/Yz
pykzMl5fiqz3TeBRzgrptqg3xrLLJkKpEnPWn5JIFrdsZ7moN5dXI5Vy2RaoyNGtFHScLMeIgUHa
Cb2gmF6nx/dlWjgmIudNYDcmMJM/vLZ8bsGJ1O/10TGIaePUbLOj0qUzYzUMsdeMx5xT7vf7Cl5J
1y9Ub5AZ1+W3t8ypPglY07j2Hv+smI6TJcBumdWoGJb1FCc6JICuAkAGQcnHAT4XmiDK9WRC+Tuq
drbPhLnZcsZDrMuaktXMGOebYnfi6i7PXSZ4Xvjd1SIHkvaw3Oxru23jL/evpDWWoi0O/l47LnZT
LE43JQ5p34I7AhU4wQV42w2CpEfq9Ycz2otLQ0+G/0/vbPpMmKRUwA0ArxbA+BDvkZ/VFZG1tpPI
SYUsVTBawdrwmaiBqibn+/HoTfKjwDY17Kevj+RY/Vd7+Cxr/4Bsl3QLPjQyZ0armJV0TPNskQjs
rUSLIMtTNyDmJb91rxukIEYWSQ1BbaxVyjU8MfEeUJS+WjVQvahA5AZsRBoJn7kGX2zDjAQdy+zf
WzSywjSpEnd3vSZQ+AErNPzdS/I2jr5+IPArSbD+Gb7U3LQJ8nZAVP59utLEcH258EIGVipYRG4K
0xdmk99KJb1RSlxH4DfvoffdAQbGjsU8r7CiBwHHBO8BpvyGclsx3Cbtk+PqdQ9SwX4Xz3uYXshz
tLMjwpwcWPBOIRc1u1112Cj91tLkMc2QN/z372PpHZ5AVaKeb7lpZf2R42drUvXDH4jSEbQ6OOUL
gPJXGpUnIfuu++ZQdjsrjt5GLEvrtQ2xBWJLIIVSCSeX/MzuBFH6R/aH8oTuVM3pCXWtHd8eCMFQ
JoKwMQMYwdKiwdWVvDTAvmpzOoo3S2hDNWlBeuaLvRwWIdmYKObocCGJv0FniRI4JuQea+CEn12s
B9oadEp+/QVWvEzEAWuS2pOpkSI/vagMyLGeFR5yS89+0XcckLJvzrfEvpvMEvVx2oWsqezHUYXp
NXqsc1OKGXfcsx1l50PgxjO9f+LxrlJ6Q91v3F/fFa8H/FHvLXLuDZfMFs9jH9Z8N1x3CyvEATzi
1RCKpANfZZP8K+CWbRX4tCRfnhTANI74QlRBBJwi5b5zc3rI5bfcDQ0dP2GBALPKbXYOfbZuGONb
qdxwdFgoAS0E4gk/G3lOArGGKwMVPFfTR91bhgDcC/Rqoni65wXtYzQyHoiXGVDZV5+tjza2t8wl
62xKyeBfq+jxH1ggi5Te0BNf41AADPs4iYXiUhJvn25Uj5+X8/PWw2nusfXW4kUgc05yxiHOajr+
N2Nkhab+EB2rBO+TBXyehNAr4KNux7tTtg0+wdjblF/ADoan++iza9DHMJF3gBbTDEVhJtK6AFgy
jEeInqLevgBDv75iSFDepBwMA0uezwQRQRqzhFXZ4eWNNs+F9T2FfnoYfYUK2h9LSCoqClNU074s
bWG8gFR5E1gyHgXLtK04rnNxzs0k8BgCQf0LbX+2V2OkBGQVcq6230WxGIS7sPCzeoke5W41GppW
aMIZyUmwP8Dlp6LxzkRkoBl6Hr3oPFjIJ3sYGpqJkvQusEiHJ8tbDWQ1UcqcwL8Alx6hsDwPYV0g
fMuOQ2Z1MNW/RmFOopAHAm4gh0Og1E4c5bByjJm+zcfOrlzH9tz+7v1eKrwx81Rtvf+0/HSfnOzx
gr82dPUnFrNx4qHMgrkLNIDsc/5UpMAsZuP0OrKC+5mS5uaJaEDlTyCcu8jBf4tSj0uozGVuTFJH
61QmRMoHjpHwBagXW8lVIULFdcY2wCLF1v5FsLMpWEWRDCG+sQrkC+6n3QE059WQOS6N2PGTDJXo
+JITsrxziBLcWCC7+rVC2mPriILrwJQTMl98gC20nRI24Qvth6L82G2AzmLmHypoIIpKXIyo7ePg
j9xz1bdsGQdb/t+AMUGRkhN3/4YIrKGAMYDrrrcMqIEb1opHzVwtO1Pod3v04GVTWtD/i3L4fNFS
aNApz2UPw75H+1ntNxJ4QwTYsMuJAxcIEjY3ZIv0sIWKSq5KI1us17BrOYwrGCw2Xboqtd2PVG0A
TH2QsXKivbEU3cBjdOrBQoscm1ZsSuy0XT9DUydRPPj670yFjyLQqi41hqsbgXBUNpWVTl3TMZiG
qKNhUwR4XHr1hMZ+7qwTQxRAhYZgOLCriAmne/f2+IcvuYQDj36oBIOOyajR0Q8Mx8Bd7wnvcWwj
UIo44yE++uzQ4hRZjMjgR14w5eGBMWyj+m8kMgrjRiOikEuhFGM5NeeGtd/lZ2CjGILGHeOe1sH1
s6ICaRFn2mGV+K3eC2g1tAEKX8GZ7MNJYPbYTirG8N+Yv9GvMxFfQ1fftC3ulyBElD19jevYCDZb
Pif0t8+zME+8N2YqgEenL1a7NVPz87H0TDtj+7Pgrkj90zLBsaIBAaeU0OD8GFoQYzlRavySFcm7
YwbxEgaPUVhvNEOTYprxwEJLzoti9obgeVAalQs9+Q4UAfEacVfkohugicTTRD7lHnJ9P526IEIp
nmjW/oO2vTo+rm3yhtvI+22MANIIlXFjgPkdQSEx4suzcJ/ePJ/XLNnujgNc8Q1JFjvLImccvxOF
1C2Ligjl8s7fdawrwO8pi9KDJVmfFPHrpdn23OCVtL9UHPzYRVRHhi2CsfiSJOCRj2TTrD+x9o+V
A+q6Du7WhSZu3g+R3XJ466bhUUsaLKu3oySUuJYVqsutMk9hO9gH3a4I7x0JlO7IqUalTVCaJAMi
Af98QGB2TJJBl6gQ58W+NoOmhK+po/GgI0I7Qmczs+7Ytp2PCDlRhB4Q2U4c7rwNp3CVWsogOZT+
0KCrLk41zqmQFDdiMx6ZzMpqnQvtJVheouCceURQWgIBa586KCKO7pxZB+bjhT0yTFbhwXEfGqJ6
81hDFjS/kolZwEhNX6Yg4COQIMbh36RIRhW4qEraPlKaZNCOTIQMxQlBwYCIfqY8FmmafYhlZqek
OODIMAl6/8+OfqkpEItUDtUgg/WvQ79DlJ1rUC2MPvEdMWXEiHg6PoY9+KI8VajeGgaTyrQ9OY8X
XHL+u8dAHlN9XOrf0Edb1q+hu/RJD6MmWbdiJiVLYNCgNaQf8G8S+329ppQltE9RNPuK415gfrpS
O/fnF1FtZViuNOHGHQV3dfiHDYZFVWxBhoUqOsv2+IwDbDlB7MrBuI8CTsG20RF5s0nDWNCw+WU8
5Dc8ToQoThDu2UNQIvC8ENiuA6xkiNL8Pm3yI5biD+6AbwTfILCFe6motGTDvtS1cf44ci64Y4NM
5cZmc3pxK3UAMwno/B9tE/Pz/mXZX8iIGatMUePnXtNVRwPicnP9JTsEaDWum21gY7lLcmRe77ZW
9i1DEcmWcZflfd3EO8pZo9tbzgtdpvbCqycHhtNBf3w0dGstX5tAIrosm/mbcAx/IglskfJ0W3He
sP4Z5GO75/OxUUIlVT5oyeYyPYecnTSR5GmmZmMnOqhxSCYIeZZczuZ6ySTvOwiB1YfTu+GfP4Xn
Q21nqyf+vUAs2VAcLIqBjD+f8V1b1FaF++37nQPSuK1EfSTu/DWtjAce+aNZxIFkWzHf1UPCtI5Z
KAl+NLCCKrn0p3iUAYxFMFSVj6QCfmqwnZ94QRgtczbKOQNMpdMt//ErNuaAmMbyl7PDQA0o40V8
aUXv+3ElEqY7c/DfgAKskrztDsSDs/oZDx+h+uJrmKnkAZbOBirOoxHZz8h5YMx2O0RsIfmLKu1T
J3p5E2bPvalem+t90tGPVlUxKteoytXkXJVfom83hMpwCdxXYrSNLSqAbO5Vxuwuz+3Scbss39tj
ktnCSClcERdOs4mtF3D4ZXsESqwCxdk3kFo2aQIdI77s5j5lOno97OTDHnksXwGxzPAR8YiESUXP
8dasms4O/lRueMuduNdadrl3edgIoF2YhLLphqck9N4v5/+4o/Lj5DP4opJz2X78IC6a7f7QOUCo
LmGQz4dkbPbhlo3lvNfLu1goItQz23oaW8gPhxcit2swYNRtVry+rZkpfn0e2MnfXu1PU6a3stoV
Tvy25oiXK+N+rxFPIcM+BYreaCrtRAxUmy/XqUzk6tsmE0gQ7nwg3Sp2fELxX4/6sW1pdWiFokI5
X+WLlIoUh7sZfirnDKLli6VHlyJKRskay+pGMnNaY78se8Z+93O5bBtdv/JWVLI7a9CStcqa9xsj
gjeowOLjXNqLCd1BUXmdgjmzaD2y/6v+jd46REnH8ptMqddfAtTiSVtm+o5bPIsjrN5LuLj+NUMx
J8ctOehsD8ys0jH+Pe0OiWuPY3ioz2yY7PeMIVRBNZGQvwETOea5WZMZnZXzpAh/crI51PnyIRm8
OYxRixfFlIwC0HaNIEo+x6bYC/ls53Km+dq1IRQGLQGYLk7uadMZvxveyxJDdutAwrs8YGyafWkp
Ug5XRzuh+yPjQ/BzexW/vDPkAIEKAqUxOQfNVS/9VAPGDDig2jKmu6LBcnVuv7fYmNHZLffhfwNJ
Yjg0g+JTbtthRAZBps70k55qaSsP2+TvdSN+42QmnN7n6OXNLDXAF4+KcZhYjVa+7Q8qFrXZg792
o5TOIAnDlhNLzw0UnzCraKxTG8aLn49NXfJFisTcY6aPpvMuwu8dmzSUHm/BmxJzOC+0q273iCIV
CKVLQf8wTmGkpByRAz1Yn661bOpGCiFerWqas4I0M0la7u559kHichoU2Zp/gooYqGagz7lg3bCw
Q4J+y/THTylF+9Yz6w/THo1qVYP72pX1+Qsz9ukRiFd2lX7JEH4EekUNagZ177WPkZlsjShxV0Gi
zw2+99BpnvyBKrn0cyNlsROBgvHP7WLtHeF/XejjqbMmUUUOC4j24p43qlLAVO1/pAEC4JvhjXKM
+RtIYEuX4nn2pbfRimh0BPOxlDSCzY8gBZS29PVHqIdSZkpG1p5zKp91bxQugkoo2F7NXJh8Zttw
w2cyPezDGb0YEU5m3hLpWZOhpIx/aODURmyb4qTqZBrDpcWT+yhs68ufojf/FHY1kD2mdE7VF4IF
h/dvbhLu45EMu1T2E/9FO4xwNET8NlKIg7N9sChlYcskLiRgw4tNLsTT5NJS+9oSekVfjc2KDR+z
Xhb74Y1IqZN1Rh8CtcQFBcNoHo6389IM5VqAkqeXu79zqVDwffQOobYB18tFJ3zJwxTJfa5rp2wM
3tofwRx9QMB5UrF7SbchBygeVxT3HBftjbyIbZTshtv79a5xJTKYTuOcsGcB5VH1C2gdvmj0pNek
OnbsebSmnbizYDisYq+lHA8ieExuYliRD6zUbRDiVkeaZXs+WHWXS6JJwJU5vXKvaSZzRrlwuEYd
wL1BMPwnBBnJS1yityBHN9NwiwF8MOKv7/SPchwnfDTL/d5TSuETrSK/maqQNtz3DJ3jAk46qKYe
+VhFV+yuIV4AqeYUjEH1hKov6xLLUVgB4IuORpZhmP3q8dCATUA3RglC7NJrZu0PlE3ghzKiUz6H
BkCOk+gkhW0UKBAJTroa9C/p0+jcnpt190icUmQmIvuyavKlJLnisYBOZf2kvbDvMUPEqslUtcG0
vGwfs/frPW4Tx8ePGqc5DqPIPtzyQqFZS30GO5U50i4xyQCICxj9VqWQYBPtZjaOmfBtYBXTQK6w
VAog2I1jjriDM6isP+tdhB7pQGiTJNvQqCTCKf13N5kP0fEGKsfVwtdohQ4sGl9gh2kAvAWp1nqg
18KJjhM51hYjONWgUq9aSem1ISCTUfBlrPnFj3OHYiuO4e6zCSETW1S/hvAm15sRGwl89NacQcjw
FmEZ26TcoFOKRZ1YqjWYRtZkT6B8UywSaQt6QDbWkO0DKg7MikPavVYw8ryrkZpUy/yUFNO2PAUS
NfQNVoacqEBA6QHfGB1HiBGnRCKW/In4LAwyVC5PblxRzQ2hBIq+6h4Fen05CngCiurrazJ9/Zrt
zeNFVJXG9lfYQjjcUqFtBj1xFQB4rAmC81wk1Recf2d1/CSZCUzCSEJdTinBUAQ/JBwDUrlvtOzR
65JPdw/ya33T6YyyI93t0zebkwyasagPxszHiWo8snAlAYSNlo6mws+49KCgC1vM4CBNc0oreNMs
tiOG5rcPzabwnnvJc21NE2C5MXLMRrn9g19/vVM2iFsxvKtTFA0eq7emkX7LF0666O1hPGDdcsz9
D51rL4f2m1mhcy+bjEBNCMstr0MH/9s/sG0cRm9YqX9hvFQolTz/Bd0HXtzZJrDVWAwls/g/bFXo
2hsJBwLxlg3XK9j7i6tiE+JQUgVmaUce62bNBB6iaNIbOdUDN9wgg9MGTzY5QRy6qhNlLvsFBa2n
7M1WaEyh5kxMobAZpWRNhYzpopI1xfE2NWKPy9uQeyD8lZvMriXhHCtGfiin4l8C5jhzxvh6CfR4
wYTy+1ranglrg7NsjDizPkXIYiNgWnvO/VTJR5S9l9CoxqAstX77exe5AO29SOWIY/VyHlhDc3R5
g75/O6T28IzjxwmOL561drZb5R4NIjlSC/OZGpytcp5Y3uTGMiFq4bsP5cx7sozb6kb0tKSIy4b/
XuQ9ZREnMDg+BQQMb2rc+hsYP79ol9vB+Jc3w4XGL/I8hTp9ZOPkKIOxsqN7dWVQjfYxr+A/60f/
EAPSoWLeMTG8675nrKek9XIw5Cepe/o0QpzGQWoRleEYx0DM2fs5OY0eXoJuxLqXK7wY+lrHmloP
d/S5hs1Z2a36R/6fhg96ship1pyCqxKNZPK893OxRLo8nA9xtCRmlSBWwBxmF4zwlLIVRuKvMFn4
D9YQXAA+1aki1OYct87i9Iy0XfYivQlmQprrckFnarTzdGUohoZydoKRw2iK9cCKtudTEng4usuo
hg0ciiFmS5qZBNlOnzuX7SVqren+emd+j6AvpBiOMbivYVVG+u4WFKnKHzImw4fExabsTmxdirII
ryqh9eqrDxAT7UoE8odi8exJ+hpaMtnuqeQiWS6fkX0TeM7P/6D9DxVhxGsoewzypTu6blg6NFjU
oWcJFTfo25JJWzUro4LQi8oFfVzaDyT85y9gWzda5kgtfImvTNYrPyptgpEa2DrwEmp9ky5ZqvlU
y7ydc0JzpuqyGPYADACWT9iUWVGkwRuEDq0bsvambzERfEOfdKNBy+zwA6sGD4tkmyD0akxI+0nV
Ehf0zJfHgdVAp8C39riQ4bAONyyE/svGMAxQfcyeBqMZiKKJsCrtGmMwkObnO9BbzqyckKsFKMdE
td5LVXBmErlPyP2XtCUdC5ov0W2z5chrojlv8UEGajUToEpVuuTlng9ia1vAShf2anGe1KayjcDx
DWP37g9XmgNn7c8pFxHNRZBsu+Rw/YVD+vHWoo7mZXKKCivufKki0NHjGVYiHKVxsOMj/+F8XK5+
laeTS+7hzZ+5WKc26yvzIT+SiiT+uLjWq7SUfFk0eUF+fzVsSO5KEK19Wy2ckfJn02uMKWrBUNg0
ON5fG9IDysCb2AAoyHt+t5U+Dr1UpCYURdsZq/E2dj0h6qz/EzMejLCAq/bEP3tY2WuN2QtwQn6/
l9MJLJeNgFXxToKN7w880zxpfunXiuIH/+K2L/tgHAAXtNNF3XFAijIVr1O68waD0YAPCaCt6NDP
kGMixbNuriEadJ7zYXIOC8spZCQTFWCQkdMdD3upMRnmOGPDGK6vMcm1oT+1LUGIWGjafjH8JAah
9f0I1CAIppMMppnvatNiS8QIWyZwk/lAA6O+vx7hMs33Wrcw3mZCtoErtdsubSmGVP2qvvw1hkaS
WdWQuoRIXZnn0hSC4FkqS6IVgSfi6YeHd+zp3W0q+MMZ03c40PQPoxjygq+HpT2HX05wZMUxZ6qN
FUmB4iK2g7agYBgXU211oWOo9I8XS6/UHpK/UYshcBnWchtNKyfj3r9MdPWuD00urjjmSx+MfJvJ
dk4u17X7k0UdQkoK8BUD3kCq9ggQ8TLhuOSacZfAyocSHv7+kQDeRpPTE3VwXO4GcJ98354NbIPl
ZS2xALx/UfLdYoDIU2gESCHllewdsIssW0I62EyRsQWpamVyEwFfXFL5GlsUYCwRGbH3oKVtBEBV
W3h2kFIvpnP9PdKjl+je3cljHyfm6ZRgn15EFfh/YD+5b+KqPjdfONjf07XMbiNd2UJ/8rjTCW3b
QLm3OEh3cJiBi3j8SZyC4sSYuI3xFq/Y1dRkPCIZppWmw9UsinQSkNnjSnB+GAKF4wZSMN5+Q0F5
pV+bVNPF8gLKw2I5vSQREyKd2Fn0WrsK92gyPmNpiLrXbvgSmrgK3W8riYIF6uO1ZFnVEI/TW/2o
2O8ZUuLL/o7ptObsClWekBGTBAnVpSj149Lyy7y3pm63DCvK2qTWL6Rh4/yiA04CZjsGEfspu874
dPGaDhga2pf+mQfUFEAWqCMYImSDJVAxMUjfmJ+mUEbnUz12t7dOLP265zsK+FE93S30xRf7P8tX
PoM8l5KHU+qYTfEqlPQK+Qjuc1Ff52Impfbjktfp65+KILZ1gIb0JgzK0DD2BwEhVZYBsW6Xplyk
ltpVM3Ce7UWSznj9G2XBI7aIl/xREgyhEDs7awcnQoP68q8J8SMn08cY9SYBMbcp8L79QzjHoeC2
Ku158zMj4Djh/Asy29vDfBbnONSWqWEAOX1LtAd36+YCH+ZNoMI4c6jrsdC2DaMkazNnCSzW2v8O
fda5nlMZiFKtVCNvaaa8Y/FlzzArMlByLjOyVwUy3gAc6Q26c/Je6WcCSJLKsfbe86oXb7widyik
n+ivSXie8/CtrDzlPUS8/y9lH0ykBK7r/O27pijfTDdlJ/sUk97ZQrmv+vTm9kx69LqrfZP0HTcw
UDYEEHqxM6xGr1LWXu1x63yn6Z8Yjf1a7tKebXZgVgdWJ6BMQHQ7Lv6VCuPgaDHxzgsxj3phzm2Y
U0HOIYUVgCC1n/N+4z+y9TvAaUwAf0TgPv9RYqII2xd4MHMQQLXadAhzhAOzHKj5dd0wuvGXzO7l
LTYI+8NKBUeeX+GjFys+INjRMfZso/mCCxoOmU5CC4OwWxaoOluO3AMbTA9rfW+oz+Gc37phgYIh
uFsvOdUZIHEkxC04uOgA9FmZOFQztiLrZ1aIhYaivgC+9jpNn9qwmCyv8ninpUTLwsAFYv/tU4JI
6nx6zKyI1rImikw4gFlF8lSZIDNDBx/78US5Aewt+JjTpMgaXx6efaWzhUWnI5KDCsJLBMJgHFtX
sgW/c0LfYfYhsfYuGUPRtcVtCH5b7CHMQJba4dY9kSrJIzd++FvjXVCaMPiOb0Webm9hVDqoM80O
jyDtqzpROoAQmK7yI7HVNG0cgHptROEiDuEe7RddyuTZqaEApn0p4p/Yu4ahozBOW9rk6F4eUBv+
USDp1WieL/PdPlBkROeSXYK3llE2aCr20uAsKxtLIiEk3ABkpsZaSlIJ/Rhw+lw7ljCr9XWXzbOd
PwOu/LuH44HUeXcgWm1HDH74xTGFhmh5YjWB1yiSyD6KbVD2vWmrY6zHC8YCRq1PJ1fkLVfyfdNc
YoJkAGIwSQtbyVhosDoHh4/EFN0ySc7z3X2tBpP2LSnLFQ1whzI6OyEWc3C1XdtZZGNKa9WpSsDP
xFhzpGahZ8uPRmGy0hda6R+M5Bfl3B883ah18uqXMgbFkiVfKfN4e/DkJQ5WYIdal8kYq/hMAI8K
aPSCkFZrsvVVTEtyRai9CMYjeJ9ssM9rSHS48/jrV0WuMotye/rqYLy0anULGTegPsXhCppxExlM
s7B9neduo5EwUbdycKUMZNr3Zp14qslupBka2k/UxNCfFVSQWAwyeUooqopyijzv9ER2JSSQHErb
fZmDPthf5x51etUmes+WZ++Lmjex1v7JA73R+D6BJunnxEuvHthh3cx1NXKf9TK+zJamEcwa3aPm
O5V87LJ2PjU8h5GFL6/p3tn3rrbiEwgOvn1yZNC/LhJI1F16UZlFX158YLWC06MIe7nBMiq5HOWi
JuZJB2QhPLDuw4O4j+viMf0rZD8qk/RtrSwxufucGq7CsIzknC5lqn0xrcIkjniyCnvNhU857Auj
9Y2MIqAsMlSMSBUl9evMfZYu3qtHTvamYw6PkXsf87YwIdSk8QOm/EIY/vDRohH4rWmdDTlLU4Pr
0G+ZCmYIFtDivmKvpY9UlX4h9XXRaZ3uQdRP9O9HDoS/5APf5rKQ5UFa/mJgUEToupk1+w6sJ5QB
x4/1/D8Nt4I25vi5XMf1s1Fb/Z3JkS5OgXBNfGI/kcOAlKJ4hSVv0+8FKrxfoOTVMi0eDGmXBnjv
BpvdPDO+xJ0p1omVPSKtn/sZ+iM3m3Guj+DhkOSCyrLh5wztZkLdRew4GEHmZ+x8dcGPsP1bshM1
gOxewnwkR1YKuHCTA1rpng9Q2xFERUkT97jEDHZzVyNC5cjuWvt8uNRJDV2DUpn4fn3zDOo1xk9r
HRh0B34Vdstt4nGx89DFb3mqrlbkomGi4ODjskCTQQaZea2kdxkta0rERKM+A6zcPTDGwTfXUBUH
Xx829T7cZAM1eX7QSb4iB0v1zLTHGtlQksBu7U44tcsXJbPiiBKNBwtjkNpTWcYk+YyGnCgOZJUD
pJIYCOPTYE3yKd9D8UJBdj14TQoiqexCYr7dPKuSFGi2c7Ufo8V0bL5DbhRL2YsSk8RunhpVyJIS
p+PN151+CSi7wiqcpIGpwTfcOMf38q5fOzi+Knldq0mkTgKQOQLCKf4aoYCs/k71Fgwts2MjN7n3
FoMQcmGVv35LHb23l5nTgUK1+akHxp4OJ1sa34HtIYH8Qo/ibAmybqNH6G8sz2nXvotCGM+GigSE
tWwoMflQc6vfL7CQnfP4HteoXjVE2TT7+G1jHY+VEQNV+liq8mky6C9aNumWypm99VgqEJApJbnG
qd4g5OVltVm6O86t4t3Ck2nzYidj+F6a4pvqTdZS2WeLq2p5ehpHEUCf9A8NK5z9gxdgqJyQ3ETp
92Fmi6MQHpvLYji4CgrggGqKzLS80dm1xDeAuhQIn4nCloR/4v6k5N/iMRaLvJtg/TBnUMdSaZcZ
2YPec2QNnMHF1ufPb7I02NxR01LTxxpG6TKRkOm3+5CZHbw6B3GBtvQm0Bc+Znla5PNIa/tLlJje
Ehv36kykzkv7BbrZKosSgykRLPGHZoUZihHAt9YmEtYl1zBIr7a6lcnETBKvNcUxPcUON1osdTNq
SeQm6MJKJAhLm5zEAxHs+vxnxWQJeR3Wg1zZbpnSPvhKxiPhUf4K7rXLgGtQp8l3Gs2Qdx4NfAfN
/GfIVUuSOvhM/ldJXBsWD/Hj6+BUMYkOQWGyBeLympOiF6q3wLyi+hLK9zlluMpO6btd6itb9WeU
wDZGifD7aD9c3V4bESy6T76nDEF8+uoFpvUSnLPs3e+7MBNXH4nstegApSz+pGMD6HW+xfXRYBfh
cNRZ/blqJ4REOLb3TilsxzUcv8O5KEsziSfsH6niFMbBXYEOpK4j5LGtjRUmkd5U/ru/S9jZ/bAX
isE5QDkiVnTHj2TXkUD8kVDt+YWiSig2SuiqNCSDC1REIacXkrGw1jpdro2p1cWZWknaaZgia5CO
/mEW7yEpu6amBuXcS795wUp+fPaM09BJ30k2ioko0LvFxmlJXoEt/fyR7INKbIpYhE20C/0YRiJc
cKpRQJqMUy2JwL2ep0ST8zaYfPjdmGljesi/JOLLuFe0Av6tVA44c9jeePGi20A6UtEVVQyZwVnp
8sslyuMlmoxtPFRmeWtkDzya5ud/tJ2UmFk4xBsO/H1Y7D2jAf3kwrxUIkNLXZb0Dy9J0qrikCgm
ZFzDKY6Xse1obtkqeiX+3kKg9VWau3o6RX9ubLgpWVKTizD+4DV5vgCs6psepNqo9FQjbWVXh22c
6CUr7itF5Tin2KFWew8r39/duB+al2eRU/DSQAB+6eZUaALnG04PlJ9d0w4rrmBuGS/DQ6BIrKVA
3OcRJ/HMiJJdEbn7cnUbSE2HgZ4+GtCIwL20hB9ilwho8N8YNCGuyNJk9X/06QugcypRuXU6EWHj
01Q8T7JPZLfQB3bAqhl4JztFF59Bl5zvqo3uUZp0SbFkA0QSRWm7+kpdnfKlEfTEV2UDrjZ46yNI
5pD4XRdk0pGkL65/JuZUDzj+1M0ygriu7Qx/eDF5sPmU07mUH2w531zdOPT6EwP2Z+ixnpsH+gRM
jbh+ZEa+yhRr0FWSGEDiV+Dq5zz4bQ9zI+GZpCq9frstqGDcvPGJ6F38ak5zNCWyniS57Jqpa4Pz
tMOcz9dKKgXGhZLK/iCbpmqwKuq1KuvEirG/929LGFPeUlEk+b4MYEcG6vFX4cPb+Kt1LR1rGMB1
9evOmDhoVj+V64MQuR0OxdbH8z8UaWacg3iKXeva5FNwZnw1HYh8ORs4hIaa53hvSQ4sV36J+O82
q6gkTKg+smc2TNkrgYcBnW+v8VDM+5VuWeKS/VKRcogFmfFbtPw23zPLpzRVCCu4uMfvq3EoGSbn
7wxpWhpDQvn1IfJNaQaaJihUq/JZ8dJ4PjDeTSWDQpGbs88kv2u36/O874uHzzTMsAVV2uhX2YSP
hcdRvcD+bi8txBxX/aXLcJMpZjbuhMxIoUU1JuFX1LKXA52DwcgAQckFlVREkCgCZjpk6UWwZQIg
bNwBXZctiJxYMWF/TYfRpTw1vXQs3vZqqiZ4EJcjMw3X5WvUwE8DdUELHmNEgfnmdvqOBYu5YYMw
L6fkQ9eLTba6KVQ8zQiVhE07L4U5HntdqymsZnrKRHk5lXEf60x8o0ps8BOv65FuK7hdxlxOL2bh
f0PbX/95Lti7KZaIFUdOhfXYxous4LazuJz10FeieJ92K3grHZiy3zN/vupm5ILOPA9IfdTP+l8n
29IEZVvRAujppww6GckBuf8Orn1uqL8jkTclGQwT/ao5UTMjQ05OeSEbPrxc/63/XkpR0R4aMTib
jm4NnZXp3ax9h0QthN7KDaMZgsHtiblZxWCvP9v0Y2UIx5yd1dmJdwSSZfCEB1VlCmdga+uoSDFy
m0F/yX0yYLDj3XZJYC581qZZBGXd5HlOHXR11kdzYvnaAdy0DrmVcSDL138uBcu6ut13cnGdBV/P
ey3xq/cg9+usaQvsdmLLP2QP2Zel1pAnOqG7L4lzenYS6wN/PRwW4FdzI52qjf6rnlFI+KgF0U9y
PewoPI9TrDKnAfRYqhBen9sW0rTfAeK4KOw+ziOPvvcFI1xtWjKmg7SDlMJcv9HQwnoGr3bNYHZ1
+bQuibKh1SLAtIZGtZiFFeRKU4Do1A2nJEm+FPcXuQxWtgyXKrADFCloWxIuRBbJ662BuRacSDPz
zTc9EwYfVOXKkiCrujT9+3AgXONsMx0wOWfVGmx+TNTlGxS3K9Na5omwuD7Kj7H2YP49o6YIkT96
HDcgVNbokZOm0TIbH1qY1PzDeBxn9otIVP69xIDn+e9DXnc5UORICe7WvvWWjh6DRz5qB44E4HBk
ZaKtQHCJL/Q5CpCOUuf2tD1+rchalbC7nFuBLQ0Yl1/mdDrL1DVZ5CexQLgHJmgHv5Yd4jA9YOis
Ng0GSVybAiB3scJ9ySALbVccTLD3iCo7Pm39QX+kQvZfNxFzjnHEENCW/i+mxPLGfveYkYoVkDMU
WEAo9Q1Ep0qN47plRTEzCEEg2AKJgM7KeI4eTQeY1T45Dph/KG/Sy2+ktotAnUmA1SG0El5BjdQ/
M0Qsro7/ggbVAVb2v9Oe2J2XdMqSePspLN7TCcpLNaDm/bEx3uDYCLteb0IW4CQNIFNPIVlmJoZ+
GhKk+XyT8Goow7hLkS6ly+pUcu6l8ddYAAhQoPuId3Fc2gq3K1oVGSNwuUQZWgEXVjEh0c4UpjHr
Pf5pCB5YCxCF7t1FsqzC9/ZbdfJHTHK06MT2A8T6e+fmqnX3xcJMxzYAgRz7YMOvPLiVlbTedTB7
03JuJWQ6gqo5nfJR4Tm1ux/21gsILZpoknGLx5G0H8/kpLkyCjHxZxIFnQVgwy4qp4PuiFnWrhrI
2fC8aJ1sEuEXmiKfZrmVijQujTW0ANL5Yw5vDTsZhSxGefgAyySBrn1hn30J1vj7fkBa6j9HQMsr
WXnEC9AEszVKucYADXoRKcy5AfwHJQNwqeWv6DCJBNrRs9X+rAuG2lbfBW0zJGh4t+nvOmxToC4D
IJ7HAouo4A32GEKizELoDhnet8EVYwn4IzmsKveJJqw2ImB6ISuHQMfrDfHkKS1rcwoGHs9vAtHr
4YqAc/KJqoWosd1X8qycjo+HjOHRZS7HXuzBP61TNaKyl767tz+646MJ47jY/bM8T3tH6u5mCS5W
GNMR1ICwJG8lQUD+NW43N3hLkeRMl7UpuBdCk14VyELl4VXoDHVKkYRmePrnxaYkDdMycn1zQ2Lu
IejLuV0jxljQr0MM1YR76Low5uguK8fmGfzfbFn9Gp0MGk8XV9YoZxazhpBVPVOudPLsqrEdV9mI
cC655v9qbqoYljwVTyAQSIOTZFC4zo9PWnBUlL2CFB3pXeA/92+/pvF3lkHlwpGPmg14fcGsHUx7
kQ2iI6x/4kfuggi1x3aXRpayItK2Ud3kGMzM0WYGLoc2/+DXwRO5feDDHZSpLXREuYLWVT9Dyp1f
MG+BNWTSTBP2uMyIokVjMiTMpZro5lD5EVdZEIwFGMsE13YyG/Glm1u2yZWKV4KgQzD2Y+y+bMef
VEBqH8WOPuIDvnvSBzfPvjTvj6AUqiR6kbY2SVDl7dgALg3nHgiT4u4tWQ8h86nqDTdoI0H/q6SQ
virJIL26tkOu+RAJKvu7mm5TQh1rUGuA9H4sPM6Vpxz9DhdLkn3qC2UgQBW5tUEUHjBe6nZCooRs
GABYjwxrLFCvafVX1JUvO6tx7y30GK/vH7NgSutxPM/A+ccUZ/MFEc4gdQucKLS3ERZMhtIIS0UR
P5qc/lxmjziNaBYipXWfkx4ocf5fOhNTceVkA7k7ipaatAVVl9CZ0xwVMKoSoCIZYQFxUfmRlzTK
tRZgFu4RQgdI5PtGi+mhrOyvCvKWbkwBwwv2Nqh/KO8I4kym9MN/kSEUg2M+NUMFoQuwTFNd8UkZ
ifWTlgB6ukFCSJRmLHaSFYth+Wjb53Idi7ycD6vw7cAAiQDHM3jd+ic7/uHUIJ9sNMWiTFom+C9G
YBasIYjJiT1gYMk0fOXuE7l++yROdEtpdX/1wQTm9PfmWIC631zhJ95yZRCbPYHxrVkCD6cM/HNw
k/WjwvAtptbcjIr3uPdjYcJj2R8ZDQNJ/sGoJcd97uc4uK9pdbLI8nwo90RJOjO7zKGH4zRKNGMH
YhB4WzIvdsjD+cekvVSfAXHBQh0/HsIjU8km0goH3sgCoph1Vf0zdEQdp9G+3wq4h7KSwjXrT2mK
IyLahc9hZ15OsciAn/6pXVSq1FVg6UifsO/sUDXyd6WWwNLt7cjDysf8E0X6MKvpKA6VRMt1CN+h
qvJcLVb/OCJUH8qLxpug/dqByGe2DdPRPKcOBUH2qot54i3TLSlLcn8s0IRR0B0wDgZm5b5bMQbx
MP9WgN1h1ot1TnCo+vR5kmYNgzFZe2jOTVd9+8etMJgxMStGbYPBM7QwasUN2MBq9VXEntEpDVMA
gBtzN6QHXOiyZyTo1VQvujgCE8uxHo/d3NYkjnRWbOsegQ6NYqUbJEyGITihApxhuHWH7H6L0gMZ
ub0kyagRC8mntOk3ccshN+9Xkly+CXUaBJQ2IPSXiIfHhEqh6KBPI+91GxN+OqxR+d3DEJ+sxTEj
dW1ChdrqqGoFCavosV9pTjOBehzT3Vlom3OOTWVHZjidLlk8ta4CiMaMXgSf6EiAxdmwpM8Scxof
gS3Hb59Rysdaos0x2OwUBJo1vsXjx4Y/qPux1OGs6+YSeuUVfWqiRdWlo1bWSNIA1jNLqwO54edt
q5c6NwF2dJAXhBnA6g+Sfk1mvKvvJNdTVrLe0415qqU7lxQrTzsfYncYQo4ph9Qfs3dD/XJGSKjC
l4TSNwLCXwIE/m2tmHBLss59S+riwcsPdSDObJI37OgBKaCmYLSiYDI4mNtDWeqtTAp5+0tOUeer
eswj4pTmYEHS24oOtnXd1Y6wsVOYLrkr9991pz4drHLovRNDbOH2kWYgPc/+Ms0lNRnhU+Z1x+m/
/HHkDyymdORQSATTy9QRm172iRvg4/UAYFBF7dNTnWFkURi0dhqkBMTTBSTgJqzaVhUoWQO1lkfj
/yFotmKYYNKY9G52VstmJraepMHuL6utd0yTL7PBUq9FPOvTuV1n+REArlsoXD8kvag3ii9zruWh
NkhCMPp+SM4SEVbS3IByOjlP8hqwouTPTwRt56emdIYhIsXZUGf9aP0kF30paU+f5Q8lqSLGCFc2
CxWEe7Tz0bySLtcbnsXWPR6vLXmiJt/TPYYJiO6cFRNZrFiK17vs+HmTSjcF5Zm089L+7LrXJoVk
UwXLXvVumbJZ5SsEEjGWo/dJp4CR0kDqDkk/ND44442sAC2extM9ZQ7yHeXyxBobx8aLAf5DEBtI
YHQxhAsu0e/H46P7yJRUPZkmUYIQHfpfbd1ZLtyUCPnGnm/1qu3Th6N3oXpqvlj5GGC0aqzJSINB
BvyP35nvzbj1EVyI96AWUDbh2QmlN6uHRmIaT/CIB9byxluc2hFA9muzufoHVeCIDTwrSJCzGRwT
1NcZIBhBc6EGyxlS5Tsd4jDw5aBSNP85mis7QWbpOooWF756p92jItERxQcxT6xhbpXpvXRnndEJ
bBX2p3eDawAUFCCkX6pWB8NreeONg/HKKTFewQ9GYIv2KbZLEtGbF5FhDrWNeIWEjX+FvU+tF37E
6MlU/ijx1niY4WY3gvaHNfX8X4dDvVSkkJqOdKTEFM/JfLFikohtRlVJQV1umsngoQ95wG/mmQ8r
OsYcm1nG8Ofsr24nb/avrL8bEC9by9P73zafik0xy5pbpNe9mcuGxHjCppKW+d5s2x0+JpNq6sQh
T0NMzHNa3z1Ing6lj9wQ9GO0jKtanNMHWsKlhH0TopQSRY2RGtVaCtgfQ26MTvT+xhltZMD++EdP
ICb9kDM9vmlDNRfqRxOl5DHfV3d8ZPIBb8h3LhbKgnur2XX+Pb8gyaoIGRK05vBnwBXWlOaDienr
0STGU+CKuhBRbDT2sbIRS/qs6bPu4wXeU1je4W+xKbdfX5ze3xYv0leIO4aN9Y4IxqiA/CkmMafp
MxuDed4S/yBD8W1XH+i4BLO4E3YIMAA31Zt40c3KGR9H2cmEsGx9rJmpxG7y4nO5WQgyPSdkVxkq
Gb4E34Jfg/+chzeGruA4eXdtt3Pw065iIC9/x0WXxPWnjhqFeLP53AFPrnxEjHduW4bHY2vfIHyk
SDgb5UsInNj5L0/XbKgcUNnkUfvKP+CcEZ42JqJo4Js5NQ3pJcZCeR8Zh84ZrIvUORgQH/eyl/iz
IEa8NoXiGQoGllgqSh0hWr2DKNER+/ZI/jDgFSBxnTwgG4Gyd0R4V8dZ7Tbr9wiYBSt9fWMX//rS
BFAZHQ27az5pX0mr7yfkIBcelt6vV8cPPhFL13yF2TA76xXZp0Kpw4P7+tpwzOU5+BlKpHZEnLr1
aRGviWcrDTphne25pU37w4Px0QDkhV9Xbsr4bYmRWPJzyw5R7HCw93LAStelMfAlMy15KZ89jom1
NP9g5ifBeMvy6ODceDT+Nw2hq6gDdOw442gbCHqLiVWhoeHbIHU4b+D+SZQ7xxRx2cU4FxAfCW9x
yi1DWTSjU5EgVtjRq9M9MqmHFCWJ7BixukHpRSl6t4di9yLUJM0BDJh5dzhNWNNdIPU5JOEjfrOQ
W7tUkxQWZ14BZz+aGfoyrr6HjJj0jfERBeLk4f7lI1DIiVVbtKFU7nDfJ4uQs9E4y9MBNXBCtIPg
gYP6vrosKzBoxQtMy2MUthCyFXRm+6HEw2mrapitNuqS1/r16BCknr83tIiD/6xd1lhUuL0ssslc
Lpz/2vihfuuctlhES8+8KVPpo5XBcOgbtu0u2liYYZLEh47N9ydIug/TY/Ts01syMVHcrakXBg/B
CQHR3zoq2xSli9K05QjaqStChSz8LNPQlPdxgv07Mf7+SJSiYOv1/fvr1pdF/eH2Uv+JGzcIbylV
wWJLKdCtiJXi1fj1YAxXgh3IqksOtaYrRkMxPOXNYSVzhEcqy5YaaCNEJNNBEkBMW72C+QZKLH9L
KT0Vny8n+DS5R+kAFriJAn1+Kll9AfFDiiZe3MX8wTdSdnfrOjq8OWjkJncpzHLmvVDU2nV4ES7V
mPm3HweuqfheodJcMxnqPqh/6KGydBkUPUNpLOqo8qnZYsPu1zDpzuI2Vavq4I2Vpuvc/xUJ0lOZ
ZAVVS4hmPFiAlnJ25I1f1Eq74XRSlUBKuLmCVn4TWCXpWjohKL1RDUhuTbQFHOy3Kec/Y7fvOUNq
8S6bhZskab3ThuYthTKs5gLCeoUjU8FBkSnjN/xLzvbCnwkhmUCNgMz6+Yie0Zmh3zakoFtJjFVh
BiyhXFQihkf/BXNpct+JeanvF2oORsIJvTQfjK3rmYgsbiIT0lI1CpCLWr/gWCG22jTthdusggIv
oZK+WkIrSNy5sE20asdd51QAKUrrWB/xS8Rns3zUCq5dHRjtLoCd8MH461Mq5A7V5vu6JsrjZjZN
LNr9LZA3gwW59LBYKprzbcWEnpZiw3bqe1YbjttA5AXqNHQXwLi9nsXMmvl76y3rMcTwcSgnIH8d
l2u7tokKAXQ/OlGUK6Cs0fHgRuwYGstjZq5d/BmcB08ANylA1T1PDcwnIyKmoUgCmZ5SlVYD/Srb
hyMrbTW7a7ELal54d12TqY1CCUl4UYwwSvwJHauoQDpXyAu+woeRnZJlYEt0nHPeRmSOdna/ylIw
OzJPiyeRZO7rIM1pcj/P8wuC6T0WI902FqhSvi2AeSZqSfFzYM9c3GtRgBIym2ynXIiSHrdZV5L0
pl2zAEyX0IP7tyW8rbZ9BMsC4wVvl0UpS06/WaNyNsYvSEmL2FBTDIHTt0xsrAn++b10ssME1XxI
5UNIgxdIn2T8Z+F7by40/OZOtdwni0O/LERukbPAij0TbuntX0+HCIYhxvYC6+szr9tPjJVg21CB
XqV+kzMarfX9jT8L3uOIcZoFypKJhKVUUatiZ2ccxrIZ2OP/qjQaEPcoe5U8t8x5EZ84hhMUE440
Tgy7t6caY/AWJ8KVdfhKmn8+8GYAJa9EkSG7EiDlIA/9/4dDoV64M8Hk392gTbcgdV3L6/KBMFSU
vS7kOrocrTwqvDDtCoM8wXLDniKVpQPWjoA9FQuHXRH6opTbS1PGxnkHwc1LudWX8YZR4E3jvJeA
DxQLmyfkg6Lv+lH5KKxgG9Hua2qnwcpdpsrRo0dKr6Op+duviz7we097yOXtztX4g8INuGCdH12y
dPCaoCVIIbkKUMlG4KrGPci4Kz2FKkrMWwp8h2Y2mD8FtaCxebb0kDt9V3eS9C/nGTn9GWXe1U6o
FH8r+Z4lPyhBP4lSz9kk2XxriBQ0OK0Wn5x5MbQAzu5RaBc2IYZTyeWJZ7EoCsSkDZfWPMsxjYQ/
rkVc/H694DBPLrDaLC5p+cqEYdu/fx0CRIBzahNy2/PhbD6eim+jrUl+Q1nLfDLnEBYDjNjb++50
gwgFF/udpmxNvulr4VRagnWqUkAmqdvn7E+Ispvg43/Km0QKVZN/GTefIc9MhV2GPgILla9C4huJ
0hgouqr92BMNWiXLnxo/virW3BZvyPkzsHn4ubS5q65O5aw+XuuKZeYZHrLQ+llrU8h6VM4osX8n
CpebBDB1vPHoWjXMlLFgL75QACoYTet10BuWLP27WC0FL3rtao4d9IsLM2p41s4xL80l9Fq0yDoP
pkzh5T8drFHlNW57p3H5Nl0IhU0ugI5NQ3f+pTLWxqqdCgHjYc2WY7+gZ24NP07DWZNE2BsGubov
GHpnLB1N7wqVLiE8h/8ZuwZVOUltontB/vPhVWHeDdHiQCs4WMBG/hGWIURImRfwuaPNK9m4QubL
+uK5qDfLFskSnrdEqfCTQnEYFLuKocLJ/2BMqso+201NAezqmOjy9Wc74SLmad+4A0DcYcM4hGMj
CxrcE8SeqWR5Ht/Qzb3LkOfpShTvVoCu8YD/wkmLzm854dETTjZzgPUAz0rfCmXB9Yn3AXM0pYoH
Gl3GFzByKXWY2r/hl0Uq9HbQZCYVvQZlYOU/Xlu0OOEwC5teXPIVz0TvO2z+EGv4ADl5hgO9crLV
IueICz/5Cw8Lzk03IkzGU9aWBr81DUgCjwcUXpyrn4r9zCHa/4767Xdr87x2Jyn3Egc5NKrxJuCq
BR56zl4gyF/tKgDR76mSV3XmJ3smXTZWYH93dr1roHEJrnTkQaB/OLeXswZP1I1g5ADMPxDra6fn
lxa9rzsLwzoKfKxLY2OaKJ9KHabBOt4qipw7SjdrVIJ4dS6vbcCNmDtTc/lCHyQi0AU1dusr+SIC
FbciYMVjgovmy+mVw2eD07AE2kUV0nGJ5B5qw3RRN9aq9FYNXm3JGlmFpy9bPrB7dYs0Xa4R2GqD
uKcdyLbWrTG90kKKxV8+hdM7cYjMvGOSGlN8cxeKRuQ7HzqfD+hY99VOYvod3WsvUaZpRC1fGWu5
wbhJq3xOHmt/ts+9kLkp1poK9tixqpvtMrU9fjd4olRJmI4bof625e69c88aXp5ChcQETr0czIJk
IVn4yxOXH0ohj12n8+eAOg/lswU6wF/J2hAVIopltG8jbupFEPmFWjtkX/AGp++CnW6bE3z13V+V
GVSKgWxUyrLYn5oWVNMCdV0JJy6tDAD8/F4g+k5M4+07fSJydzAdeYJcefOPgTEYlZh9O4vC4oUg
wETqYD4dX3GGz05N8SySiOeeZx+ScIPwU/LKeeFKbSbqkBYMACmGzLujlJHskVwTcr8dBYC+/0Z4
stwYTS44A7HRDnGJRZEReeqJsEaINU0Lruh4BozH6XsQuuy7WQWPbx+Cgbr823jPYFSHh3vv7AUY
FpJMYW6L99HTghgc2b2PsUNV+5qMa4faXbsXKUt9M4Pf7FyXIOM/McoDXIg8QzDCEYN9hHAiDOMT
P1pGx257p4WaYSJ3cyV9gn/YdRx911/HjnESKqDRGDV1v3i5AiIWGtNP27Ry5Rirbn2ilMr6ABhr
Me772hMsh5A1ciJ6oDCs+9bylzeKxeXxQiaV1DlUHNQw0JkJ54qhIaVCaNP+tHnImtOe3FE8xFY7
MnCW/uNBUskkxAs0cnE5yhXe+Ffnc5xZi3Mi9mWWaI7gPrDdFEIaQCFeN7rEAeFmd2c6/5jWQzqh
EQuj16lLYaKmqwsTiLsYefSvn2jqF1nuET6nAjIGHfYhSlVXO9jrbGlbrtCKOlaG72+zE1yY9O8o
GEihSPDGpVSD/wc3YidpBiL7dW5sMJfGAzyNpkmq0mvo1ZIoUQMyTESnFWHN9kT4aC9hG1Bzmo+u
ExfaIXsbJztv6k76PXiL1xXh+MGCgdlaV/xxYXAsLhLK3Jhm/JJJvdIpDc1EZgrqRArGXId3Ktyp
IxmzBaZaXci4QMmx9LNd3uk1bbvvQqksSppZMJ/ssyK3oZmOaOxt8nvxv94H1VPZJUw7pQqXj86o
C7wOl7rquHGNyVDf/3mqwwxXN48x95C0GYEP+zSZckVPorquwnXQcj4y+d91+UicqB/1xynvp6Yq
boMmzTpJUkLI8eAlkvAilxswVRcUq7WxUR6tuF2j/Rzo1JaMQHIkpvsb0f5gGypjWKMpmYqP1Mqw
yRLhSr86xulfd8XJH7j8Rxx/6xcV4hX6KafllsCk1Vt0mwIiuTqhtrxfHqE8b8Kpzml2pjXJ0VKI
dpxVzleYHVaIyT6i0rZPufHXl144rJqvwFFfFa6PssFyYoGGudpPLpiZKKSl7AtNGOTAOmbAmKz/
4E8VuCxdfqHPPSlyWOMYOC06igb5qGkKUKok/Yigohpx0fynt5enAd19vp1BeG3c9waYvpdubiiu
f8a8Oa2mV8raK15X1mDb2PRWQcd1hK/r28bQ3oQp8GDE8kVgPETdKY0BsYiDVi9MgSpvQa9VGmCx
i7kvXoF8io8vmHoG9Dw6AasfUbD5pGFHOAhuMsp/xVGvfvNUXiHCq92eOx0bPQ5UfQTtSKDHHRBb
u9+5ObF71UV5GJrJbk6/2lHV9ZhMb9JgqCmV7swvQGqt8WY7C/c2LdZp98OOM86BksIlB1BNPH5/
ptgHRlNfzobd149eXAocH/FL9x3DWSl8LXh8YLVI9/WmSaUZmXg+xC9AsISh4Nfi1ptm5lmwH0ha
23OrilrMusDDleNe9yIfRJICMaqU+y+P+hwLCrVQ/ioDbuxWgG6hqsiNKTy/7QGiBjZt3n97TkJi
PQWZkInnXBeDtlMKIoujmlEVM13LY/4SCAXjeWTMn0IFo2VDUrJVU+11rFR+I0L9ypnj2z9qHYV2
yRqQjTHlshkw6q+8TEs1zm7+dy13NZHVE/D4pF33p5XnOndDfe9oa3FnZgjz/B4Kw3PR1h4dhubO
uyMkA0fb21a+9xB7gxY2q5jPHjAAYNGxYp1QvKxBeWCgOehWQIWJUCrdfWXAQio9zuvtCWKXdhP7
TauyAAhDJHWGn3ReyHcQt9fHGgASmrXAL21/d8JA49gauA5FvCTxz2rqDQBU+cMh4P8LCkHQx/NX
/7spe1BnC/pKAjy3Hvkwmaru3Xo1siXWOKTDQTq+WKRKYoM40dIN0abJaxtqweXS+knCLgtPHPaJ
wpiHY+dhiNXbn4578CUj3XNirvBOcw62RTXw11YcMpPXLZU6n8Gb1loetnr42mvm665LCnaeahDF
/HoMqSMqpEWPqhYJfYXNdvGTxuU9SF9iJxVzvPXYz4c8EK9mDp2EhmbPBbaIJvIGS5bACn5epCJq
AtR5d43gMOoC8abLiWQLXeoYbia34FzKRzfKicyFl+0JyLdyx7RXZb04C3JQ/not/yg9Dgx20I8c
3kIAYeEt6vxGPFyqo0/lHXeCTX+a1LGJwjMqk7245juFWWpOWWVWxZYIw/PXBZ3yWeeNE3v+j+Lq
6z3xUgN/TqWMVMskAHQAHSb5u+alIcxKkae3ty62w6CvHchGsyzfzDssllbwxnDJULTyqgbbWmQ0
DFMtEAu9JJ0Hy+gAl0oWogpbYN4anP68bhG35n/nTPMPqzSrpg73np398rlV5ITB4WrpnWgMP4Ev
S8fPoht5Y0EB+6LXAr8DyD53GsCKjSl2HQ7oiZmP2loo69Jl213okSJkGK/bnPCFrB/8e9f9bJMW
IyWEv4OKvYmxCpZEjHyc7gG9ixTVvVSI85q1P5yBjUcY+lEZvT+1no/EmT80NYdRNN9/MdvrxWD8
mJM45IO8nqMFP5acBxiMPkglVMgkkRFKoSXvs45McMGrJJHvw0qXbV8LAUi0VFnb6niEGTrnYWIH
X4P+laP60ehcFOanMQA2zMThxM0r7ISu03da34uzRbStUOM62LyWYIevmpBAJNkclRaYYGydKqfP
OH4hSSdF3GvpM+cfWKHC4DKpKFXU88bqiL+vy43oDmBiwwjwctHD/ACQdb9E1YRLY4GBUj2uuS8D
GXj66b0wlk7zOg1sxx8FBug+B122tSRavCAHgRRVWQIvakSpNAivW12/21eZwirxWVVtZCQoZu3X
tEhjm64UuaBe7u9s3KNiMQnkyq+waBxKtU953caW3krbeLC1xtkrTCxeKNzYxKyfNA6WsU3StMNn
koMd4md57UlRET9kQYPAWqwuSPaCZzibb3aGZzoKosQtrEor7oMc8bef+OWm86dgRlinBD7OlmNq
sPqnW21Pp4ucwaeI8zUwfwi3x4tGGtHwQ5O9A77NglterS9oN1V+tT7B2ZUjCGsBwwBtnn8VPKhx
O9xaiu9p+qTjBkr0yBvRwIPOtXVFKLGhjkvS/ibdene6fognV54o2OxARqkpXP2z9bHd3WrNw77P
uYkTxFKlBiiu3r0ue9xnB7oYyVuVkpKT0d4XE75yP10X8kfZmqApWlTYdJ2y1kT5mqRz9g6ezKkR
VIE1UWL6036JYvALNSe3QoRUiM/l7HVLX9M+6eILKwhyk3XciJ5/ol2FZGjITL8bfZ6qfTKYRpU4
cmEjo3gKbuwwidf6juAozVS2BBXFNneWNOnrYmd20EMHjzxR/Fbpn67SROojRb300nz3/r7oD7Wk
qNx30INXrsih/CVHJwtVtjQJPZZ41l0r/GifL0mklQPvYi+0N22ZRBrdtn0c+puqpAqv/5gyt1M2
juicQTiiqVEo9DvVn3rxsLdaHd4HqBMS+a1t8AssOlZNwF9OUwPXBoyQyi/mKQyxSqMY60XuA6ID
/jaxKzZMeUUCzjxtIK/EzoGd1RGQEl6o92n77ggCNWW3iVHvdHWWP0H0sgLS1X59X6Xqa2eIVqrF
k0w2/ZtVdhpy7aW9raTiiWo/ctdpwMg62RBFduMZAT2wkc2jmvCkK5QRs2DM5a2gVgBUOOOvW40i
mSnIUHJlenOIS3DGd14nU64kr64YKHEVH2uFDJxBLTMK1gHAfI0IZSx5AES0u4n0Iz8ZeRvWBPn7
4CoyUljOBDCPXb7g/sginDt8QogVTErKpY9OlP/PRPWwbLyF29RNWp2vFZeLO6vM8XOcXe7+U5+X
EbK5U2qmw9Ga0wcPoDChSaEVqYCgUmdANawywUHJZrbD5i0lPREDxAZliIR+M3fjAFhUQD4oAvSs
UjhP7eZ/ffPbkZzHJoyvXQwhsOnIulzdvrBrI1wzDPxp2NdrjudboJTrSXQyC1GAGVR86p7vyf7O
WFho9k5gibsWtXcyFsXEWiqx25NL2rwM/QoGn+0Pn5cPmd7VOHtgeKEFuX4aO3lJDJWs3D+BtHON
+eDuHW7nJMTx0IYDJGnX9Nj/9xL/OB71BdwP7csQRZEoflACpm2q/pbvDVjM5+uP8ETOeAB1Y5IR
lwUR56dP1sA8EjJftXbSsg1OCF/pZRFfJIhczBGi/7b3NvN1Z9H0uXjET53+MionkUmRIc/UABLd
61xYSF391keP0kfl4n5uyTueBV4BxduaeZVipLJpgoQkiGI9k+p0H/zjqCH0Ne2IWDN2mXf8V30V
bu26EbgfH6ppIlcWzXjF9OsrOchjC3wghWUGaI5hIjirvGyY42g8egHD41ePJp1n02s5Kuy/LI/m
XHVLDV/qlBSB4WFupZXhv618CSTgFVuwxO2PCqy9vyfG9KPNj751LjtZ02OOXdtjkrfSzL16uCbY
qtW8y+LrC8FqQPFggWodu8470QOL+WVI1y+uiQ5PqAb6T5Sni+EqyxBKd37fl2uP1UJywiDxnBSw
3YUQStgougnQoZ4J8iQV3Q+WOaxPpCRDFTbBg5Wrxt2absW0rn6UiIq7pLveWcsEp3e760c1yxKh
iC54Y9QPKbvSCrwlv+5kf+qqaz4lRThG3dRkPgYGHkUwGJd8PAUnJ3WSmQFLHlaYVofG+7RyMDAR
e06rofkhmZE2f5lIl3tGyllQlvsU4dh0MzNXwviGDz4BS0wkG+K5aW5Of6Lf+hy3WZq5dPcWyrjc
D/8tavnhtBRX6J9FRNyESRN1t7QIRzzoR3329nBkhhLgDqSBI603Ei0hJQi/QWlo0RbQW6r8czR1
2YcknT3Sw/mI374HuzmKvinSXn9JWGfH5XAv3cDzI2T1TmNcL+TEA6OXX5sKoxaehx+rZ3upO4PT
ln0vsY6tIPiI+q1haS82R9KwugVffEhsdptGqfm6/D/BcPK93+7kBQ4QCKph0188l0NggH/FS4ds
6Q5k0EaMSKtrXZAIgR9VVuUbwOzbLSX3ro4aYjlvlCK+GNy7pFKFUZ9a7DJadd8BUXh3UMUhKS9o
6S2CeTRJ8Ekx6D8vA3kvwiDTX2/HsLgJO/XeO5wAqHWZMQXIFhV9gtcg7AetSogO/PW5nMWEZg+f
+9v6Qq9YKhb4z+owdwZY5nO+IEeyGqhN+4wAY8PekDsz+vHuvIvKnRDvk3AiR0eo7M5Rj5rzag5X
2YREcfquwGHebLUgqf8s4r1VHPE7z3eeDpheIAhuwShX/6cx7H95N+gaIj3AllNxOBlkP5Is7X2N
8dIE4Ov20iSVSsdS7YCPu+fU943jWsRLZhSVvpv1VZC/Ia+0PS2/y9mZoOrCMlmv3QsQRBPSgtGL
wmYx8TsJ3KTLTEq4dBWRL6r+iGsXGZHhODdlwntZ3PnZXGwBTCOEEEV6y0SKsL84nrZrR84+/9dS
eKHN19GakAtxqqici4A0+JBOg4I0WixtlasUtgabKtwZ8uWhz9QWfKuDpLFZBD4CBS6J1u+3yhyC
NjpwpO4Gy9/i0woe/GosLYhKxOdbdSen4igX6FRLHXGMpZduKGK6ueTjFYT6/jDYzyGa6PzRJ9VI
/Zr3rQB3B2ZoCrpnFFxgOCQwqSHsEMswB6tCHBWUbVPLIqw5OG4Tqwk8sZE8C/6NIqhnzGCiHPxf
RpH8oF81L9Z0J9aa7uyUTHTdID9FV5ClI4hlaHigFzMDzQhLsg+yprzPkJLSZeTsbKs72BLJaIKg
0UDjMUDJn61Q4a3tXRhRvYXXFjXtTl1YMs5e1sQ6frBTnTPhUKp/9RdfHrYxmxYOTjA1UcyT7r+x
8WSdrkWWQK19dI0TsKi+0/L4Ji5j6EpgqLxYDYJ1mNMD+9hlqFtVeUNyYkxOwyiUugksE88hkef2
n9Pw9Qcbt/1ZmLNJW3h+dKi3//B+A/vIpud30hT2QZNatWGEFoOVyMiWfnJYYlYHn0FY9oHAw/WN
KC4GU6eIN9w4sXoB4j+uIKv7QwrsLF0A6uoS4q0nOT6vBCMbIgMcN4rnW0ImMbptPK9n/9/1NKuw
Q9t9tfdU/mdElUaahv806kwCsZbjT0aSQ/F17ifYUUAL4YQih1Ks3qrTvc+IiTGqCBB4bK2i1yXO
ut3azm6eEwsgRkYJr+7bGnaOlaxL694EMSAhwxE+vCe4bF1r01f35mAdOvtw5ns3OfOgw+CTxmTR
2sOFBCD35yTkTSMmkAV4+smxMWhNj171B7tK2VOxluoLLI9PTf7g3mGJwnlfIza6eegZ4MBEc0Fn
9LBy60QQCeGDVDnuQXfQu4PdwYiONfpKUZO4ejb+uUEauoVcX9wRM6RvZi6oDBrNF4rZle3wwMY2
LXOrsJi8sYd/Vypr+O3eG4QCgv9pfiJVa98e5ifTac+ARcvolxW50uMujfBse8laGzlGtmOZLTDT
u3oEPU6F0+JMUZ9c5zIr9zj/zG7l8MEXiUq4zPSQCT3oEbI0y2eGYMSBTtegmlu+37VQ2T5t4ryF
z6mZtetPIaPyVowPURv7rpPXCGLrCsgPDnLP5w8McHrwXVJLUGaF0baJkmuxkGlSpcjBL5wjabJf
i7mmhgNnA6W1KNIZYLwCIU0dsBuFovJxYJeF5F29tRJ8vdpWFDZNWRhLm935b2I5rDjME83txpMh
jUjOFmxxnhjOO+NpCdQ8/pjs7FmEgrl80LXGTPFu/lTmye8/xsoU5BvwxRRh4ln78dEErFcj9VP5
PLvUOHQ6hycDSJ6W6NmtLi/Ayy0Alqk8rFkUKu43t01hEOaU7D+hrUpV8CJls83rUmQlQMfOR03K
O+2gcoWsJQaluP9mNEJYB525CHk6Mm48/zgUegN7R1BV0Upf/NwnEnv47+dpvg1G4pSXHdR3ngdt
4PJ1RN65WxLCCk88lz5j/fTePC6PBcb4992GyPdBk+T1l5fsmWNH1WmymEJyJPg9Q5kllNy98LnE
fbLb59zuzxNxi1pviN4K3qSCEyfXCTv+PG5GXUTjRWs8fM/4lQPuC8FI7UOZ7H07mHcWUJa6vhBE
Cso5VKi9W9X2IU4R1UY6MwpMbnFp2jsobFv3r5dc5Y86d6iyNA8aJrBlskmh3/cpKxkrQ7DkwK6w
qh8blWzFxqs1IydwcP0GpjMxKZmJB/yEtk8wVViLE6BsGlmXM4zTPcR8NuhGLN4fVsk/ZloouChG
mWz8K+p3B0AMg5ETffeOGdBbHs+mmB24VXbrIbaLDE7jZNInk4pXCLKxQeJSvdpywSoJVEYPvs8Q
6m3sIfH17KGmXppmfS6gjCP+id5t4Yw2MkFb2aQRy1tmFR3haAJ1dfPnHwwYnNgd3opGWGPvRidL
ORAc+pppWBqV2HGMLh6hutYbaMsD48Br3GWoK2DEkMV1ZhccfCK9t/e37Uo9Q5kK3msVF+6tXNR2
2DUgw6Glj9AGbRy/TekESwjA+8aKXB8u7SkqboTIhVQ4UO/rVQw/D/WbWlDk4uuqAXLDsMS/WR4k
TEXfVx/dWah3HU5oLmeRtNTbVhQ5eKlZV9Ql046lu80fvkryxhblWmTPYlMv/R2j1gSezLV3NAj1
5u6vd66V4LIcYTdzI4XUZFl+P6PE0UZ8HjbvuIYAYJ45gDQsb1f9CmcRlWLfw+s3hKIfJUslyiNj
DBNIbA93yuhfRQxrb0ERtgfjstCo7V00/BIx4jz45eIqy/RxIWmWMDFNlsR+bXNOxdYhjk9+0nRl
3/nihHGkjBhok9ZG6ZSoJr0Kss10BOgX3BJMnGD3CyJKa6riXYJVfueuKx+LRfG3LwhcU5AKCZAp
GWHlLbez0OOTyW5rHsEhOLmkD/spyidzeSH5pQbBaNkt+1TB2FyfhQ/HmVrNzVvVi3fvRphgLwI4
+5efF7a5YkW4OgeZNAB6AFznI6yCgTn87vzBAJv0F3ijeErGSfo0Bvp3kTF3khMT/UH1slvXELFG
gOrM4zXoyl/0nyCgRuWUTgppgbiJ0MOoHPs4+21OT+b2+Yzt3107EOoXtFwsa6yEvzfUTrouwuvx
f8sx93IPfNLLH5s+Y5uotcqwGZEfIxuWYPtuTaktNTfpz4VoJsDS67VL8vSfMgDSBO8nrooS7FlU
A7wNuyi76iLcHvl9JiMyJQlmv+yp4HHJgfTHzBuFUnJZadvLfgRIPfTOH5nfbhMIgI+OERRUDoWW
vLS0pU7V7SYUFdnXBb3EAJbOgFyUS2Ei8NGiDfEBgQ2nj2c78kGBxlZQvIXMG2uAlANZTIXsw8UO
U+cpkBlwrzYASLsMsDyQxTZfc9c9KkLhk/xLkQKLpOLnkg2p45hBxwC6RCjdpP9NM0RSHmtN9fxD
35F/+fsPd4VxzqQUY+OME/b63hcCNwjwQ+V+TqVeHuy/s1U58FwWeRZYHOE+hTon6fa7CD30E4XO
ZH+3M4V+WicA3QSOdPj+dczfB71knTa3Z/3FaqdYVACNPIdboDjEz0LhZw/4oJrF60qNvedg94JX
j83vg9EpZPyk7icBryW/ccf5wRcasoLx6CNs9wG83jZmhczperPnrRGFpa1gcTWTMBRlOotLv1k/
fXkt0nCotIIVHTdr3eP25O0fszD5balVas+TYXhBtxyGZn1wsywMY7ZAtnGhy0ObA7FbkMr5z+Yh
U0B1fyhb6TH2lqOGBgNL930VL8RL1A9VEQzm3bBjyt+3qjl8xaFLRgCyDy51Itr9Ns20kHQbkmVe
CGMrvTbKQcxbJlLEA1HF5qa8zSLOdhJh7752EUr/u2U4nhZjfQAxbP3+Baw7FxMC/9P/7iJxJrzq
WELXk4JEseZnKOr9EU6gRA5o3gXu18+1NrnqaD1Wb6KdtfiuVPXn2BoyK9PxzabOYHmZxKpa32JK
Mrcku5yJY9S/nkLuEyVyH6vHmRkzX3t7dEMu1zVD2Cc+2noNtNF6uUrHGIHB8ScN7baSK2kxu2j5
nlbnFSQ5go+Ako6yoEJeGGohuhtQ6MtdsehJ4Lhmow6kFTvxxzdt0Ic+ZGLjKeqIOwpD3f04OLS9
b7et+Bgbybsk2Uphi3lZdZZas9q/M1OSBxY0tHd2ekuB7qpyhTsovF0WBBjeXAPynoZ6UPvpGDRU
00fESpOK7EpmDV4KtEWFtQukUFkmRWuKIFAbj/xo0Pa/yQgE96+GdvZH70khbeup7WoMyMKpqvBg
GsA8Ss1pUUabqIs+KMQD4LVQ01gL/gFNxDcO+Ojec9hwrqevjp5hlk5Q8fwlXE7nR3Nt8slb4b0s
jjWgV1WMdBIv6GuJ2SgNTF2Zz2541kgWd2QU0Yw7j8PgVvi9SshN05oiAOogJnQByR0kruaJppwL
9N1FJyKYItac5f2ex1SfUpIqXVmOEdkyvZywa0Pa3ZSmAIXOC+KkAorOR2X0NwGCSP6douqgAoxh
loggUxqBgs6Ri7qf4kokDTfYHuLnsAkw+cuq9oBZ02tifQmM8s/wnDkzT4cDodcew5P6ZbA3aO2l
xk/Pic0e+2wpKetAmCok5b/s/65DUTR9I4klFIhy8PNVAtpD67XdF62tlwWjirHh6n3PgF1Xwfb7
vb8SRn2pKSIZKrA6uvwPXWVit+fDmzAROGuitoG59qgh7WAwtZ3kNBXEpRhxQu49SFyJy7SG8WOy
beCeoJdC1/yiscpSj3cN5+TwIUpEuF+V/jCWwXxcDaaduMQsssqHN0yQIEKKoWoA5GD8bNiVlORk
/pxplKmEBh7WKQi5Lc/gvHndqIBd4i8EkBI9zAeKewLHv3xLeirBoLSJiki1l7sxxraEHiymMJ7n
4fn2KHOJN5QONLB3bLLZlH/T286xaB6BPKIMe5krKzeTyXdXS9h0yabDy788Zb+TfblUcwrcP/8T
PWTPQr5rvBD8Kfmm1Ur2RM0jXr07e6DtOnOB6fP3uJssM+4GioRIPbsB/a6qwrtS3xIZqR3fjzHW
bNpzYAmXwqMt4eka8rTxSWtDYbV2cMEERppxof6jrtgCDWUAg9p/HRgZQx1WuVMVcvk1WlYbHp58
wWvpTfcIW6wZBV9hgEgNvEwhq7heGk88mWuVysT+yVs+lQbw30zswRzFy1GNbKej4UNwrWM4WfAv
w/ispDOkjN+9h8Tmgtxy96yLuvagAMbbi4DsldRy6hnxX+hjS2Eo8kZTRI7/r0++MOlrFgGtO0gT
oFu0iShiE9d0C6ihRAeoiTWy2qkYKsY2MZwkApS/KI5nchj9A15WDLGliv+xfDSZyLxdRGuA1RbS
ykGosod7vYd4cn/14VcTYNNKC6by+VKhKH6lQXcCSUMxPzNWCDdGL8OW2OpC/w+SBtxl+eTw7an4
xwXZ4VBxL/qm0dC4yysH5n7U9meZ7kLABit5r5JsdQ5P8Q+qM/YRSJZx63y9SAto5juUMbDdLcte
1NU9ad2Kd1cu7sDvO0TJF9SXl/04q6KnuFIMUE6rWVNKEIVTiAWh3FwTOxLW+yOxdJxPiRhJRgIV
WUwa3q11Qy0ZOzE+SEMRArbO40meig85aHU0nYPWtNDPyAGXaWbuse2PKCVGzlxGvZOeJ0fxMZ1w
KwAn2d/vdBgN77jIvAnd47+Uj7ZFXrGl/4DXtCPx6w10DQZbUQ+HiidSjPMLhCxGcw3mPr5hw+3e
rVVvyVj9mf3wbyyw74q8zrPui8/Imy9TOSL4POmPrBC8rVzdGIf8oKZP797TEN9OdVn7WzqH0H1L
T/F1vXlEhIvGF3dhklHLJ7e3rSSy9rwjwXfCn9QuxhT+q9mp8hPhg17k+LG6Wjg4YJ5Bm8lZXhHJ
dV1BLVHJj/WA9p6VrWcS4JrXfFDV7QAEf5EJZkOFH+67+bxgPPlLQBM84Cie5YRD/7u3cSZs9gQ/
e21NOgdR5/1X2n7FeXxyDi9J8QTGOzXn7en+O0V65OWd8L86+y43RWIiHcBo0c3AUWpQlSrWoIoF
R7kdoqkQdrih6c0yEXLDtMFyJqwTODMDvdvaXK3fn0dELBIifSfXljLane42MVf4NAv5OgSv5non
3V1DZoKITtgp4DfoYUSzS+kIo6DKQ+545K0JqXhvv1QBeNF5aWnZf8lvaLgDrXXz1mp1K5phxxR7
zqYcjfElzd+WaRXfd0sw3FsoQYOzuPehtE64zL4HSGcCFobDmKivR16UKpHdvKPSRH8zHrFDV+HD
65fiECbm+pt4mopgNd4xj0zUfXpoke3m+vF0KYaPvcmBUzE1RgihKj0TxOA9mhELRIoamygtFg/2
ZdP5dqSyo+7ouzVBs4rv3WjSUgm4lnQY182uKOl1DgAFDh1cVvmV0lIigJ9LgTM0cZ3QhR3Me9Wx
SkrdYpmN+/ire78lmDa5OOqF0LkZ4ti64gwDECCFVKKJ4g0ZIrJohConTioElLAvs7Fhfyg4Cb/+
cAXdm6N3kzArhoI3SkR6OEqEVoUqN0eaRd7jgIyL4OHXX+Os4jyRALwdTXvWNBQrxbgO4seNyENK
XlwoCy/thwXCGZP/S+dS1ub0yEId1+gSL3K+04whft/n1fjeOUW9D321dy2aWhjsAOyiOJ/jVbXe
5C5c9195JNlRHoVQq9GqnumzZkmnedFPgFhUtgWYRx1esKJYyQgFZ06gYlDo6KSgj0OClc+3WoLq
r0KgWFuMOduCcFOLSHAwb2kuidTw9+dVWbDuBiYjsoNoWYYCmDE3p6dfndXIP8oLROvtioz5/OMT
FoD9WASqxcZsyCX9JeEp4QundPECY7xqd0GWj1T0v6Xe/Ep6hiMAcGVwOnPHMNYPJiLZAlS4BCVm
lemmCDX50NvhLjftOHKPlhol3yCxKLNjjDjfmQJoSaRGNgbn+uaY+PlnlunAipWXoTUXWKS70R/F
o4n/gQSOHXPlrFKsZC3nq+OPhYmrFqvXSKa6da+EfUzHHUImArm8+mRH/r1tl8F7yPBPVyxIGpdZ
yi/8ElKSBpr+wV5jqVxZIodiUykQ3OT82+FcQSBx9YUdUoc+zpaoqmVT1D2eP4LNSp40jHtTem0P
ITqF2dt2O2QT+5ZTdQoYnKS5K4p7T28OyXqv0ATAtYP6RludHoEBr2t/Yu7pT4uIQ74U+PdIk5sS
JBAwcPDah4QwbhqlmzLY8JBN3vUD27ZQRe52zpQsAzXY64VtCjkT6ggvsaMe6R/WZEMogSHWupbs
WXF9q97+MWrdXU9b9R07j+nM+QKnv93Cahu6Ziv14rqifBlSu4p40ZxkEcmZwfk5kuWsI1NvzsCn
sGghKx9zycISrYdIvmR6nOiKoCveaeZB+hAOzDrMfXtgnGu2wZy7uVRNuat5c7c8NlRIJmf5G6L8
QhZ5Jh8GK/03yynIQK4lusHauHwVtjjGfAkkrvVfVMsPkW+xK8oFN5oWPTvi0BzZpxycyUb8JS9V
vKmAkdKw/StDLalalwGlAjYLqUatvwzbCDk7vnDnUFw8OIXb0z/5dsVPw/BM2RjFVR5UCmyft5Nn
WYPpeQkbraSvWvaGb5P+cHDHM5Y2W4AQ2PY8WD3xoe2FCfEdN623jBmak1BkiFoCATEhrLKr+FYk
tsFTUN9XRcUo2zA3NsBSGjrWBSqBIV0lFdnsvKuspwz2vQ8Pi03rVRccTEZ8luaztID/P8l7IRKm
MykDiCv5TS2Pbh56PSHQ9SXK8IiObkc9wXZjAUQJin/jqeEwyYP0EBHF/rSLfwMBeDJfAO8c8JzL
VYI5lmnovdUoDVih+dEBA00z5B1f58rMIHzjFIGXr9XcR7f/C6xOS6h8Ss0guOQL4GmLK4Z1uzIj
R2YQ4UF4SPd4o+PLzD1xNkVVIZkFD0W2zahkS79Hdk3Ef+173nNg7OD8ZP8wuYgPQ8ZseohBwkBL
3v74tpzKpYAN/R9++vZVjYce6R4yHNUglknIbXZp+dngIpSwwovmPz4XqMuE5wzPs0Z9F6l3VXNZ
viZ9KKLt+KIxIzG3a77dnj/r2xMo0v6PMxIQnPDS3ReO/MgzuXjc8OFLxNybb0J1VFB2PhLRRNhB
BihL3uIX8wcLrhLWE6wxiG77QHsDxpaZzFP9X2gWjXAV6ZNw+/e4RtQQbXDuvPnE8FCP/YbfQho3
YD2GfHr+XEcBdMmuS7KcRqFQypahx/WlvvVYkL35+fwQlWNz8IWQNlfuU/rj/vnu9GvZcpWcIUHJ
Z1H7hrQSepx5Fs4NDaJglN3aIt2Fp+qBrD0GElQU0q34c8nSdM7QVSz9sYdDc1Cv5/ive84v6KAP
9PFMAw5/UPASxO/wmade9iAQoMNXlZ8uTXPQz2hxVS7vyn1YgrKo9up8CSJMJSLnOHZo53hhRnYH
28qTmk7AogZxABUuNEzkms0E+h5+9mfW3eYgmOyNHXtEaIbTK0qI3EJt68AeF3giYFSEn8LYya7A
YMWreF6eoDslb/70Qx/frESfpUfstLcSO5yG4HC4LcdJUsHxlhle0qd/hiqCapMR26y13v/3IUsu
AaP2NejI57/m5k3OULYD5Sz3G3PvGgOEMlOLzrX/E9s2lz3D1iHZnPH6f6r3mG474URtikUMXwcA
BO2QgEI4kprfXULZe+SG+lvJErlmIgXLp6wA5Ll7CONBHJfFPcEX5Dt2qtDYqncJnsHNt62FWdKG
B78TSNn50vb88Q7CuzT8g+46VTo3CEGJOoNApKWKCTcJ5jZRNiB+gY2hyH4HtDxrTt0UOJEeDY3G
+joKDnImYwYEGtRT+Am7bYhqOX8TLm2hr3C0U6OtNRWcnH+yF5YIJhwxTF1i/zYQhOb59qm7qqEC
UNcjSEBlykGHG6yl9qOBb/UQgg2jQzMCqs3Yns5XmVUeuPtZFVRTiIA78Jsl9pcyEKyiyL3rcBHn
RyjZ+VPu8FqFqpVGgqiMNshDSIEZrJMwoHEDeVlE205a7x2+kdAAj3+DUHSRQDmatUT9aTY0fkKP
BRzNtIQW7gBmJoCNW9HO9sIAZiFWZiG3CwB3gIbXKeoKup9WDkJZWwYAah0aUS9jqRVLV4w4udOt
YgVgiLj2sCyNiKsGgXOoMsSUeymtgr50zkNknm9l/q5eq/Jw/W/8cjOTknZYot87Zm1Qv5RwXfXB
bSqvpfWbHWRBEvvIMfRiSc+bIu2vc5wYoYCoXOstB2ERKhrLHkba5q8gxwQIo6bDlHgOR0u+sK22
FGcdb44V8nKIJjCUFGFt+3lt37h4dV7slGn3pdYzZNePHhFQP+ErKtBWKcKr/Ni52mJWbnp5I+Ho
8Dv5uzYpcw6gXTQ3oDX+5e6cYLbHDUA2xWP0OZEAY/rj/LPjD7HOay5UJBZTKcRqGrflFp4OrhDL
5szU7QC4TqDcXmmKjPhDmpjkDEfpTa//gnjKAqb7//RXhOau1gzUlwUnaSSAXTcOO8bVHcGVnptv
TbGBOvhotZhN6BI3iRGjISbp9rCbmx41KaognFOP1DemjjYCMU85YVGJOgr12AkQUqoalSCPylf6
4qgkOQrlecAbfgku6LjiVZbn3m473KMrdcwdZx+CjyVWceYKKOkwREDZxO2NrNANf2tmDp9UEZQd
7Bm1IIl3FZi+ruAPpk12h3sxW8AkpBSMjlefs47ynIt6MSTUbfxzWGnlzVDFRv1TJh3yBXyvPs5g
eCKRF9uUQWXtAUY84x36foLnpupo423Rm8lN0zTZ3cTWG8eIKZYP7gexysUrPB9uPW4ToFRGw/wv
8Ic4Qy1T1K3B3Yy//O6GX2MtjyOl0r4YnxBp4hoW73tj+8WCGXfZO89IJqTpzpI4inF5f1bXrNK/
T0+HjQerdUnmGwK8t/rKDxnY2md5CENGNQce7GXvYwJ99kwKz/pbwlQHRqSmAoZBFd+TkVrfTY3l
FRLVomS6e/zNef+C9p3q0SUXOQHLOAb8J8cEJ0gwFrVEDnG8nLfCo6R6jVCGpza0+NiyUb2a2dIH
CTjpbShiht8iFIbYhLwzd0/7G4VW605S3Ho0NXZl6wCNJp32XBUBx6Mj/92BF8q2lMLWa94yKOBx
zfApyu9RSFVjMiekOejY8g0b66CWkG+heEUv9+LPCSzZ0EOPcHjUNAuU7ZD4+nSL1iOCCHZJ61RH
f/rppGLTynvGPkxc8dnLFfjh/I7HAx1Kyr9kM2mmdnPB2jks1G9OefBteLoFx4PeeqFIHQyoY+Ul
FYq17os3uBPiTlG1NehwukgpmK4FwO9dImQwXdhDWTwl57orfdo4q3EyAqdvv1bu7cvmUCH6eGK1
QBOBnQgY9hdrjVYcVYOVBABZmQiz1dxq4xQhaHR+1/z7z7u+fZUzppEgRH13QDc/PCaVLdlcnw/C
oPbc48RJ6Rzj9Kl8o9P9QdgIFkeli5mYualyizGtFM+QchYye2C11rzY/GRyQpbigKN40DX3mpqP
xuxQgVrr4ZRhLpGbbqMPWP5Wz/kY+fTkfHKgvQO7ZEDhH84mGX0zNvWIWXQ0lJJw1dMt+s5ElEtk
lKlVUNBAcCjyDotb0wVHZzMfyr04So/UbnAYgqcH1FP+KFPRRupM6f6RwFAS4gFAafvG/+oqvZ1i
wqWBmXDfpEdofiG26U6q4eZ1XatvcgF/Ok5Glx2fxvMEJ+e8pLALOVxpcUpibQdyUym86eQI/Ndn
lxt+W4V3Xfctr9mHprbLbIFxOKjkoH5u2CzJpitOorNEA9sevc6J9enW5slETbYOTjVZfUIZVgtx
+VskHrfDsf5OiFvUKJjK09aQSjIHsNEmhsITdOqB4dEi1kC50AW8FVzSCYtMqKXkmMLgNlQWrk/g
kM45cOJjlsFiF3vc74yYxTtWx1z3Gd2jfDaxjGZr8+asGK7H66FegM8wksRQvWgOtZZq2JDcrCu8
xSB/3uon2D2yElLYAGtWHjf3wHzG82DFwi5GWJcarClkZYSBN5BD/3ufhmVEz2BKHamNFE3GoXRN
rb3a7UHs1KnxXrsASNQtsUS58FfbgTvMWf5p9kvEUOpYeFz2KNYTOZKXp6bSeB6KuYT9nQBTn/Ei
rxQsJP0ICgS2g1JpjhrCOfPsvTgxVYSsWLv7zfK34wNEWii5WSsX31FQL5PEq+q9BIS40PUhu3rv
Db4dhNH3bE7/MvL8idgTEYKWXlSI0O+xaB13kimZHmxHp71uzlmalEaJitmFQqCc7gSL8/g+PucQ
6rL/MTBk+K+IGuaz4HyolZNawlK1t8F2ZZqHHWTrKprg28cbIbixcNZDK35LYqL/44mON15aSls4
SF3p4MHoN3SfFKFoj0mP3MnLTGwyfM/tm0TGGyYQhkOV9FFR6N0HdD4wFWreyFva4siZqU5mXMjF
Kr7vS/NjjABq136M/jZYUdfQqRCou036lKLvZwcZFc35Zc6m+eo+5rjwssk36WcfAXqvOK9XMn+/
Whb8+oXz1fiuLcOXridPds5ESwNmnT03NmCOkGqa0VWr3RG/uDAcCybdW9t52fcZtl59QPMENMWs
J1iJS5HS10640X2apu3/sZapdhzS12SWr/mbsgNnvVha4bdoZQ6VPHks1d4w1cKBth7gCNR83ZEu
9WNIOl5fyT71wJE5u5iYWWXbaenMNNI2CVCQSF9heKJwiGhu+jec/cN/lf6rugvu9V4M8r5VsxST
7avio0OanHYbMz8e9oEpp/5kai2usSNNI5CNgIip3hT3oXyzjIKJGkDshok1ct7a+sum+aY0tsde
518ofkVWwjJtzfllC8Fb75uCKZ41GJdsY71ldesi+3+9QO8YMlq/BubHQqqUMqsGap+/9GqzmGqe
1/sYERWaGd5eUH2oVyTXvFFU1ShrHqXmq+lOOJ6xfmCJrBn3S5BUUM1wSSSEci/K3k1h5gLZoQQY
I82Pa8SpwBDkV41ifEMyH3eI+BzRyXQWYsmAhc0KSfRFn7PYDlVofRRJuGhpQlFLc8YnLze1UOtG
HuggmOx4Hf4eWeXNSMZUTdI45eSUIF3MsVc799tG/L/q/giwHaKE872zgyKaLhCNHq+2en3IELjg
kEwJ1NJZ5scaVgFdUjiT3UjNm4nZsSSH5/eb+UFbHZbdg/v7r/7o2uUxHYphrv1jccazUomxot6A
nih73xte0LkZ2aKoX/IEcMyHDgg47hYqFduU591ef40gutUkjf6iMRSvtDwzf4UJ10s97XvTXhOH
lhDLmsqoMm2E9bb2BIzGnISVGDqhP04U5JkCr/KMp7G8HrNQhCr3jwBEGrv+ndKKb4bvCieYNqEh
lwWIaFpBMvNgkSFiK2p1sC1XsRnJfyjbEsvAxqS2rILr+29isO1Fg4yhe1liz+aaFGEroOYH+RJV
SBNWve1fs4/jAJ3rLkZ22haUquflpB63E4hOuP/a/IBxyp+HdS0yvqbtMk/nor3VlRPLcyWGL77/
IYXHy0fXNbZ2sq/Ao3VJ7ZLM+lLLhwF+7ZN4oN/ZCjxXQw35zqMXpuFFwELzm4uQ20AATOYM8n0Y
kLGep+pmUK2iaRug3KgsmK9G+RMaHYNs4x3nXB5f9EeJydkkcbj6JeGEujgEIGPUAN9sjunRyeV/
uZRrpE9EFiV7ilyTaYXCBei/T3M32P2sSuoqbrW4KgQ7vw4A/nIMnzf3G58k7spRS60hIjCjRUGn
3Ey2w3p38VS8Tu3TZefIB4UJv3yZ9ift7VNepqbaXdLrEt4lpQhyWEUZ/Ak616JaVy4EVSXBL2ot
rbiH0llOymtyq+Po95ikvCG6CbvpnJdmkYdwlReKnCYCKwmOb0ndbe4RYPMBQWYPFOMH/RYkJHRe
KtQ7utCRdkVxcy57XENWdLj2PrxA54ZkjQOB1SD5tOC1A9cPohvVF2cwg+U6bFRSV1g39y5VGv6t
3BRL4jygCtLWlaT03mH/kOw71KMonl6BQdT5Ru3bqY6fZuEYil22DtgL4Wm6Le1zeQNL8ug4tLS1
KZX6v++JjZE8m3oDoGItKTDumdHprRsXzFCQqLGj0tl0vlNG+4AY9WVc+1CQZKQOAMRk2paX5l64
86kQGb1IFYOC3VL/kkiAwRaaHE3nOS9wtSuuD0GakMwKQVS6tKR7A9IFxuxcIh8CfCiKSu4PnE//
hA7KJU9nXsblEGuWj9ZDD5ENFe6uQOiYI9/SjPaZpAmq/PtOpBQr+da0bQV6u25Zr0dhwluZuRcl
dbzTwF0WJGNG2h5lCXO5gM5CAAJp9a8wERcnzfgKfrwkirVOrWmyR/D8BJckg+Ptvrbf5ve9/04b
aSowXzZLbT16gw2y3MwxP8PY1DH122Q55ZyEYaFzY++r8vzzCFhQTjzx+dfsCIF3nmYu9oYidQkd
JAd5k9MoZGgpA9FSGX0XaV7Ol9h1YII9zesES5smAaRYdF3QwvkQgZ2Z+VMy9Ooh6kQigt8Wvq86
Q7i6tza7/NdPQNdOEzX47rd9PuXhe9ydbXmwnx0NF2Iotj8bZTXRwOAV0vqLvBKTICj6zIN/Y0+3
pGdaq8rIAZeaLf69Gkbhc4kA1xPHs+5Duhb2r8NcpxENSAspfhYHowcg6DPojR/sDI+L0GbjQuFh
mbQ6JoBpYbWdrDoGvEPu2wNnBuAvAvVgy2iH7mr7QJB7Y0uWO5sYINsauTCltZ1Im5KsdScOr0Qt
yTwJ6iZ0I6geLVrMOjr+XaaChegKq5HBeGvAloByfRXpfFvnjliQG/RWJfhrwoKqdIGJ/tbv/7xR
zyo5wQDwmByBqijzwlodPSoIFHux4sE1+00XwQqUbVFlQip46lSMLFcQEpAHRwIpQWEmRyMm4u3s
3icpFK981gpRETix/lZXqMjQO35TQ2kjBmw/YiQ2YkMdntLh9Ofhd0AmZwsomG+s1SpeSwEX8KzA
DKA7qxuDcHkFA4kdne4Af2e0otEo3pohGEUqoKPGoYvuICQ8Zbn+dPkAk+n05pU3qF/uSe2W4A+g
NFupR1p4Uonhm4gxGP7CBCCELmd7prdcpGANOL37pHiD3jNl5QW299J+JAqEWEhVJw2pdLpbb3lT
Y70GlcPMqkJUaWxnMq+vD7W+DgA3I/tp/QjrswGe7pDSw6Nq7LV8aL+6FtiFB1OVdDb/O9IY6n7Z
bvy1pz9OFIAYiUd+EwZjeyUfmQ56NUc6GRZe387PxthcAY44O9Rg9PIY+mYJuF9wTXUoDxhN1VDI
+FtiDemlRfJ371ZV8mO0sJpGbjhRkJPyYkjOgPwUrv6nRPu8Y2+LNok1sAZ75RsX6zDXmiqdgrw8
NBAD3wXNzx8BjrQEM45U2iDAS454yjaR19M0X3gFsk3lym9aYfd8dNy7J7PFklvVWHl0PTUrSxfE
3DeF1ME9vx6hFeMK6XIb9GorYjfJaWjnP99OzSHJql+1Kmr52YZlp8MVCMn0HYoIxOyKBEpriOsm
xvBXl85DY1AxXMVwZOoNOxa8IIlhNhUMbZ9qEEy/O0niUl0PKyvmTo1bfIyzbp7jD3zqWGL7PSkn
gWWswGNJpaQyIFdd66FBCQvMUUK9XirNk/p4/XfhxrKqEOGngylPY8Y4otaW06q+87mDJC7q7RwJ
7aFIDZBfWrrHV0aBIHGAhdb3uiuhjESdMcz5xxdkfxiqJjFrBJE5DLiHoPvJHcdA+AHIvW3RdfZ1
ULWaAEcZElwHtL1Ui/mu5jtCQNU3uB0omOT3s0rxk+7awuekxs+hd4o3EtgO8grZ/ByzyhyiOuYD
gwbcfb43H4MW3kfYTdV/CFz2CoDdp7J9gP4c/299V//paYqCkaOi/W/aW5PIiOzkfJMvvdDZ2cPP
d9UMOUqgjTzC2esZDunf8YBZGrSUipYbv8fGsZCRZS9VSCABTTPtIa79P+DrF/HDtcqRpL4uFkjw
VQav/EszIRzhZQ6fJDh2m9WHyelJBlSg9u99K+l2sBRt3zM+VYU2jN8HkxyfyDSQp+tZE43GsWCE
Gv8treMefqRq4GUqjSSJNpYx2hZRf22zGYgMQ+KqYgFZiviMSUOepbhpFSqxogYcbZpNA7UysKbq
Ah0XTT5GEegRIzH2kH/BsNN+06njYa5Q1Nm8QQuWPdG4C8QWc6Oq/10/u+imZt/l74yxygmP8YrM
FrHjuCMD9x/L9RbhVdEY3/p872xSXSiidbv4W7kD9J6jtuBPTnUJfta6vYzI9b/zcZ0QREhUfjgV
6fZc8FTbcw7e1COHxK6jgNPxrLBjqub18uYQx2xfPRBe2m91qCL8A7A84mGx6FQKSN1JJSMnhlwD
jlPJt1YXNbSEybCf08xUTWeDDJLg8jdKUBfP86eq5GOuSAwXb49wUwxllUhf6VnuMuFLZzch2yDv
3e2Hf9Q1UrOlOrMOZ6oWQUrDfSAcXI1vqHQMbhGUp8K/ACsykG6ByseUvUCKShqDZo9DVcnQR93f
TX4khi7Kh17aF9CG3NNh4nGgc7wAJrIUcskjb6B3DjTBUB1ueGWdpbJSURZeYQJU349yPXVqtqBm
laJsBVo8TOxUdBXMvgqSzCz3IndfsFpZjmafCqKxGmkLx2oHlgPYzwdYzks+m/iCjYyC0F25LcxK
6RWSUF5BGwYhS/Wfk9Ren6+0LgyZrtGBrhgW85hzmzVY8/2cwh720uhKMd1yrhm8tKA+WX40tNf/
A29I+WlM7GKYALx/3r23iBh+W2g4044i1fGqhRCP8C1sBrm7rjMitwQ5nngBCCUwFCVt3fjsJQYG
blTyURhgSaS+vb7xDXBoeDpVXei+LRNQpn5JlUbaBIR6zesA3Fn18mk0uyvMnOVunNyrFAHK/7c0
hzQwejG50qaknaCRWwzoKee2Uf2PnHESSMAssDOmduhCS5B+g5BBwEincebVjoV4UrdM2rvOxgqF
y+VZmlDsHpAQqMEmtNk7b/0dhj6wCuANET0jQ4pkxI3F/CtKDbWqwLTXkI9aOVSQdhdjskCCw/1q
4OQhodnPLX81eTe0Ur714Q+WyBqdB7oblXuWliW+rMLxJ89Sv0HU5uH1WzS9it4PqqHNEFTvdAeg
v8Vgd37m6dvx/XMNPP3cHkgXE+UcaQkip9XZ+rtMe8C3Efoir9qYYe1ZgoSS9+fpxvWFxZfSjOqW
oR1uc5miCqAGxzaARZSqBPqwE+EWTZPXsOxfFbUE9Nvy1sK0lCj2L609rlMUjWCCaIJXXrQw/90A
C1qLNpcqRDM1uVz+/dE8aWVmfyE0hoef2KiRO80xXShDD13p7ChxgR2Cuk6wknbjRAiHtFfe4tNd
qG1kka9ySl5QPbeOklQP2H8PiXleI+RjPajOOe1uxGtYQWofrOAcgPy8f1IRUcshq7Qpk9gekEaI
Yfb3Y8DQsOjaIYO/u8FGZQiLrnCdz9RPEcBtiCnuUMoXnIw3cYEU+QXuGRdwyUdK6mv2BxsJU46U
RdydbkK0JWktGC9X+pwS+B3f1TFQtF99Sy87Dj6Pqny/1XyAaVBDrtL9qaBaDjrzbM5uvV3nT6K2
mW/K0icDasepY41PYJaqzGv2aDTQgSuklKFaIi1t9RNmd6qBqIfpKkigwnlxvEWqJcGM/ePYGOOF
UUltMAYlseN4TvIxnElo0x35t2QSYnv/ZQdYWOXCoBuqTND4VmjQNWPGXHIUFzfchRukzu1AJLKS
qcbz6Sb5kAIKuIs8YJ7JM/nrTE3gV+5LmxVdkOkq0bp2qDBfw6QAPau/iib2WsDb40dytBg6gait
p5Xgu3A0JSqWOCtSHSCZ/3h65g4XY4SlpQ5/zIYoeYAlfkWxv2mFtUy93GI4avON6s9I1S5epPlf
IIQTNfEuVbE7VDVG/dEwA10SMqo0cyY875jS/qcqlsC/YJfGS/hRwGpkSIBhwEa0ClAGUQb2JOT6
ryz4pLh/H2jUYzp9iCFPc/N5Cs6xOD4MxcXd0H6tVN7qaxS1Dan08kmPOo6R7pJ2NfselZAkq2v6
Xrkq2FFbrXRCQHk033t82iH/maYab1xmxWhULf9Gairb9qxeKVLDgw0+bbyGJ4YWd5dNJ4iy5Wy9
pjOjgPoXN9RZ1zwVkP05EO8n1GabXzU5jfUSSN0+ytZRS+9phHxWUp+ENbMiTpt5cN9y7fknbe8O
RC17QKaVb4fq2f9gacPzA5H18+MQeue/MgOUlJ41ATB1Qr8cJPXoGeeRgytERQJYoO39i8UbUvRp
3mekeKgP69atDlp3/B1LJBuwiZQSZYEP3bV+4Wm4/ANCg9QzBoK5Y3D81Sp9fUYLDa6GH1j3cTh/
rgItF19oe63DYAnUfBqTinbfy5fC17ooMnxmABKV0OSt715FuFkYVOwdmt+bbY0lHZDvReybu4nC
ZKnNMNY3RPzx0Ns0/ULQQrC78wlcdUpcq6OfBMAVJ2EuoETcS1HOdMIk10yvUviIsTs8+6sZ2pF1
37gU8rq504IPWxi+Q2XI7vZAv08bwqTDX4kTDFeldQVyxHT2cLgebjCndl61Q3hzMwd8DuTA0MQS
WxKpXD0Nzx0abIb0N49KQtbVT6R18nkr/J6zlaLNdCS6ETutYNgRObsgdMOzuvIuvKIMs1SJdDGW
VpDy9TmFmSplfAuL8zu1Ov3GgFB4Uddk4GnsktJdOSjNJiWWjpN+yOj7YArchpmjD3vKzE+YYGok
K6YF8QzqEnEjzYL1OvTmTizAiCboFI3oFSde+NKIL5v6VhfXZ3DQkCCj7YOWhE6XnI76mF97HqLr
qhg3uocYrGuhuKDq27VdG8g/LuZ+J0ml81T1/7LGmD/VL2hl60RL0lCJlMC7+lKcfOvsl7iq81JU
mpR2DD/+LAtH3fLbCUafm7QoZ4yMopj1DeuUF9shZpS3YtNHYEZjtInvfJuicu6r5r0fbBYODr/P
xv7Aj8Oc9Hgs94nGkysZzNch+OzLJShw0TGqA1F8mim8PgLhmDfbQSEOgi/fcARTNJEH+VZjGd+M
zI4Sw6opGydzdzmiZE/K2a7Cph6sUPF19k6qMxEsUPGRV/xKkWU8tAMZozvWKuPgGVzzvEL3wqAW
zNmBNSkDp7mlrZ+/v3S5/+VXSmSYwWGOuCxfw/lsGseD1ZQ9dTE6a/PszDjILSrtWrvP+OX+y4D0
c3rvoBBQ2YNqKA4LF5WuOWjWdjuDbfp/7pP6lLvkDczLLRTf1hL7QFtfJwcykD4PvIPkuUJZwYcu
DWGSi9QWIGE6xZYRE/wvUB74O+akjFzJhxoVEiG/Ej+HHIfKWIoalZnB9DjPlt0tw8PKddkRXyga
fXH/F0k89PU790D1KwE3yd/1k3SliGDGXBbiuEI+DNbGhawFfHc98mkTXKSKSGe6VTpYWgWH6X7k
ZyT5jIlP+9CGvWH6WOk4qt8RgHLJsOpUibZ31fnYkrsXFo2kG4n043x5SF/3RD1UhxEaYDvYS7fu
yPSK3EO/I6M5OGdlwGMMTYdRTOEUH0rWFhUd7hmfiOsKwrh/29Umc0qZxZ/TRPklJWCrGji0Lbvl
osLPp7+A0IdjZB4avqcTmwJOpOK4pyGB6JcrbJ5PGEAb9NmjN9aLdMl1FSfosTnKgKJqDBlKeNX5
vVeDe11/Nl5FJRwDVZs/TpPhPSiifmr8hVHwgWVW/WDs7QbzxWW8snHLuZWFMFTDJ2mpyu7S1FAt
ekcH98GNLCHkOWmmNaMw7hDt9/T3RLKMU81kRiGMKJjqf1bHl3OpGpqG7VjZoO9WdaG3qHK2aQPf
ttPiQGPPiwAUQbZeisSwTiuOYBbzgCCqwXKkgByjaojTIQfdB4lMB0y8mZViU549OrPNzTZ/8QGg
dZsS0hUtlQR3hC6qOgp1GV2V5vcu3HMVL5VaPm6glmMbQEGhJTLOvaq+jxAD1Uagde6hv0YTo+so
KsustuL5RZmTrX7ca5BM4OApaEK3W3zAMzdbG0W1+SFEYskH8kCD+T0t4ta/i4SggEPSmDJSNJvs
brwHFxiW4bQ+B+s110prK9hGEYGlfvcqYyaM3xr/3GuVK3a4bU8JHg75iDyjpY8i6v8iGnayGqKJ
KQZywrsUBJBQT2DajTVRpw7CMP0uwWVmFjzL1q9rQ01KjHrhOrRcdopEPcLv9cUCdGGNKunHOpt1
tgbA3TDHJ4RHACPfIOaSEb78rjq8ig3UdxHeiioL2FX2/TSCyKJYYPnZh/LHcNni9rCySYzpYurP
ToMEaPuUASG0az48kvLDFgUJYpuX62jd/lek6UAqQA54qFP0SdBtWJMsvBHlm6XiHWDhOPXt+3F/
NsaKVzibgEkqaf2TNqlCXBmlePrYnS+7tXdyOeVXRAMBkIgfmgEvCtydLKYampdTB2ShBpQKl9vM
U49evM+Cu0lbeEXybNrjsrXbWuRXQPy+OA+S9lVtHXaynx7JpJpneZv64vCTFiv89AVJw/TN26WE
V4KF04WZJ9ebCMnfcAvrNF4E4KAYn0meIAswHuHNIDUpHIoxXT/tRrTYJx0sHTcd5H4KW5pVIooC
COgOAp4AxuHseqUovQ2K8GMtW/naFarjFff+O4uxV+1ct2UJ5yvtDBURMrJTfUsOJdZkSXOYFg7q
EBZSTgVvk/BcPIvBRlGu4ke4rUO3SOGpE30kMjtFl/5uVVaE8lfEHOQJk/EEXysZOpmZbFFUf8NA
AUCAZEPv1n6rs4hJ5+c69cV3mCV0Vomm+xcys0vUyXyS43V8nHMhM8esNZPNUP4YMG40ze4EmpFA
rt21TgBd0KF6O5ogXkUb6QQNpNOb8RO6rzJVphzEE5mH5IX71ftmZeSudlNBNgr5T+5HwbbcXv+v
dRPHwF0aftnIbJY2+SLH5D55odMoU466kBQFiXafOBCyZQ6y/++B1ySPIdHKuWrOoSbHX///lxwW
dzsVWk2Hp4S3SR6AV9A2QFmWtvtndS5+nll3snUtHrLZ+XuLgCmFwqSmlUxE9Uw4ojSBXvt0u8ao
tBCJGFsJ+mTAwP0KyMV5mLJHilTG48ReKE8i3y+sEWhCTnRsciAJgIbrt+T59orn3njKJk26vwT3
loe/XIVnwtkPZi2ChBL2pbyWNFpFbr2OA8ZEvoCz4AR0HiulL9PCFnLSWsV1WsvaxexoNYHS0jL3
CeJxZJBX3oGi5XlAyMmQXRA401jkZ0IdqvCc+/zdax9mwDVBzKO59+q42H7/dJ29h5RM/gFSk2bS
JuY94r/d5IsqcJMvewk1+XbRzPDZNUxfzgUqFRFXrxxByk+8v00zegRytv2G6CyX1HHpd/PeoU8N
fTw+d3i+VH2q1eFHCvWsqkMXNeF6QPhCjIcIUYrnIzdj+C+btqMGX/8VLvMg1IdUW/9yVBzmWvhJ
fACCnfWqd3zyHOsBcEATxEMNtlAA6l3u1QlEj7vhVbtT2CaAqcd+Z/KYVoes54VhYiEFR7ZL8EGW
Oh3FJgcfBcrTqLkKIvruiOBVwI7c5I0MXgu2/gWuWu2u30hAlNodrWAU7ufmxpaRuxAiGwgxpQbc
FLJSOufh9fwOQXuVBFQhB/5xDEesnMuF/jrZWVctcflwHkJnkAZGTZ8UI5IgOKTWbxUz4xkxpur0
RoEiHXgh0IpNDdW7oWuyW1jpdFOmgE41FhtS1nMeOfLf2hV4y3bSmeY4Xm1Tz2ldHhlpVD6YdI9Z
oP9nl7JAMWG1b4mKywJYTZAN1/Vi5EKQYfe8jgU2kf1vBwLhQNOIc2Msm8jJ1mgm5DDRgXu+Baxm
I5SH1uP+QwTxalU3h0wexF7PPBuGo8N0BHXAiLyv0rk28ph4Xvzh0bvrG8HbLH6BEqcd2/DEOqov
OcbG+nbTc0ltXlV5v5meVY8UegJo89seMJjl5pvvcnxLudGCYj35dH8HdaNVkwUWxuJavoFg2hrX
WyTOBVvUSa46kocpscA7VXKMZv2R7ER4PsdUBiqT4WM7fx5y1dod4Slmfgx01YrPAJs6Tg9TUT/Y
azm/jIjMpr6viJ5tiquy9UywDwSzH4MkdpKZHu1631hdx+kVJJv21xbqT/RNjv4xRMvAaueZSqhs
+aqMZUx2Z3PQ35CTG7oiqUjjJifcVrd7XQS8cFYdf4nwExRmo3cgZZY+OpZT9amx+WRG3C5xX/TQ
Zpq2QSjycOBfjvibynIeLTC7C/ahYLH5ZhmZsuTPqV0pne5caJXb/6Ayh3juQusQugDKIMyFRHjo
0FUqZhsKEbCJF7+udkLyXwK6vesDYk4LnDhC/mcK8yHHsFTBqFMNi6PQMz/Rk5SXNC6qo0jXyXub
RnUQRSUWeJYPV4nnX/qmsISb3K0jJmXiez6FidQUAdA6SXlxHbXeRdwxgTEEicrYRbPHxdTcEgix
CVUyUcPU7+gaNlqIX93A1NZehk8ZzKtlf+6s0DrTnpti5eXYgMHnxVdLnY884BcWntKOUoDcmLu5
UWQT/ARUohfGauoIXDhAPBcdhaBiVtmwvQHKsJ0R26yZjD91nFH4aFMTduGOhTs3cq6SDIzryVLK
Jl2UyxAEeArgEeNzH2AJe6cYtszHdKqPu8rw9/kgApBEhKH8HdnPQWNnnj8Csfb3eZB3UIczpK7C
upS4fXPhx85980nrMxu7zQ0rz0ug6sWS4773qx4Sz6D5dv3t1HE9FBI0cJ+Goz8NiuLxrFA+M/fq
Y0SjnBcPRJIm2c9+MW/YhMsTI3YYTC/91SneiSraJYDUH4za+21bZSTSWslEzkRQRYBUNYabwR+P
snJnnAncEQlp8HBJHfz160evPX5CNmS6jzh5E9HIQwZUDIiXNhtSkepkmh3Oktr9d7DyalHEJOs9
pjQHRQTbs8dJRhb6Et6GwUHIng/rh9iLsTMlma42otINybBv04dcVjHfA9aFEG1hMTVLdhHEGpiT
14AZZyoDpDLes2xZtVH8MHG+UFgNlp3vnrBnvsBIJnqwaygECbE6XjEUcOYGjcDpBtzLsgUS0qx9
Gz9jYfr02Y1Xs5mBNI5rXY4viGZAAV42Do7/w0HjjkwzohgrLZqJhVTzK8kgtzNX+CaJXzA/7VZQ
zFZ/sofn04i9ih1V8NLcINHGrajSMg3mXIEKUNYJTv6cv6JJQcaTZ0JUyw2D8AC76/zojEFFSCEf
yLbQT7gFPWwGNYkWyxiuh+RXdqYRZ0MNTZzqKCyHHTNviaEO5DZd2XkYLJrnYWOhwPkXrO/xEiHU
PXfmCsrpPX5Hw9quoj4ExfJMvftNNamFYsBW8riDidjs4se/eIHkd/3jkL+pfkf8hiI9h5tekj7G
DKqXBjeKCXWzBTvqeN0dEBOZ/l0Hs+DBCralENZ3ldO0snU1eJpCMIjO8OMlB5bSZr+AnEo9vQGx
TV1eOKKDRKunLWxs2mtl/uRCT7PXMc4u4nZ6rVrETJRCzEoB5xc3vJmeXpvMlNdiSKAbUZ65g7mU
nRMewO3d/2x/al8VXUTuhMYvAK/eNCOJyeEfF194PstW6xeiyF63ygeW7HdyaiS0NVgQw+tdA0sd
c3kDDHH3IGLYnwaSt5Ph4MWgBAAc5LrYh87OEwci6SU3PFx8Wpz9dReEYM2RF6hy4vkEXtlx2RKx
9KyEONCTCqvqXBVx5eJb0FWHt2/Jm7MWwN8SDuRU+tJR7ILdLAkcK5RVTHC7zlQqwZ2d1CLRWG6Z
91aSsVHLGbJc4St+iP7YF+xezrnMrOQeYxESEN2pqLPhd+RSAqwHMahYg7fSNe7BrY3Ln3SP5aYr
TsavMsigCq/LPpSdzL9iRA9wLH6xOqZM8lF5mAJoRBnJ6s2vhacx4CeA8QZ59iFLt09L8gBwME1V
uGhLbe6fQQa6hVMRokFtFcTtUy/c/gq/AjeWoGwdTFG3LdZBz3SC2YW1vu7VlCVZd6a0T7WOrfum
//iO6kfUrBME+te/NrpZTDH7/8NnprpsffEhqxM55XzIdlN1ne5L6elLbYC2cPQ6hCWpeYnsppT7
tcv4S1AVOngawNxS10x4qxZcr1fT9WfHhuSwjfTz9JIiGJ8eOAKW/92hp4YjDfFfE6Umhhhuz/CT
KpS/tyUpajIcGYOdydMMfTR0vngU9lzAaGqX6rn08c84+Xgp4ejmddVV60P2V2OTLY+Taq+Pdw1I
H2sfFsKEF565z8jZ6Bp4S016fh3EV4mfUYri/HFKaAk65zYtkrORCaTJZzCnnxDdiv3EkIoOTSCm
xV+KkA5vFVKmm+VREWnqgvy2MXYiq+cCd1ggpLge9UTCoRXVfe6sy9PjjHntBIwvYhhqu6YDXxKz
n+VLE0ffpG8rwxPCKF9WlC7Lbkp5rjjckb5MW+zZuFa6f/is6V7JN7JW1lm5SPe3fmYFpb2p4/JX
1z0P/OPDzPgM5Asd2j3SW1gZHX1QWr6BS1BvRBukWunXJgMSFjaRd/R3roi2GdcT+9q3AYxJRVJa
MB3EgWv6MT58ZV8Qwn5pS3rllyNsppUyYaMoRq4Yox3k0mQCJoHYKJucbv2amiE9sgXNgXfVpx+0
85l1zF1mLnypYj+Y38Sa3DxKZ3kxseQEiRYl2O4abOVoVZOzK5Prr5LarfugYkUZCh6tRNm6sKUD
aUl0312RanGmFFEikBULl7K4imprnK9GPZNVfKBpquniA8+k9xXSbhH+PPk2Uiw64cM7jQrDWCk8
NjgbhqiDPOJHyU/oX+EyEp2bhpyLopUS+/nGsF856xmrMAEtHfEeVl4H9VdigjQ8zbnGL9CMfVwG
VGK/iD9Pby8VqsqKq3zPNbqafih78qGBOiMW4lr02jiKlRPfbv41o7ylaWX6FNYuQtSoSyU79hgk
4YJDf5fol4eM+ydA7h0mnzTIujxPUT3jBSWdOHqk20BYtzZGeoTIPvB9N78HiHQiNp3W9dP7Eze6
wRXQSUWZdJPTvuIhUh685IzFDdMboM5l2gLl3RljRTEkGUVfmVNxxgj85iQu93o2zrwcSDmGXISU
YYewJwdLh/Xo4qXmoSBKS5PCSgo92DxCGr8a9dHR/5yvi443E5JD0nki2O4G700gZJiALDL6r6cg
AvSgcv9RJwCC0KjFQFXREtnn+leTA94JVYT9Dr8NYdVxcp4tcfrH87xiH1Vrfuu29raP0BAFjW9z
Y/Pwf1iyMw6e/FDC7Xp9Kb2L0PFdjU4mPeVEXhb03gMIWBbyj1b5XujeLBC+Py4RhEiiKLDSUahD
s1RNKeIHPWrJM6EZ6y792r3PAcDFZb5BoFWZUpm0RTLDm2JQf920+78XYiQh+gAbD9oTpi2I4UXS
CNNHQDfGKI1q4v0ZjUIwUBqW7lSm2bT6qRpK1ANq3YR9e3wK9G7QKvAvwc6IjybO40NMUY9GOcNw
JEos1dYsNVhpA86ccMa1DAI5Mlvx+IqAUdHEgEeLRaNSjTeaUA1s+Sf//znHV1qoTYbzmZi+q6ge
EQ8cUpa7OhSKXW4Y/+r1IxGh6mJOoS7Mdzuww9fv3F5kw/mEQ0LKSk3fJswkzAJk6K0QAjyT3aa/
/jmIrgV2Ya/nM5QP8d7yAuW/EgqR3ICjx3eBPJOdPziPejYLiThMZEMwiASP51Wk/KvNO53Yg2Q5
M2qInp6plnVWEcYF2a/gR09BPpYxCWV2w2b3mVcMNRoYJw1AUgdk1QPgnxFqxxNQHXp3X0oIzBn4
4o66yrqfg98WBmH3p95CMaFbeDUefRfAunFtmjf1EaqjEWvB7naZ8uZaSYS7q3Q5AvylB+/VcrOs
vjaZ9XH02zoF34eap1nYE1QyYB+UttZsRsJ6/37jgj7PLYcxw/RekgiqfVErf/Onb9kM559MXo3g
OJcumR6OuLs15EMRwoMQwahU7McUD6iwQaMzltfWY8e36Qj6pOA29lUvp9eZ4Ob8GKSGx+ya9ofV
hQNkvhoZ+tOtx+2rsVfdfj/1W77qD/lLGu+CGT8aJLeLVIsNxK9gYDxYIrCiI3ayuvPdmpUzV132
AbgKwvkBi8knzbw9ASLiv7558c5D1hvU1+D3aizVLRIf5ox2DXv1IPA5n2cUUuA71R5Yu1KEU0YH
9/PLqZkkqJGaKuCZj0u5t30X0XcrLHsHxvZIZZiE3Ag9UVq8s0nbKKgdMoNvW3sNPu/aW1kXpU0N
zWTeU5Xb5nCOxzW7+IkibivgUPsfOxQTQoYHP2QUfSBXPZjahI/Qevys5KoYBRDUYOVBWx4fSRDE
Ugr0q4pf8A9Lgg5jnXYJG1cvvt1kO+Y0EBLRAuOOKTCticU+xX99NToujZ/f8DaPcNfWI+4hkg8h
w6IfL48dPp78myEvXy5zz8BBLhOgXQngUEChykrQXwZQ0jL3XscX9RycxeDqp27QJDiA5WsvR4u0
F7PW55jY1foDKq4gycdpZxz0zs21+1+Idzi/BL5mgOPKZc4TPQP3KC4L+mWmJlbdma3JTWfVeRFw
qVFiPmD/qALCo5SgHjTBD86PTh/Dqjm5pRU1s634vRDqlNgIDPgh/YRJynuR8V/Alm4hnp5/sQRG
6wLt/Ujq8jd9Tnf3Uewei9yRVbKTv9eH82hSCl3/Zv/RH0mSiyrEk1Jj65unyyNRd+vPdajruCs5
cskNdy2is8P2N8wuTJIvW46KDiVX5W9yksceTPRj1ixQC28m56KsYQ8tVg7+igEiuwBsi1SII0x4
hTVWVHBQjAxDawXhyJNQGo//GJjsTy3kqMqJBp4PzXhBa4xODMYSJ9vkaO24Z1jGhq7wkdh9twaQ
gDIlQ76BUbDaNzicNCvMkfB5Lgwz4QEsSdbTi8wiqI0fJB2UaBhqob9JRoTkoRP2u2GwIKwADyV5
1+k97SxMsuesvY/X7S681BEWuohwsRBoaFiKhaNeD1tg3rJ34Fx+iGZlz5+ti4IaZ7ZSODQNf6FN
rGgmCDyFipmRIoswnh/Ueq4e/yBE6pWqtdtMJVVZCDjec65b2cqlj2Apqj3AGepsds2jWcf+Khny
foXVML4mMWNcEhwfPCKCBHcw8KjjsO2bDLTeEvSLJAdCFjGClsF2nELqvTw4FsR1XM1BcGxtgywJ
tVxmFIt91cN1aULwKAG6rVsklQYMsvnDTqLiVVxtOSVPWe5bPS/FcIkYrQNMI8WT7hk9ja5x+AVF
w1P5X0xMaoKXdLXehN0TecJnzZVY5saTfH6P+6h9X4qx5nlXnMHQNJae1yeqVN2+PIdwOAifmd5k
toD2BMydz293rZRQ70i0awOdvruYruZlIZt/fFjMYyUgWVVeURwKsip20n56E0Xc09Bu4paqbDnl
La7EdCn7Fxvj1nvW72CFLqcwKvnZXAdcLY/c9IijC/0IJFzLoJPId+P4pnvNbht9XC4VlJ8AcXc6
B/XH5B6zsTTf3Lylo+qecJJ15jj+LAzaJIQ2wFKV794HH6XqtT/o04a7j9wd7BS5oxSoeLS/fWnE
RYmFILhzCvB5P4eoCp2STDL/Sq0bvsw+tIjL+15WizVn+BTNrDgU3Ze0KHgNOxEgqsf1qdP2ROFr
ibh7e0Usi5SHdM6L/A9P6NqkMB2r5eawuGiYXyr5xKSfqeqWHVSMt9iv/jaoItVMYsuQuJ8LBxZc
EePZAPtomjvcqULV2CsZqFzmtIL0Z9/NqHjQ/bw/lOTK4FhPaMl2EKOCnPIl1Yz0lCsG1kszIQZo
dj+P3jfVpb3xbYUAfdGWSnu74UHVFwRx4skzvUzLkundgIUAS/La/TYdbnaXMVWuXnSIB0ImCz6J
jogM1cIwxfP4VyMUyjwr+VA4/qrL89ar53xjuX+n7gnqKlR/x0KWlGO9LmT3uOb/TyDuyEELeJDq
AGKu0BkmiP8eKJbAF6Pfk/QirE/d1yMegUDB1nTJlu0UU8RwnHh6b9IoIpUoeCo2tC+alPeVzOHS
8tD6koWJDHhfLiOgQbhFxOMuyO5JSABAQKluNamV6Mp2X/jI1txGqAN90fp+Y/sCMqVaIIX7JDnv
NKo27k/g8S/w4Z2+SZ96f81AFmslJNnoGXhjQSN2TzV3oUgdZqPeKiyds7hAg6a6Ey7YiyppB89T
t0BYtLDAr/3op17aBChOQ7a4nFQIXu/r+bTmF7SuSVxW3v/v0MRJlNcooSUMF06Tx6PT8BtYSqag
qtEgYU547IYLGJfNjRg/Kb1M4DClhwamTVBKEWEC7VstqV/EDprp+CRd60ff3gp8ioTXXzu55iIS
eMZPBNOVRSnThvAqsstnsuTHnbzCTiNPsFiwz5t6fnhDSbcWUZJReTew6Gpes/vlOoKZxQYULAQJ
Nc96pNg8ngv2qASfomQfRksfWHRf0dmQ45E8l5wXt8fv/dUY8b1C5HLk5A+ecUDyefGhok5IIzDq
6dUF1A7jAGIUbEecgd5Y/4tqoFjFz0l2pRedwDiNxfrPd9U5HQ6llCgx1L8z2cdgQMS/1Z4Vv1/M
THmj5FJ7zBhqPefttH+ifRcGNdh9paA8tcP6MN/0ejVWjiUnnzb/baqq01ojTb+wCFH4pjW1Q4+z
7WksdQsQNy7DiT8PQtcCWgPyBqYAEQHsS2n+4zrsTw34axGdHoJmekf8fHcM/mPPAB0dBGIDckXY
+BJY9UmPg4YxhN1YTa3dsS7cUvMdbf6dQddPsX8ZjfnIUvkvM0eUcL8JbqWFuPDgQceAESiUa6DC
nQUAhyphj/m8UX0mrViJgTifFmsRkxntrMjxV18kwguUlkHaTGsVtEfsefD7xKgMLRVhyrmCM5Ys
+rwVDMDlRV04Qcgi7ST3X5FO55Z9jRecX20QDxVLbOKn68Fp7P+9d0/OeKaS9QT3S85d3cbDofr3
X6qjz2IMaWxgq+BmEwMKuWUQ/1Q0d06CDxRuZdo65vkt5gMxZU4N3mUWzgwrKhbg1n3fy19BuQNE
gbY75QbYSf6Tfd4tfHzdzii5R8HMSZBjFFFL5yg1LNP3lj/EDzPuVcM86RoG1Ye8sSOzOITBylo3
QifaOzSMK0YCvlVLYrnxm8Lua6Tsr1IX862TN1qgl6bYqJPko9zsyBuZN2TXo0hG2XeA4jHieC/L
SkayuTrPckGtbBy4saz8oslSerOoIb/k1bgw3CiK+A1FxFpqXatHTMphM9yOSghPidiTVUsG6QZQ
/o25qTenueCmUM27Gl5KplZhWQ0fHiLQ4yRkEbFKrLq5I96P/Cf4KWQDtoVF/riFksVx5IYd2WWF
GwE9ACUbfcDNS8g9ZzpGsFFiajrrgQgi9uFNNe8UzTpN/rmr3+npMN4/6lXQcCkuMM6j2S/oBAxU
uLdlJbkOQ0pK+S9CfVv4q0+KkfsEwpYZuhVt0a/7RZAm+s6OCphmLMIEQbnnnqo1tMPvNfH7Urh6
FGbVNDje4z6LBqte+9tuO/cKIa/he/Xz/dSGViiwE/BDLtBBC/eJTc/waJQHhBMTD2XJq7l9Uk2M
+vUBvbEP8FYSCZdma/IvziWYJHJNoZrgafIzGtkpIZiVRG62rAMV+c3E79f6199XneX4EsFBilkG
dJ+bg8ZFAfWSvWFeWrvbs6tXmF5bMAFNIeugY6AIfZNmnsBN3SmAzOyjwFua9mOANzajo+s+Mc6U
EBE9/SY6EFxYZwlVXoT3oNmxbsVE6uV3vcOc9lnBlS0bib3QL5zZiPlO2CdAuGuxftE2muWI7MLA
vrC1h6NG4udSDLFVnsNEKqbKkUnj+nkDobtRXqFrZZrnhXvusZJyPviyEsKg6axIJXj2d44tg9kx
fkCfB0TMXpIVLqChAZMunILvSvs2qyyqmXCGTo2rBDACJOgNVgVjguduPsrgPRJ+zbet8kQdRVpT
Spwsf9Dsgh7zr5O5LRR2zoqaMdf3CthOmqRF2j35/kVsaAm/s6wmB2I3t4FmXNdCZ6lxSdxjJ/h2
UbC9ZTQn0Jd/EgijmuUB7a5E3oYobBziTFOHXMau69fhh54ESyse9fJqwGeQWyehZe6MQ/5iKaN7
TtyS2DYevZHbin5iBCs6Nn7KsM0SvqXl/IAp+QbmDNzTSAYtGq6xjSN5Ojgfhrb2HNj9D2I1D5iz
wt0P3uCXaWT4vzF5au50r02Q7k+EU9gZxP6uriXO3ULJ+/1LBgfKzW4pkPAGXaVAvi2c4Gm/Eeho
On5IkciARbeAGEqC5P9AaLRggccgjksiZG+LDN8et9R9fcwm1EZV0W2dgFybyetYcuD5QQbpmdKW
FmtWCS/eavafk9JrItCl6kIRGPFmft9f6/ut9dAfQsUHfyUhqcN7dJrr8nDRkbiwqf6YIRli2OIY
icSOzk6VHHgxwpL4YaKX8Tz4KDZmdegjEV38VW6PMjkIAnJRwRqrL8Y8QxKXu4SI34oblvLz6LiE
v1Gkswe+u8okikKtt1YGjBtAMIVfFElgP/q1MhErb8g+rSc8riPviJEENW6e2RtY6V+FutYfkIhb
gHv2wDU/4vHAWAMdmxUdvQR8inuhgo7exePKYKFgj9gcFOpwZc+rkUNkldc7SFSfyrYzcEbku8Pw
pkPdO9S2DT8TahLyaS96eOy7XW/5dslvD6ThtZ1H9BCv3CiwJYCd5P/pr40f6HinwTaL7WeivkHa
fzn+pKIPnVlBiLw11fKib/YFc+7yT9+6qHmbtEOjyUTx6PxYRrpSuCYJIdJhGy3ZLhbqVpY/WWuB
y79ctlaUxMheeh495CVp3Zp/+0rdZpbR8E437fqJcccBUYJRwkulR0fJdlhiX+ht6S/26sGxyt/3
YVqGSqgmU9NobJLtHjsEKEBoN8pb2+/ujXBfRoosaFJCOxMvv1VsjhhzJ6lGEPPbFY/eDdfbFbB7
Npwzn36msFUhB1hckZRwEzh+vcKjCiJhrMOylAbGwBOSmmrStmp7x8yCQt2YlHgL1K1j8ZrdT9Yo
Z/82QBaxwb3JdvMr2rsyq+s6JBxBqrjrJoukVHDzcdeIQ9QbSHKWcZbUZ/H9VQJ+CjeEGLQrSLQR
EOhmEvHFDfRFx/xUcpv/I+pncYoFXWo+Mb2TrSWNfRd4WVcFdfAGJWPuUMVA61Go/aa1Wi8BKmRt
Lbnp3PME7om0WccjYILCDgG3J0p2AjAb0bXo7KH9Ks8P+2Pv5yZVptPdo7jFrqLhySH4hQnlw1b8
YfsDcNUfSewT1IPJNJNqF9ZWrqG6tV/7JzWdhhcNgb2FBhdt25LKCdkKHi0UmQyyzLfOW+gRVopv
cIU0xAFLvjTffw37RQv2RzMnDe8uKkDO+FRXiAVygZQtABh1Yje1VbVYudI9c4ccRcxB716VyD+V
r88gMtdgdCnjcZjfIjqMzMQPS3LOK0lo2iLEo/vQVkCSH6b3PzlJe3aPoElFjV6Eao89NFbyJAha
zByD+WSFj1971E1qQMyFpQXIphfyWpFTc7CzaEV2o9GYHBUypT8fB/6HBcRKZwHoSZKPujsjGK05
jZzKKE35U+XA9Irtgsw8ZDdGPqeoKdX1+3Bxoz2kJxbYaNqW09vjK6pjrjUcc3mLDefSc6II/Wsw
oL/FH092DV0zW5ed9pblYpG693dJirUs7k4FeUd5hF0qXP2qBrVlYlbMjwmLB3bsX/uMb039cYrH
ai/e2taBHAeB+1nwM0Roz0hh4UDthBugKR7VnTOKpMb687w1AtSHOBvPO9cbsbYCwpDFLsIPEMNl
m+kXKIbD2vCgaE+znWPG8pCICY1BDKfTBQ1D1cGhDV211GFqA3DZl7MD2cLXBwvWOcw2qwY5ir9D
Hw6xnBFOVDiJ/vgGiSpLSMyGo9owOeEWf3Fyg0S0WtbLTBtRy9e5D1HVHS2J9rsvJty0HwVqtim3
mfdjLLx/Q7zg9b0TMi55b5e+4H/aMBLNEykJkWsq72HETfWBNOcH+NQVjmEjSV1e8Wnj+3LUABOF
B/MnQbkJncc11ZwUnM3tFWhYYlQgQCia1zu4K7NpR6aI78dgy7+YfZj8xSPRngzQAevu52LNaXsb
KgL2dEWLzRO7gc3OoVo6ZeqVafiMP4pftKlHky1dsf6VYMRETcXbSKTfR/VKaQGL39FvVbHO+qBV
eA11AzrxZfNbwXx12ElE6qVQDGF7gAU/cwD9TLC06pN8xaIJd7tXpLp9xyfA7rbSuMYFcuOLHCCo
J3zNReewE4YIVJ8DRZrxsQeN9tBxT2ZCDT2GzT7PTpS08/+7M+VnbxIPlEeFlC+e2mT19wjd0OzL
Mtis+fJgbO71yxFOoVEQGcPG4wRlP37pHQ6oyDnjeawQ5iCVbJL8KFVd5N74Cah0BJL1S5Lnxx3X
SqZ9yE0XrscyUpM6mwhUdfPAxGMEOl1mdlPgBdQYCjD1GG0XGlSf56HXlE1thKhJE4JYqwd3t6N9
jHA3OIP0cchBhWo6UlDXZD6kJvy89CFbLBjouNObVSMCm3IH/8y/X6Ayu1NiLFxMHl3BGY0fFICV
4pFsWoK1Nm5hBJqw0nkAB3NbC5pS7yO5tir/3TPi92mL8LUTl0wrQApHWZiP3XC/XLb10s4a1JSJ
kxjOxVvJtNBzDmChbngbOykwZ2UiVD596EH45WSwvecUdda+qHyWqgwuCzLQ5ngU3M8N/bRWaHOj
PLuawAiELZWm36t0UElsosfFzaXeKa0j/ruqg3J9CFVqQigplhTc34hxSlnapnxrcocy+KaU+Il+
oFG7B8/pCLhRC4IWaWFU7HpiYhfKqR7V2DPSdjmNDeOZC2lu9yAmMG/NEFwXiBRIgYckmCUvfday
ehhV25aUqZzWrCmUMos8QgN7TYxSt8r8tXQ+8XzUL7tvGZ8sQHojPxK5BeGqu25EXtH1Qj39uxvm
k4QwEH1JbdgoDqcqaRmgTI8mD32l5h8UV4i5LCclACb8XLru9CdcEb0YlAPQh+f9L7nb0cUxbBBw
YbWakyPuWgx/mhztlWdcEMrdbvDN6xOEBIN+LHFuDYQuuanukAWDCpoI0KM3SdO5MgjWtP6Yu2eq
8erKbZmsZGRuAJ7BY4F0kKmJDs0rBq6EFM/UGIV6lAbVHpdJU2iFwpDD6LnJuS7yszEaqkSDtGXt
clldFax0vbwbQcrBk3Ca/pChnEwZHJJGUeXbnL2GhJowHK6gl9vEu/ARlFHMoNX/M/NBmRI8v6bY
zs8+KBhD4WgoxGmPBXXwo4wvYLaIwLA/vZXJwaHz6VA0YZnEQXmpVKZ7r2icfmXVA3FAsssnVgwn
5eodwoPjU2dE+BO/kmrSNvwl5NJxuuaaciGNndoheIWjTYrlGScHJuah8I2msIeJC483PJnXL/2z
kWpVxnuQsvB8i4qHFvoWYss3f6kCnVMJxZsSsKGefk/YDdfrNbnhishw/dkXdG9t9Cfl7uEhdA+n
VCIt9ysO6A/GvqdMWa1igDwb/Brh1+X2K2ZeDpJ+cH2NF2WNGGqnTqPmEr+Q9Oz4zmr6wC9y3TKV
VTih7548ssEneEc/ezJM3r7cU2rKgzLxW9MxYzps8wYouHDrAPiVaX7lItv+gfv923G7HxWlN4uF
IBXUzJwwyiL+gCh+oRvqAhn7oGsvA6kKG03G8oARL+byR2yblCQsaLBk3dCDPcD2scsI89y7khXa
2HtKSAoP1RFybDUg/gbNSn1KMTgTwRUFa0f7/JjekMa/FZH5cZypYBOtGH6tGbEKx8QoKSCM5AbN
oAZagAl3ueOdDCkVe7O/fZFN5W/kS3yVytapyF3WEP0bX7zAzKssLBv19tOBdpUhyJ6SbayRhgDU
Toy0B+uWoZEel3E2xMQPHZkH4SgPCgTv1JdHxU3lmt0PQStrjgZ1MI9ffp8qycVAj78Tyu+ew02y
yl1gxDq3CJvR4YY1x2W2uRa58G3rIpV7wrAjX+FUzuEhL/E2FSvK6XYpFLbWhD49VsdGlB0SQ6mM
tu184+4vD+YRwJBh2d0JNdSUl7uuy5Eh00ilRESCsS4nQCILOdgXkISOv/aK/3ana9I6K0xSVFbw
MPU7JkItH3TvyEQYJcRcgz54GH44oTAdRu1XHTiN51qlKKZgZjBmf9b1TZzpACYeBtuj6xrsTrsX
tImb8WhEVWWOxCVhvfARSpFAwlRkFcrlDrVZvp+vdB5v9f2UvT4JwiBh2VAB0EHQ0UaIzyUJxxLK
7rCaZYYF3BDTPKzDVguNJ60aVx15kxEWb0rVOI31uWaqFHJxGxZFLVgr476JleDjlhvAJHZ9ctf5
BRPABbT6xqCPT+ROclIYLsTlvg1nPYg1Thlq3R5PJJUikWVSz+l44I13io2aHzUxIr5pleNULWlR
8eCPIaadprI9KIVEzdFR4IHF0zQmbTCcj/oH2pFdo4YEOYv36TQYEPNH5/6PRSuoolnp1/D8qbc4
1XTC4DQZAPzcxFQMMF4Tp8CriWGKi1rQmBkGd5dUg8rRAIllRLjtN0hHc+PlKU6yoPIYISbnDksc
v4x6YBr90sZqyhiYNm+Uu44Zj052uffxi1hIYZ217bbHWju9L61WMtRB794ezjihYBFtk9uSmdXg
H5riVfD76UrTcWuKLF7TXg8ipV7SiU88/iyq87+fU2gIpPlzJGVpQA0B0O3dDi6sAuCf7sVSTpCO
qP2+k6C2ccXLsduaXPFANZmtjUFkkj7gfjuH/344vrkdoqGgsngA9ZzbKUxh8UxXEQ44rSdQ28Aq
CEu8NvWxH9N68t1u0KT93lxYxUYhOLK0q4NIbQXmpPdmawheRv+0liyKEmPhtFNA5T6nIspL6Vfl
1P3Fddlw/zqBbEu0yguYisafQ1dIgX8tO40QwQ6kzpCQXhAk6i5TH0b/H+VwFbYRMEaMyYUDaBzp
Lsu6dbGlyltju85VZLJ6NsRrrMxnWkDcgDPvjexIoQN9H2bTn+ySdqeIPG9ZCZ2uhaYnANsOQJbG
bwzDxzCyNFDDRBgh4jOMrC5Ti6HsmZHrCSy0B7vEZWDBQomqe9yk7h8bBeCCWrFS8ahCwE+88OSB
HRkMiT2//P3CTcBmUq17a6D+LQrB3lMad2T9WFSf3WzOG/IQRezG4KojzxaRoERmJRuzFexQ8990
x26YCybBTlfAquTupmKXGV0G1La941MTUvsQ1owJxjxX2GQ2YnTJOoMkTqhhMeC5FWsVlcGxy/va
uXYr3xxJ+eF2BBudrYlohXwbhLprdkb4K0MHaLSLsCMooWrhEtaH/6Vs8Yu4YBhGUysSdlGrw6om
5oM2xoVGdPy/GiQ2E+GsWNoSo27gLdf/i4lMpPG9ESUvUb8NExn9IDb6JHRIVamg88DAQcIDGn3n
ikwDflGxDq3qvQHgsEOjl7G1VrazH+I4VV+obcN95dO7bRk/Q/iG/1MzzVch2Gcg8uwLY0I/xlOL
YxJSaAdgQin538e4Ht3K410zmkVcgPBOtZexMB12FfjDOsKgb6katf1kTziIAizBiQdD7YR8Yf8x
o3j5xPg6QIOEZZ+4j1IzYJfUcruMI3ap4N3/ytYUD+yrfThzhtUXisiMYUKlFNt8MAcddyMfNEEy
50JV0K7uD/xcONbj+5xgYTqKyPUvmbTsHaL2I5EELg92Gs0DtZ5nr6f6z3KEu9YvuyFSXM+nEdhl
B5PcWsiHRDcm5FLJvqDOMB7r2TwjcCxHCIONAbEwnm/B7unOD5TyQLurRFb1yfESpmwFdAM5FNzo
S5GA56gpzQRSjVwfU5XX/KqhlVh/IIGtZwC7ogqYEYpZpBfPZo0vRLt2HMYJgphWkfjWzKDmWL2N
BqvlXRdOA5SH8XVZ6jh9TuOT2dbDrWIQ4NEuqG0RBk6XhCzvamxB5FRQpq3apepYe+4xW/2R7KXK
TVATW5nImi2cHxO4h1WCm+F9szbXxWoBvaSfuiWRWWvKahulfgfUQvZ3MQ0aGL9AZEpqv5b35QSP
Yqf1I45CI1m/qp6bHzN0mceCTuu4HegTVe5T8wKB+/hE5/mjYcWYXBBFQXewWmWsRDCDl/UnYyfi
i2IkNCKxpCaBFkSsUkmAvmZIReZdP5NvPsSP7hmgzXbETxcf/vB/UqwFCljcrOd/+KktyDCaRZL6
urSMHpyDRhbS0GUiP/8G/1hzRd74LeGOZizQ0jOzJ98Y7U66tfEHVfIcJ7UP/NEA6J0PAdDf9KrD
mEYAnhlWPqoeHWyD4nAk3WYiGoJNgRQJHgpS2MSTjmToCeF2cIrcNF1QGnLTX/yE7VAjNbS5jW6H
Z6DurZfB8s1sWL05GCklZ6dPlOSCZBun65rVe8Ui/2yCCzTYYt18MBt4FATC8HsNN20v1x4agPEA
P4jtBJKHHCxcR7gmTKJIcQq82D5l75QLUmn15qwR8qJE+UMEojvhc1u1/z5BaUL7uTr+lVWnvHCM
DRQeFQbuGy0cGjDvTI57d3fkOFORQ0yIBuwB95AijqE1baH0yaSnwwTTCKXfoj6C5WybcwQKLUrZ
ctKqmOMhUwK3IUHQg0HzaLznQ6zp2QKo2+KHSe51KxBPBxtRi4H3Ur8kkXz19owYC5h40Qgwdthw
/DrO4W1N6Yd/nXyXvt0Lxaiv7dhdnZcrWA2G+SUnkEneM1zY+7tDS6xUcaOsD+wz1IJj26wAJLy4
BRM3ufgBp0YBSCu3rRBrKhs/gxq20BjpLmGFQqCxZR/G2SNiiki9B6pjPs5tqnsEsvX+a15snXR/
YaBX/7a+dMPVK9js9uKWJmauXbjz3vZSSZS4Kd4+LX9tfLCZbsvhd9XRXIXm+CGsQJ/8YT0zRZA/
8DKN8xGP8lSiGvOU8MZ0pzH+sFn9iFsnZE3ZEB7u7gLJ+xD03bnV2rRb5A5KtbR9epRopydqIbMk
A5QvGT/mh7AOwAXYyBga3bdrmhmT+sYBaGmNwOmptjZTzb3tk8rVH/WwC00+WLpBHdgabzG7ORVC
51McHiYAxH7LLsLE/J/vaBvUh/DtSzXC+2MY5H5Y4cGcjSOmA7tzNQSdMjQrRw1ymsMDU40Q/qCg
tCFDslqNGiZD35PpOCukveM5SiAdm49wiHGCQDTHy4xihMIgTwMSawqHqd+dU0lzz8ydFzNNlxlq
6RC7kyGBNfMYGDG0Eycpbw9vsi3tBAFEz4CJNz8CME9YUlnk110kAbuN09H4N93WEIiiqpxkTbTZ
MA8hTj5kZ5doiwXrmqmlvaomX10tzmxjo2JpuSSY47GOjoau0HIM6ci5X+GlskAjlSwo5aujZ4IA
RDlS8NxtvAcRto+HugteWonhWK1NYTFjwjy0c4dW3hsJSobZCwGNKr9RxXtuso6wv17Ip2UZIFOd
Is7kHufdUSg3+4t+SXX4Cv7lgnTP6cmEG0qS47kVN27uGfB15oBE+P1ouxAoeYulWqC2DxPa1N8K
spdhGSKMqomxXaq1GJWtcZGeWbcVskltbLR519KX2QkJt2VAHgEr/eYOtBOSFTpIBnfxuKe0Jh23
b57dNWHpGWcTH9yLZ4BG+IidtZpUC8+jspm/dWIZEXH7PWNHsTwIGkuNRhlVH0BbQ2KxxdWUgLiD
ISxoCV7WWYXrnhypPQLI5QYXQR6XWeFowK9ac6GMhyONinQO8kFLfBr58vvFh0Wp48dFcjRmrwQq
RR0HPiHuQ0u99/rn94Knc2mYGmixqaaon3BtPixWKRZK5M0bMZa5DgE2ZHsB5TP2zyjxNk2x1bR1
ExqBhna2AGClodR1/IeY5y8ea4aLyhuc9HIv1yAYAWzK4+1kXASA04yw9rw6Fd6WyT73UOU5iOVl
wP9b1mIjctdcgSo4+sCHqe88UQfU67IgIcUyI8Z5Q01Ctfhlbw00COSFZv1dLAp5FbFxAio+9Aji
cM3Ov7NVIHi+wghgDojF1o/p257hg+dVQ3nqRX25sCX24mfunZQt+5t0p4YBe88nlWUWbj/4Hnst
euVJYZEcnR2PiGsSdMO+HSng5nN4NIkAzyqyxHRNfgebW1L5IoUAb5Nt1C8P+z39+AlwvQa4cgkz
4H1Y4WsoV2dSBf/toc+hzCPLSAuSzBwL5Hx/OEWNTn8ZVwDQ/RzU2e7HWG/5jl0TYYkswOqreK+6
xc72ZHIcVza3VfZOK6PTSt9JOKBqwEbX9caP0OUTppW09tTkz/+EK/9FNz69HMdbLHhH5pxS7euI
40fG6zxorQJFeBDWDJA1aymr/9m7vH8tNfNuCkMNEYMjbD0o6Z5hS0kAD30A17mLr929tjLfxjWy
OPAlo5ztitELc/B3r5G5PTNuzcOfpO1E1s2gnwQJG3QXj8ECb++md57kI2Wde9AdghGkY5PvdSp4
MYDJNtXAQORCyxF2cuDLElD33qshG3SBJH5rG3MABqPg9efjirm7+c3U0Dn8LzyuwP0yZcwJc3qj
Bl27WpBWpwlS9HNcaxHsSZ/isLAndhN0NjqSkjDUSRxs/Hfxd67dVbVK0D+jDGDLmh8q35VIMZXe
699zIPQbJozrM94vsWkSz7p9CuFOIhQ2JT6KtnR/wfUwdfGDbevphIpWzUQYQ5v0KcYxOfg4i+JT
D2fiTasVpk5mpVJ7zLmu617POz7mOynQKMqm9T2hKQOJUxkiZNV56ylvq4p5WX/+fGUQdti9ELzy
nMu0xmtO4lopLtHtHe3xGVG65wh0jEX3kWTxaimznLDNjCYMIXEX0aQs7JSHB8htKPpDl35vDkUz
KC8OgYxN5wh/2G0Q3qLruONtscJuIkegvJtQGWvvzkvx8Xc/0tFxBpi6KzGNPiZI5fhlIQniKMQl
6q1KJT7zPpyIOfia6WfokoYFtdvpYoL2oAdcldAKdUsuOLLFm2ey9Hzq9PCndKxc5q3qegf0F4/4
yx00XI5wTy0WpcJ06ZsYJOjltYCoq1aVnVqSAuNNnwccAs+21HRoskhc2r3c2iGSjCz6q151qw9q
uA2lx0yp8809W1yzZ/K/mfHZ4iFBmS03Xo1L7yM4NY7m/K29sxlrZpqZq8ReWhy6I+/LNm1gzxol
xNt4VMbuWCjwn7PsrZv5gW/EPwqP2cB4pohADbnbqne/peaw5g1cR6dMXZMDl/6P9Yt+xdxrDOiJ
PtGrgdkzJGp77nHhaYxiexO1QFqsknMYvpdmmo5oNCYYcoaOz2XaEvHIWg0ciBhpF5zuEqnolfYp
2Fr3tGAhRgj5fktBl1ydRO1eYs6Qv15LBYLDzzrmL16Bfy0Y41RDQp/A8I2nLjVE7t7gs68Gp9sD
Tax0VkQLDjhIyHUz3uDK+hwJ+aJr0zx1vMQKQq5iSTCt83023LSZraJUCBJ+ugemBqYnlQRraWy7
9arXd8oqihfhbay3FhY5OTiNYnnSjeDn3R3HRYSr411OGDVYhotljCTYDEcXfkxmSO1YW2E1isk8
v7A1Ul795VqEChiKtxLXLk4ZzBQXvvQGxyjMb5osan6ZZ8W2F3rDNYAQ5zKqYe27XcOwhahYsd/S
wYl6Sd81JwmRUenYnLFTeE2MLnA6tYwJNjicNAZcwkVaMBENkHd7q/YnuOnc7OBZ0LUy7M3iE6hD
QoObXK48EeYohLdyyVNU1BLok+92v1E7hkUsmr9+kZIY+tp1gMZneI2CR0ZQU7Rj3lZ+X5LIPC89
XtjQ4lrGejdIjTRot+yW9CB+aHv9V+pZUSINfKFwrO0d4gUNHW+BwADCc1VswrNkI7BuJmeQe+g6
XsPGqOYHsBKLV1SGdLLlrg9YXTmkqaFrkZIl/J/Goic7salgXrXLXelHVBFixr/VJArdupNQgEyG
hprf2d789gBm31MiSmWy1Yoj7OTTBL17kdVDv9ZEeEKNh7PtDqx4JCM2cKZfVGJcOXr9kN3mAM5B
XAsjvd94F2fm5CWSCRdbaW/0Tv31YzsRg5PhDenAmiEd9ZjHl0vX8rmfCWTcmoj75MHaRwim3EUY
K51x8R+itw14bOZPN0OZ8/O2H0qNYOv2ubbjSg6b702z7S8oWS/2oeSSKuHbjwnSXSscNR3w0OiT
ztxOLzr7gExnPLLxTx7TRdz2LT5FCbqlqErjI+eBJCjtkQije5sq5Uxn/z5OZDyCuuNkdpzUPdvJ
xKcodH3LhpbkbJ8kDDd+qXS6IqP0XgPHUhMqtBlVp7g3s6aR+eocZvgora3bKdqyuEqyf8K4J6pb
U26ODvBIyM8ItP6RbQ1DlK0Y8uf2qvSQClT1LJpdR9KF0/CV18nO4b7MTjGMB0ynlqOOOi5M65/V
jtp0rn9EbesE85cwT4VIB3KE52qWHhx/YcZ2xwKaIDhZ1POsg/QV5DHKGPG6NKP/FwrvroqrT1C8
6WfPv5F10aPmGLhLOWfPz6LgSKWHvTPVMjfEmr8DEtOiXzrXtgTQN+MA+TYqUrBXnpLN+fuZ//a6
DMkBK2XRb+HrPS8Fw/nqGzkfPtD5EyZItixOO6CAwdGoGgVb1OtEN8ltERqYHSWjJYzwcRvmHN0d
e6v7hskVEQ6rSHhRXj4ttQDNbY+UyuzJRrZKmzus2SWt1PCMiS4QSjj05ZO4Wt2+roYoabwwjw+I
6QLdQn+hd37zefjhhnQuqickCdb5LaMhFqYDDVpY4Cgt6Xyvkc/mymB/UBrCgyFDbq8viWawps/m
XFbPC/HJyPCrWoV9LdgGy795Fyi5K8WXSO9Kr4bG7L3aUu6KXkRuAmTK02VbAERYuv2BMl9RNZDJ
IGDpRpmkilF6paSv1BmO0D7rUnQN+vqx0nX8mWQun/yU6WTWzwxFD8zseGYHQ0wztK3mJiSLNhvJ
FIZFfPSdjGTSW4am9CbHHeiS5CGG9RYs08Opt6szX+KO47Bi1UCYvNdL29vRrz2bhxjPsn4Q0/Cp
rMklSaCz2ZBD5gXQ2F3PTiFIhWG/wS1pMSwUaR4cUSzFTGRAFMvbda66hPd/pdd/A1QD2Qbyg/AS
FSBtUJAIruGpuyIxXmNmuSTG6kywHBadxA8zMdJdOTjBovmSpnt0C8lw7Sw9hggY0VPPHhTxjUBk
NOSbdGJx1KfbUHnh+zPEPeVWlTzQ+9wJETSDdRuCUStWWugIuMluSIbQOhHLKL5vUwPYhpIYSA3C
JkWk6a3zEpqlL1R/EfI2brigq2gvXCkKEJd9u+zzJiqG2iAkjsyzbsKgwtwLMB0HbYxAM+J4dz1V
hyyBbC9F9WwXsQNVBmFRCp3COvdtAaWKoNditXIDf6R+Eaq+985EnJzx3eKaQVysbkt54PCypZbI
uGJAB4KI/uNm1IycThY4gxdA/3Hw28VCCaccTx9rVpfjsBfK9S2l3gVToWuichruXWca12i9VwCU
EIrbF0UMzOVHng0AG7LKQ02BHsdBDz0papjNucY8bASssnf/AxaUSNZen34q5hgqwm9WXOUJUjZm
jC+mxapvJXk18X+79hgqsmxkJnYk5KrWQyoREqGGx3wr823+WK/KWUzTddXY2jl8teda1+kOx1Bk
msy7B8jl4rKbOmb5uO/LNepTmgFAY9ZktVWdOD2BKYjVMP2fszJoBgylOYbYllCIctkOBjxvsLYe
TxyY6SOAOPPdtwd7ztVD7VazQix1CCxnHabV2QVH9nesQiQ5+zZPA0UpIlGp9EBAfv5Fb/e09hUE
PwYDcyhLInLI8mQfSQvdSBTCmgO6UKr4DCi2TIDaUjbEbwI37Fm+iDXN5hX63IEKQpUqcOvPZ7vG
zWJ9m8Zs4z7nUSouxBX/uuyBcAamWHUmHa8jLebHiiNgN7F7TcGE9+VvlegbEeWyfimZtrxcHLG5
mB65um4TRLtaiIvJoKDRRjNJK/UTa6tUmnaipUmCRUfIrhETg855X/dVw4XclT5qJeXtTAE/8RUs
Gv/OBChrx+eNQWglq4RF8KsazhfdWNrgUfhHoDZpMP+wzH0fFPItSM8jtlT23IaSACagkCC2+lBj
8JLaWinxNT5a+tZE0y+k1GUzH9amm7uVmHySSQVs/NUy7XofFmQv2PepAH9mYwIJlkYRcMUBtgCy
uY8Np25s+zjLAHZVSTl4grUsAiz8hpR3+mahJ06xJ7WuOZSR+WjXcmzK2B4wn8lNfxf936BP6yeE
dohFidX7b4swLe4rNHZJ+U8VuSw2ayyd4+MzS6R+CXmV4SOQYWzmkj7XYk8dOAIBRcou8/0b/gOI
jOu98JrUy7NnbVorbR+I+3lhaEhRrqYDTbEKj6KnqFnCYLxP9QtL3awWuOcgu58GxNiG5m55VTyq
DQkTtfqGPE8ggYCPJnfwKiqzB5NOUMAPrwvgC2roZDGAFgDxTmWKBHd7NG4pYfv7RGTtuenokxgb
GopR03KHXKlgeqmfh/C6f2dNP7Pc9MXjASA1L8601cm74f2X/vmvEhuolM2qDniUI1Ri7Rk5vE5X
SwPtLPzclnRb6QrZwlE9yP/ZYeDcSn/jFAl582ohMl36AdbVPj3zZN2kEfhsokBe2OF/gkpMHNrm
qqMqi55dbGeYzK2rRIedF2yXkI2apXxiSP0gdDRno+gsVWRA5blmTiWUE48U25gTYhUtv9tirAQb
lf/Puo+65TfcfjeCpPfP3IPUflrNPpxFbkajV0Xn3jzpu23y/Kb9MW0f56IscjuKNVuVLkhzz2RX
wpvTxTRPM52knPILoHl5/xJ76MtMrqoX4Z9jYoFFkGaf95Kd2oxA9HPCjyiP+6LncHYk/Ql1ooRY
JBzCXjn1Zdr6hE68y9rnE+xiI/mZu0kYoU94paYVUCbjgKVj7s7u96tUdFGAVUGO6bNO0kz+tYQi
Cefvp3nzvC2k9Krktk9+Lz9QjduHpYXuQktpwsGob6hP1NWb2hnSYSmNwFt+oZNpco8aafHllkEc
ltK9iQiiwUJ8V4Sr1Zv9ACmmTF4QKPjCgmwcj7G+wWElYSd4S949DEaApiG7xBGyO5+zVHmpWmO1
hOR0vc8iid33O/qaXFGaryNMwY+GcVVqw23qcTMTH5OeIVvunlUPDLWSFMK0/I+kISDZH6SSaI12
vlzyvp0Co8XA6H4Px4yciqGoG81+fuD7xWPjj0RrsF2auIKR222RUfimXurlqsC6pHBQNn0dwn8e
GLtYo+mzZFzWJ6ihOpg91YaPeqAdoJqnWT5L/7kSYE3f7HLk9gvuoiWmEpYIfxILtwvMcKN2D1lm
LWfGcUB6nH5wlxTEUDt/4RUOswQjJ+opmWnXarxrtZ66nBGRFSZsQEQaFSDc7M61zlZzefIkSwtD
mqJlgvadl3QkDUpyCnhc8jRzbWgJHWQ3TIinfIuPvIh0VO+fG+yeQ1uKQOHS09l4FoT2GhqTAe2z
llmkXaj+/wZQpjzyDQy+hlkCT0dqAxTBpiqopdGgRI7ZsGyaYU9OL87qT/ycpPMcYNruJQyqrJlF
0csuctTUxY3t/FnUyWq+WImoA2kSl6EVvou6i9Hgfb7HI81+p27Xu/U41ytVblFA4wtiV9D/yKVj
/NFoHJjc9nywrKvzXtCrrEJ1PlF8Tjznt7rUEmmeGlvStUbxMZXhOkOLBEJmUOf1VgCirq28Elfb
sJ8C3xYnHcTEOuKjrY+EfzxXJIY/XdenFjp+Ptm6A1pe4FryptAPo7IR76wH32Gr2w3NrQlUNye4
qFg6/FBL+O7MwnABUHrjDCGkRt8AfMWOgdOUurxhNvku4mhAyDa2RX33gHEvobFKLQOPenj+5Pdu
cLnW2MGMnGFQgcRI14WjS8efUHf8J+UqcPxGA3tI75MT2+aAjH7jJkGPc5w9WcYW2u/yj05J96fS
94iPR0oKqoiJKhJqSRj4BvtUXAyPg28mV+DPF9m5ZDdSG67z19O0CVoWd8RqV0hdir9VcTkKdI3+
6XEXwNRQKrolzLANwOt3nCZSXku579ldOginMTdT9/T2fm0/TmyQKtM3GIHE/lRsNtcIz159c9On
QGgO5VFvC9qKwq4ZaSCLwgyE0XDRS73NzQbBkEx/+mZNqsNfue7dFppn4w2DHbYVwcsUvHNvkKAs
2qrQnzXSvstbFxx9HVFRD+tyNpbLJjhRKXGKriDgt3hfZmpOAZiouO8RH+gvChSEa3tTyysJh6y0
AmP6jaUMejiSprY7XLCiHUlmjE68rQAiuHp8/EM08wNEmn0RPxBEBFoKQC+Tun9uXujWxn6RaEgn
uEXJhTnM/OwBFOwxDOp5Bwmk2mrw04581n9ulZae/y65HVlodQGBqMeAt4yzOYcaPEAk3WGDTQY2
P9/zt7q5HQ0i7EZumydWE0e/EqCdoKXiPBDi90xwitYHONr04HjQLO1HNVVZs2TwGjbFkNuopi74
/nLTMpqzMK8Vm/aUrWVN0mWgDXRYqdVYBJ7NtRsomesrvzFijgqCIzffIo+4xff62oJtmbhXMDe9
lAx/tyFDeWuJLEHR/yjDcDoXUZZXkwMNlkR3wp15iMkh75FDqSFvkJXGR7t5h1y6CB9uLgh8RihV
Ys+i1ggeiIKBtundno+WzsDQ93n/D5NbDVc+UiJUiQMqncLkfWrUdWoa4S2JMjJeGT0OAD9+EKcH
DJuK8XIF07e5zMFmqtUEFwzCkMVoAP1RgIbNNoo+2mhj/K+iS8BWHSj9Roqx3BDdDkijyhbisD8G
nwVYkr+6IggPNx/BHOyn7LttTdjVM09Cxm39/0Cs57aLf6c7OpJ41KaE8/pxsaJY9HCU5JpCH9VK
C0ML5fAd6O2Wf011NVMSrihRJ/SsnA0O62n3pcaE3DUmok64vLlzs6XKwXIyds76lME1f63+gfB+
wmCOlTKCPi9vqo8mW9Beu/xx6wd/dc2ep5tdeg7geHAafNfIdyXUtPJ/JKM9FEF6Jl33dDWmBC7f
15n7WX1mc8/AXZligbrgdbifWquEnDasFYpBP/aARUhOuRpHZnEfl/ZqCSPiJxDznrZFbz3ABKKe
dhxJRB4Ub12WoOKSEXhjQZzQgNucrU9hBKj+k5QiRkKx/SXRB7FszzIvUB/XlBxblgM7QBK00MFk
jtBUDbz0bPRyyEgPyb9n4+koKgGC2RLZPXjXSsZPUauXv9AnMyQo4C/QXqxe9vtvl50Zg6y5yfHP
EbDJ25WUTc5tYk6UE7CefxeBLoxbDmrUQi1dRDW6pU0F6XRN+3uyYCW9gCp6OZo0tgqGQ7F1ZPM/
s94o8ow3gTP3YtYk/LH6iP7iQAPaC3dNAWfrEAeQMVCP4BUtp4fh7v0kjIR/r5tp/GIiRHwtuMWp
KwID2P2WsrFFlO4b0z0+K2itUxMiht6eMGNxfV4wgyG6bCCoX6cnVVxqXGZ0+LwZ4MqUJbQmFswl
+qMz/XCs9VhnCFQ/KAW0EBYMDJKqthqa7xpCI8gG1bi57MC0gNpf0G/WhQqF2qyHTYWZdlugzqtD
79rFAYoyZobLBYF8H35wPH0NDdv55blnl2TufihDOJrVJAEuWAfgyfE3GtNj2goRHvAmgZoZBaCo
IGKYgtuXd56iT0hydW0zw584Pa3z86xfar2gIU19RU0XYGweuonMGp1aTAW3qyKvovtuG3CSsEtl
7dt7BNlRruF+Q8NobBqLXIuYmYH7LZoKG7QkFB0gf8+LOTDjsRvnra1f+LNB0XbGuYtZXNSepiWb
BqCXipibdhNLF4fxxCYtinIhehAwWKmbtouMTUj/kvs7RWey0FhwJvSNv1ZNovDTPgGEhMIYITae
+ZvyFSPBHPAuvVujKjk/UcWgvAeCz4GoDYphhA5Ecae4QRhMJsLSdWMRyYdKy1aqOsIA1iuK/xLH
MX1Il1Wb+bz4ZIillASFTsJtXJlt5H/wcXwQSgooF7RH8C9ODUzlyoaAPQkeh4ggLT0KP1HCJhMn
be4q8CkizitcFfcX9iFP04IWdLneruP330TNRDxAAsCGCZ/FvN9s3JViz1HY8EmzULjlt5Yv4C/Y
U0llp0jqa1fE8K0FXQgUGjU2F5tBS/k1jPWYdOIAuNWAkvOHYZHqhmmwHG6BReavjwNYyjgPR3Wn
eJ0FzLWj0nH1nlIcq9dTDEGMxUrvCwhvJ24EUREj10uXLRnl1iW2UohxHpaTZiGlpKWXNGwX3rcT
d9ghFZjUAfwU06jQyc4Y6edO3PqahDeQ1cTXuy7ibJgMDWSLFSW1otr6IZndnIh85cTRVu9xJ/9m
U252P1pW9ceC27KaEctL0hAcwqq7JdIKZcStH/OCqQsmqpnUx+ldsnrY3E706Ynl+aydirTY9G5s
coDaJbvwFBNdFmdbGLFYb2jqJcNcWTsCEut6UssLNxBzvuWQpss211Sdb1hH0EsSk3RCTicB0w+Q
r8yAyrOAd0ucodB0KUZior89XL6Q6P0LVX9Levm1mhKjq38/STIOmFnFw+swTZedN9pnaDc/3hMC
/ssL75E2zZD7No8k+8idqlg9b6qRx/xGoF0fs2bE3yPZWgh3teRuBeBkoSonp1Ku35Etn/k0ZYKA
zMd1Q+0n+pryToKCbuSEDBASKdVHyMrpynyrJq8QI5w3TpIUy7G9Yreg43GiK0Eo/jJkKJyjykMm
ZA8K7MCebWemNjSLahySfYuGOIPoIZKQbSPg8JptVcVOrW1bQfC+uHWQaAJSwOqO9y43kRLw2qYT
vX/Jp7VRHiFkv1AjkOJzp7U9RQWNtbVNjHbborif9g0CfF8TyXIKJHQXa30/XTUaLhYmWWVwhEP5
+aaZ/XGRt3txxVtjGcWu1/TiHvWy7pHOzkXNrMMpWdEyUlOmmxspDmeOWVJPx6xe+vYK3SoQzQ7s
cMttm+CGE1U/Zhi/t2teg8dHwtsqmvuGSkF07y/0uBVNgUVTjKKT+W0zRTmHBnLvW0ssGryBh5b3
HQvNoWvbV2rNi9IDDOZ6nBLRb3LAQBxkSjN3gG2qo1LLzLG/3lXi2Totwr7LtfTi9ANslSJze3gG
3plKJnVHstNdJjWp6NN7L7rAU30Y+bCPBc9GlmmDFd01iue5cD7kuMqgxpgmEcEdPU6pY/Jstpkf
eoaTaeGeVg+2y0CRcbLqyZP6VHjH2XJLg3SXKC/JUyLdT48BtGRS66+/j7VwC/bDXKiS/33qrZpc
i3gqqwu8+byJVNH2+9f2xns8C35NH+Na8OlaiH5bZOkCQ95OSWct1/vr0lYy3Tq63JqEYqAgNsC0
8tId+MhN4txYPpTD/KWOV50Qbn0FRIxd2UISr7D/SAj832G8taCnZ20gGFU1ueKCVskYL/tBlEq+
FVA4IURbBbmJ2Ps21cAUDE9NqMjHNumV5VZ4FjiQ6O9R2n/Z0VEORK1+Id/EQCDYmlTk7JkA7rwP
iUntmqNVEATyzfkdCoCm1l19Tii4/ZxACTkE4D+TXyXOh9eyoYlJvtSZhNXuMrqYMtNY8U7ZWuRw
v1aGR19Ajt2uJBN/4KF+IkcJIQW3m+uxkMURZDGCRDeHZLhHy7a28RrU1KRjT/XI3vH63myjLZuC
EPzI4QhjRAOwrMR23UjfnQvT9DzvORJyXVFRlYkmpx+FGqvBKe6ZYqgfbSOwaTAHgXXAV0VPj+JO
ZvShIemYv1aXzV9/N5ChrRLC7YF+OiKVG0le2CawrmTVPGgizvHtTX4vAP6ZQxJBoAjI5ff0DFBy
0nVwmeOYTgNcSEK7yoiC+13wi9tiPvK8mN0VXFv1HxPaPp80z3UlxeQg+7BiZA5Lw9I466jrXosp
OEzs5xhnDkFKWUm3f/dtMEhvUwSSOWOpFzZJLma0/Ls0rWPYm7ehgTF8tq+Mr0fR5mQ5eeFW0kdE
BePSo7grm/rWkAPidVY18qqkc1aQcUcu9+jXPZY6oRDh4s5de8cS0s5wsm1rc1QTkSN+eiNeJZ8g
KIm4Pzz+wesIlpg60pAbaOysOnqwbbdD6i+JVV/vxpkNaCt017hCcaF6OtgpN/cNTKuDlGtVi6JT
YH0LL8w3qbAEsShxoA1KNjVC5yj9mlkY/bFkuapbfDgUO0gYnpU53JbjPJncuhMxOXRqUZNMBEw7
k0bkvl/3u6aS2AeQs/4kZKjuiKVjtxNBaOnefm/NxPCpjMcQ94YTSyvMTcV5QYYLYPHL7zWO8KfD
oPp2dHVc/SWflD96WET5eZ6ub0BMe3eAVuLAh1/5DPXO0dOHY2DwSHkQivwQ4hzE8uKLJffswLRP
QymstKkb01yVHBIjtsUhwfJUPuDw6gAB5tES2OuwZx1cSzbATLvkJ0IhIpw/kOhbp2pp7xnUD2O6
VMBNY9xkKtuAbJ1Lv8n4stYK9lQE8zFinpxAph8tyEvEphrS9IlSjwSr+Ye4gqyUZHeES4wh8zZO
Biuxe3RYncb36Dwd/o8hT+1mFTuqt0Z0s81ys53I+PtN6DWBFBkEULt2eH8aoOtz5HCBKMtN5+u/
hiLawb2QJ2sEexAdHsT3uRJUrmkmSKozCMNFsq4Q5e2qVIh88TR6D8/9F/2Jt85qFeoZ2SdFsSiw
9sB9aF7OgnIVqIH2xwplVri5vQHslTUAZN5E4o2TFTKGlzqy2i+hzxNQWl5DGoLOdd0qz6U4tTdu
8oVDk+/5afZfJSUWX3kybQv20VyEjrAaAsfEH3io6WiYnA3NaS155kt3UePEwWuRCCfIoS+7IY/n
IxYtxAwPE63l+ZI+k+mpptWyKWim63dcWDpFUYW4SI6CnDELuvzcgcFTgtNuPTsKNDnD6Ion0NBG
TKG5neosW222DWSUNF4y3hHSSRvByUYPgSnwMHQlqCESnl6c7T+qKdKUK3hJpadVzlfd5UoFY3cj
tFv9y8nwilGBi3Q6YXOW+9HPp7c6uR1FDsONAc5h3NxGcCeDOcBJWP6Z/sHWxkFiPgIvwZXjEVvF
GxKy26faEyR7D5nz6xDG9OgruGHuIUvSJJ5CSXac0frknh4bLbmBpDmGARpHZkYw1vARsWKSBZAL
4pbSqPqjW3QKYCdeKTJDzTm+C0Wq6KucHSoyBe4xX3GxTHU2sm44flpzwC5itSFoG/QJi9vTefNV
qt0Uyw+vO4aIFRVxz7o74+620f8EDXbafbcjG8GRopiWpnBSD8kQv16s6hrSNjStSl5vtOBPHHhk
lQ8T7t8mOtT9mTb8iQYzNxNJCjedtAPslkkTa1/ywkbKHzrJF2NUwADVPtLZXYMj06FzeWmI3yev
8FItozOvzNbd10ZDLAB76XnIzy9V2z8aLYcVHkI7DT88lS5nxgGVLOOABR47WqLj0H/ky9hMNvJf
D6j5xluqCsS66G89BW+OUrzgRg6GqOY+T4nMTxaYKuvtiDh4Q4nSli5w/N/1hRCMBWGDTKxB/74s
Ml+liG3RUOz1E0rBdOY1Y+zvjmWgvzlo1pmvF4p8z9PZS/qEHkIrzoyomHdToG3924iLsL/evHBw
pTd9jLBclaGFkUu9v3JpLZ9R1zxL2VPaTsizodM6/A1qxiogGCWJuy2BA3tDPH1+boHz/RHT8L6D
1Q85v3GqOGD9hwybXmTafIdS2Fd6gPFy4hkl9cZRCk6HMZ4Uggw2QIDbjNNtLkISzcK1NKc/QAZY
FR0vK/czBfYyWh8K+leUYJ4+RdfPz9C2EaL0VdLOKERONx0v/kwGFDDUpC0hGGgBZdY36Mse3Q62
FsnLfzECiOy58Znr54vyV8mIupAjxtSgohV7Tg4xRZpQ2K63AOhIdz7o7I+zbg4T5jU2JjvPU9Fm
/gPJRhYEsa8yiBNTJR3BD+Rn3VbsDRfzJ5E2O3l2QorX/d2IPV9Cy8LarSjwJhJmEVDTjgizm3E0
ho4jmbBPhhberGQZFGBHwOTzF21yE1ljtLUaQwDLxUJNqbdINcURiWXyGxqokRTVvl6g0Htvn+j7
lYwFP6qgQxK29e+jwLRfpInXiOnsH5bjdFb5QMppiecmP0exc0aUta2ORsticKCDHn5KlxyUWUDK
xM/t4+DRdaTy/jHclh0tEaKo4jwUvJvosVCYNq49uF5UIeTs29HnrtyExSCkwuatIyH4chkUwzhK
1zHwVmfwi1c42KMJVnY4DoZXTynonZz/MdbiQExud7/h7agUElaw9GJPxk/G5WKX+tFEHszTkasL
s0jipfhmvBwNxBXlVvFYTBVois2SbOdZjxvC/i3dJ6R5m2Pl+boNGMT9Ihc2wmGmE4b5GlAvL9Uc
zhLlrBFnSx3Rq8xbO7qkfbGasBvuqENMV1aJnqzLDbVtsVsBh+20wbnjmRuoQKb5GnzJEUDzdXC3
ZeiHn0hco+Fc5sEwyiyPcXpjTdl6A1n/UruPeeGP5m/MoNfXilnq+HR0pRaiaugEZmfLU5HbRwgv
VYUyAu/pkZzs1aXw3a1Bl5mJ5ZGheGsq7K/vi1kQqVaEqh38tO4oJRkAuzO7ZicMyJlgHwjFaMWA
ZtCI1w7b1L3o0jaBa8BND4gQdRfKsi2Mgl7/FHLQjpHQhGvKky8BbOqMOkHx16BKFJEtEImXVhm7
fuPCN2EuzggZxEgArNenjLjhRc5jR6UlkMM6F+Bj65LIyouHRvuMd1j3LwaDfXi2ljL2iFRw8ZPs
83/iF1GNHj0G9lSEo7JdyU/UU2mn8tjveInxXYjqdgcg+pnxsMJuiDCGQf0J5D0+BRhSJAOVEhZO
imbFvrR1WhsQtVgysjj5I2ZltGGwbb1hHiVJDDvpNtldMgpgenXHqGOXhHy6wFvLKSSEdsnjY733
7uARQ841kDoF7Mn1hO3DRmPIkXgpi9jYBqKQRKEoE+7Ep5FcJyDeaC7lPwVsoSyLuxAhz6v3PGbH
7SiCNvAmchCMtctZ1+SfU6KZA8I9m1WfyxJF5d9FKLbNs7RXFuzo3dRxz8lKzVxP6fR3/wpjkeLc
OX7OCALUGd18CWv9GUQLrWSfTA+xJRjfUyJReeDQg56KwMhBAGNTVIs3W2nxaEjpTeM8OFXMX+HQ
p0ImENlcMsRBFj4dEEt5OaoZjcuYs+EO0ToXOZmR4GetbMjAo+4uLkpJlen4ssC6+EPEUZAgtXmE
1+Jz8ceJW4KslX2OFQtjPIZPsAPsS+RZsVduRCK+eMo94SpVemHY8/5Q5/1YJyeYJPHBpLlD0Thg
Pi1Y4Z7MQXZh8C+uWlWs7soac/YdE21Nd0FYhcRIMFjlHYW/GhEU5L7Cgtp9GbUnl8q1vQtuglIT
hEV+FYs65KiyQkrsTvURXwcoHFbfWl1OZOCmXDPffcRMDTbs+TSfmt34NlJsvx3BVOBHU97fHs1C
T21wbpa2o0U+e1pwvWFLJhrj+tjviNOuGSRJI8m4259xEu6cz34BsiV51g4um4QohstqOrfxVNIs
Ym9oy7Tf6uyl6w7sQllOIaJOa98LbQ1AgLRF0VzT9MV7uyJK3B1C7YYk/53BtvuRy3SQZ2Cs/7k0
gUqvirNtxSIXQIKrBiZEfoF/DxmpqIzsRssXqQf+5yIkOSFKWCAWafhrv/EcinDPydG3UTdeMfTs
MaTe2rp0kgVBLRx/Fm89Xn/q2u/bj7CPoIec7CUSCtQtSOGH3ZDnUUzk6BE1cx52RnKlZPxQbNp+
p7hnOiB+vTw898IYKOxC2VCEaEkRPavElVD9F7LTwP1gDdAZIxmOQaXxrxn+2yzhuQdLkAyy9BV9
uzXCqffuS1UCCJENyvBaJE7kMojRnghtzrJYlI6/+2WJSlLCbuIopjux74Gqqil4yfnmygknuwHP
gBfaY+OgyKBBaax0PbwTtppUSETAccJNA54WlCa2V3l9p1pDBjHDffGlAmvw4lW/9/+fLKYCEnuh
EMap3GO1+OKgvXSzdBsXugCOj38NKVG8wWe03Z1ojrNgFYGgKb2JKjkTFM8k2mJ7IvKRgN6zI03V
9m3/2telOYFbo06gU5FIIO/X/TuY5d09iE7KvJTK7vSaTQR5/UkwbeKrWYsxRpXKerf/mjTOcsE9
X9p5RJSSWx/bw+rwG5lkJIBBQoWQ3vVH7B2ImvQLUIImcKhj5ldKjgVrNyLA1RmigIGaud65a1Rk
Nmj2Dnh7YAJ+fVcvfwwCO4PqGNW757ARxNsaBw5KNL65qeKMaWZGSgRXq3LnursEF0ahzE9PCX3e
o72ZJk3oj7z6wdykdjOQIprQbZmeCvSBHm8ziCa0KS/dDafXMwBWZDP8cM5dSBnZ8WqqJNG/l51R
J32+BXOljiHVzpjMydOPPum2G8HYfVtgsUXFnBUNm42RzNe/vcVXJK2E4BV5Uw7elGYdRTW3gc+R
Vpvy4KBVb2+SRQcbgcbnPY1aOSkyZhUKMesLkTSoaRU47+1/CjpBMCZofujR36svBB8iKGybi8wm
0Z+PlQGnsmyixR81O3xUco7qcv2OQf/xSkT4f5nCfk1cmM7Gw/RDh2sMR6qCHYv1o1EN8G3/75ka
/SBeUhavE3QEvw9kZ8nLBEOTIgSMI4QOOvTrvcd8uc6Yp3H6+3hpTnIku/Mq7B6gIUNYnzpQ/WfN
1SEd6hhzmK5bVNZ8huci2Rl5QlfOaQveVChUnrtProDTOXg6v+6D8RrolsesUu8SFu6WqVtNmAUw
Uxxw8/HTMp2rkWZvnC2Rzal/KByLBRPGKttAHus4MongUu6cKfHrg/2W4xpeGcxyI3HGKr5aD1a6
lseGloTs7ZHuJp8ckcWt28wYrfda/71vxtnaMXPxYJP1ikRFOvY8iyqdf01mgfHD4MP+InmmHiDl
HwbsmCSR/ULDsM6L6QtyUsNPP+4gXMxN9Egjd4maxwS1h0A2O4sbt3AfdlE6TKP1yukiXvmH76ru
EuCtud5NeSg1pbVAGyRZX92XETxVmdrGrISBGTAsH7BIcJccBGHRnsUw054a2K8uCcqiP4b5Aud/
iVPxEsHrtsEEtez1fYXWNeJM2ZCwX78fSdvczRcYLtdTCJbfSUHy0J0PXLJzE/UFzQfTuTQujVae
BN15/ORVI8o1BvJexe6rOt3E695fMdwGlfeV8aSQE0JGtvb48HwZy0E38nBak+LrQZjgMoZCBbov
TkZrl6gD4IsBlJVycC6xWMXwymq7rlLx371/Yb3XNZ/YQ05veC1r7uW0T2C66cf0q3OVc1+FjfLh
mSRkbouFcOXgOy6XmDLvTtmevOWVk3HGG7+Dw53Wc9O92IlXYs0qmQRKK0tPmbiKeun1ZcWxaDcF
TG2a5GLL3Be08iKfQozkBg8mTtM8FlaCHy9YRiX6EFdNRsw4LNaqm5iytnYYEYLxvOSqxEyURP4b
HilaY6ua0/Wtzx0Z39fFW3pt73IVgn9+0hAnGSuQE4vcoMBjGq4jd3skya9G3F60SMJ3wpXIYYN2
TvJOelf6rralvmhy01fu3Fbm8/FtlzEqCUwOQDo2NpU1H1qJBrq0hT9blpaWHBlGLr09xqZl0LlM
5/7+Bz4zhG7Vr49If4N6kM63LKpzbiDwKoIMf1IjI02I4F9DuZoaYy8RiRYnBLGxH9pyxTh3nCoY
zmEcPKgiHyQP2K9m5v9ryG935PtHFNA6qy3hxOXFkbvrFPlD7JHXZ2gTr5O3CyKaUH54z+0VzH7r
v6dzfdLWCPNXzcFDVuquRMGPruHbatMG7SV9l8X6rgtrbMfr8hzPtymTk4i88UzS3kBmiQSci65p
8A/rKvn4s1MhuVd51CrO4rg1MJkOGNFAxLc23lyXYSErszQNo/8Rm19kIgtnZPCFx14PMg4E08sC
S+7bOgomLBnQHnt+xG5JSDpy10P8k3h7syJA7tkhsf2bGCnzijBZrIH8qsan9bP4y9W5tLbAGRx9
wCnNsw5BRerSLjFCklnpj+N3DYKEHeVrELy9h1T8xskiiSUoKX+x2omoD/J/KinQj/PWzOrBvSmf
NrUMXOEsNVgileOlH0yN+j2/Hq2kNgTc2Q2D7WpnsdhwRAIPIks/vfwx4HGsmiBiszEXwf2n5qnQ
5SH+6SVg5k6l3q9LpGC4tfYYHwV/TcDmMqhWc4nY3r8yXRx1nVSWC5Vq2CwDJVZHRLUICV76BmgB
uTD7EfOY4oF6CVYd52Ywv0RNFsVqSW9PZja7rVGCX9vC8mVqMr+tydxYc+MXKd70ZBb+WCTzrZ5w
cemf27gCEdK0t7HKolsOCFysSAANLkrnXq/Xx0WFj4SKDwBgee1WF0m7Pzmygs3OjDv8uy51LxJh
jCEajUPT3LHj9En2O+dZ015ocy3jBAjHIhrAcilXWTqa4irLCmjfswi5NFg9fStItjRHT1NkRTLO
6YzWhdr45d7byAT0QEgM/RpE0SoRJYuro6u1ARpv45o+79obFdSBb+YSZPag+N4FpJFo6SfVT27m
a2fMbBhGAc7ko5J4X3dCXBfHtSTOJOLqiTixXHo65m0tCc1+Cd1NqUyzkalcOhvK2mhh6xKBn4t8
5wWfsdmCnKQUqbXQ5V9WjfJ52paQ7zBtj+MxEx7hHkhPDDG9x1Y4J/0bMKi3g0aAqnxXcl6WYvxo
ha+K5W5oaJ6FgnFutKuLFH111PuPvVsiTYE6TaVYtYOHmybx/U2Z/DXVleQ6zcPEBOBlF60YHWvC
G3J9Qv8CfEF5bTBzcZdrzASO+nYtNcjlWq3JoiqjMIrajZANM2ca88nhjwthz9Ti5gPzV2/nXtA/
LTAfn18yQCHaK+0HQ8ocgHf2AWXFU1qGJ116KRR+kgrJ81cc/zsi76R7vyNh3EeQaMy61odmjLZw
tBswSMPzMO6B69Ex2bi932c3qhftJVT4FpvJj2ZhICZHQZw1/YFZCIR+EY4ccrgpwz+FRaQdF2KY
/ldKwvwROk3ehfbb4OfszTMP7YX9ajJGBE/m8Gr2LkTGmskArLSUV5HuPG9TWBs2w38HMcH3+DUm
SwbPOY3rN11Yt1ncjTdocnzxETn4+krIiLYRBAhA5IF5TKPxA1JPUBSgz88DrE6weA96DmWKbSFk
A4X842afyIwV9IP4Q6yd+Q+sOB/rPLzndMb7do6gfs+m8vqeyWWIwoVDUGb92kkYbYgob6OaQVAS
OheCBi98R+oqhbCqoNMdKP1Gx1NcCgkjA3JWH2S33TZIvgd2fPny2t34aBPNHButLzqloZkudOjt
dY/KjNf0jft51f3Wep9f8YQV0uj0a91yPYXWyy1nLNDy5o+4/z7e3oLfxlJoC6SYNKYTe4ISWy/4
2x4tXcPfTwBuRThyNfgwNVxucan/sd24sT6qKhTjhqWflzaiqDqB1DTXTCgH0ssXlSZ8xmBmX2eN
d3BN2OlApd2Z7Bns6rvwZdj6ZS8v7bNXWadLtyaprtXQOhyKb5ZILnqXNE9LhYsPDeCuMdvvcam7
v8Ybo8GtPgBFDmic+vF9Ceew91iB3RoOMmxbKjrvLL/H7n4DgsnynQgztwfkUcsN3ktLR57sH5QK
q26SKe6lLcnwluqqSLt94edAzSNn3Ll7z/lgs2QSfonVJhrLrx4EjAv9n9F37qirDsN7UZtoY5WJ
+ZqRKUYotorgRMgeFohrZltygZ43cBkxmoMnc3KiySkOPtuTxcwsiq9hn+MtNbi1Kne1cHoAFSww
/in5t+3V1OHciR57a+YCSrSlI0assXDh6rxljooE1OvEIVQZXhyOp6BvQNL0nVpuJcE8O45C+MLj
OC2N4fQmp/TDvhA2xjOMttQlXoUix5y60p/EdfqT9q2DNL+cdBLj86wSaw7to39uPIQx27trYtj5
ExwYuFYDzht7xWIJt56ZcuPvXYEd9qoCmE2DnnWQnQf1PQwgaCLnPLaW+VM/Ky5dKQqd9TK5TEC5
rDRUGAUdOeOMb/871QVTKd9jK8F/nYFvZJY5jtuoluXRSkVrnvWrHHvKQZtHzPYVweLRc4UnJepE
N9c2+n1PnR0vHmkxd7yBIitHJFCmsJdG+0qRxjObvcaIo42hyqZ+23xhx/0r/exCQlJOHQOI2/c0
D4FrHLyjdrxENnD4IJAjc9JxsjHSBB39VCW5QIam9Jm4HkFgfXobBEwLccAujPRT6O+z+nLSqyW+
chOcN3OffmUHtTjUJTd2KqChC/c16Ts5aXD4En3BvOuXo1/jZ4DV1gKeowbdIQcqywUp9VntjXNw
bG6vfcWOEdk3to3YQS516PE/81rceUV0hoLvUTd8k/z9yQwrcHaY70q4dZ9HpD19fNI6j21wJY3p
NP6iG7sMe/VYk7Sux0/ooRWGScbpLtGytfNrurSzzh2HbgEtO+bYL/BreGGvbopquMG+6LQrfCf/
rcrtOYuSq1rYt87uKbxZje/6JI5L5Qnawuwb9dBgY+4oP1VlBIaX/8sB1SDOWxnTYvGGNi7J46QQ
r9WEg6MHLM8PHe4zHm2wJQLbvap/fLl7Rh3kqwt6pfCy7i9MPq6Le73Xld5GCmxF/qOLHycGzEYm
UJnmydsuxNLpGC7IzW+7ulSMetalnayP5vknQl3ABOAEWQGNkgDwBseGY9gaiIwXav+tiXmKDv5w
Wg8rt+BkbglyeZ2E47CuVAbYOFV0Pn6C9L2Vye9MzH4OSU6lLAC+s+CjOLUkOCZPPuunpdDU1wYL
JWCF70JLAS375uNhtsdhWPoeEFLcwS9cAYsZDSqO5miAik6jKFXbjPwu/QfNwix31hZonNTbX0m6
qy0n12mebatmj3G1oow7WaFkvg6Wyhy35ju3rrSOw1HAbLXyO8NSioF+KinCKNKgGpvxL9L1dfi6
3fSj1z5tfndHPp7h1Qy3RlL2BwQPXN2OkIp5C3eByxdSc8vdXFszd9M0+tPQ61D76aM+uO+PnPHo
m0kvVBD6shw85yofdZKroANspf3wCSghMjml9Tj3mUOyyryp7cbZY7BVjYH0d7p0RA3YRPEq2xNU
7Eu1TBusdJ8EJkUdDlcOtTFwMbA0p6aQpLXMA/eo0NQ5h5CKK8CecuTxCU1dZpOYNwEbfJ2RQOQM
mgAN0y2carUtIQxwcGY0Wi9of35vTfnx8tjr5/HPWb0337zsh+JqRov/cbL1Jv+S4+ShUI4QGQNZ
PugB7dwgNu+ZauBDhcy4BawZwW2r7ld91LBf2/+fYr7UdT+37+4dJiC2bm2j3mjH4THcNoR2DmRS
dog/FuybSliLDPlPv52axl7wP9fjRML01HsQus06vXdCXMOpPQWYC4Cjbf126sJ4fTVrYBgcWWl4
lmBp4EXZHg+rd7VgdGize8VxIRRJ5EClUgYf5QDxVdHPvLoqSN6gOz67hVrGZJlFTGOsPtojrZRa
JiLFMFMb5n2tsKu6bQjTXiKxGd6LxgCt2O8dpHsjfQqqTJtSj/Hl2alHAD3o4Zq82LOMpcYagUCC
CPTWfXWo0sSVK5PnMtDBiB5u7j2j1Qy/BETKxyPgQctj0YLCr37dofP/EEk0YgPLvGjmSwIZCwWr
SqQOEZ2zWa/+XPB7HkWi1eZmSf+IeBtq/TDFJY1aII5IPadeJzDhPetiFrJive12UiXjBwMqzwbL
e4by9MUiDfyc6IrbKq4ENVInFTtzPGfROFVr4aBbJBrFwlF2BN/ncBTP+09tvELW9JeTJ8c/QZi9
9OP5uA8/QCZxT5I6shMAldNMXe1SOS+MK5+TgqZ7Bw1ls1eWiM6Jza9h2WGb9H11IpYc3XoFKRmE
xV20yr8oRjI9QdJqbPspVNbkZ40LwaI5kbCpdeVqNVUjjM4WDeM83sllpGjQ6MufXX8KuUER3RZV
51Ijf2cfZofPJvI/BMyYCMeuH/XM9KJNmvmYdkZmuVJxfVYttwOU0U3vTTupXGC4UBVggvtzyYYG
jgCf+BSZ6xWwVYuL0fbG2fOQnLQA5hI11EdpGEUFZSf2j7HytrdOiW1xUNqNq/dj1Yu7Og5qcbme
CD1r3L3te2TWyqH6ZIWJQj7ycMtvuXk6SLAJKmzR2Gce7COqrvePTKdg5cPmWdrOtUOUedX3AWYo
UYFyNodosQh5AGhCv5vszwKOeUf4hg+wZDnKH2XmRWQhHJOUcAq9qGxGAc2hHzovSDnr0xWOq5s2
ubHhPPfyNPZiqyF+iZuD9wStgdrkuGJM2AyNxCL8kujuUNR84FNwLa9DOno/DXvRZ57n0BVBNJyO
65NZUxcsS4+5G6d1IB48iH7eTHuTQeXmuaBSJU3/27dZOsjroaheCrp6SJ1DAD9jIIitplFzslUR
aMgB8mRMaPvHPtBlFBmLcb3iEEpYkhHV5WTnmZsRRNidT7CLz0PwLkILJVg48016DathZYQBNcLo
9BAx1FhTrqIRGfr+gF60CUifdNrc47gz+gvBgFr8KI1WMoPNHvj80vkdseQ45l5DG8zEVlPw0oxj
b07mE5hd8jdTSXeMh8gyHxKsDdbQJkeNEHWj2ZBc7vuQkmDPBX1gN3WJr1nTnM97hFtXx9F9WxmL
AxgPrBAKWlra9Kl4lwW4wzYrntNBp2fr4xUqbnwGtDtKM6WSBEnzN9QpTrUaM93J7Nq31P0/ftXw
HqSnyw8UcoEdvPrhhxz3mf3oR9rupJSfBi5pPxcHCazBRZNxZ2AWKWb6/X/P0Palm36SrZ9oRVBc
pMSXfpxKPOgTAMAe4Z5/Jd8JKGFyKUMYkEEGgEnkfw1BNU2rPoFRIqLAX2B87X/vtTlwuORbwjuC
HLP5ZK3J1dfFarM/XaePOH3GBHBT7mKa0MzlYgG8ojTpT6dQwnY71dj/9rk/vWlJdo7hcgNIA63b
RZUmrTrzzRpRstJnOmysNK8gkZqQns+BgRc14n/2zMpAlnsLxogFLlHyQEKZUhVC5yGLc/294E4C
Oa5cg5UuesNpX+heKmFls+KWXREmkMZBdxExcjtZW3LZrUzaZdvyiJM95dtU7ein+tOxnUU056Fj
26LeL+hn65+8KZBL1BY/ZByvi5aZuq4srY4u1u+fW0Yj/O9xKY+2vYZ0FkXUZThe5AgaSY752yXL
kJithZsmwRYydopogZoc7/G1XMtwn6AtScr6FT8KGT7/NyUq3AVNM1pg3RSx5dFSGwsbjdXRhPN8
p3YlYBWiQX2kWiB2PRUCujewhOmpZhrfIAk1YYv2RPIycXF0aJaZJiQuUPrVgTHZ/ctybl370X7L
be+36HBK6LtkFsXF+R3G9ihjjDbPV//WuXsxn7R5IsO/ljMtVry9CTdOqZYoDnNeAAzVE+ElJ9wx
rO0AlcMnw7H0KFtU5MmShtqO72LrFQHAyEGAs4VhnHiQJ/1bw2S/D+7dBdesbrdyzKoy42uDPdpi
XzrNWW16EhnyGSQF7ZftUkfrDo8sb5Hn9GYX6bhbhILppqAzBlaxuImpqLWITlm/yrQvB/Ibs2H8
/h8uQPdBZUiIgquT4kTzJtT6DWpbXQWPfQv/CnT1dR2LrmVAqMZaPFHxATUDg9J96YY9B0BL6Nqo
3pw22cmKamyNuWpXu+PGmaaBoKbM58d0re7XWFFS+AnT0P6oo6q8NZqSJuXB1MoR3FOQ36kbOOQz
NHzP1N3h6akekl4NeqoEHmXWziiLSRx816i4QUta4smMBB4dhZ1nvVdfMGUED8476tuXKOquN9pL
pW4+1b6WE2284eM6u/RZFEyJj8k8osKcTGJjlJZFwC66R01yEyTX5Ph/b8VQCfViy6VNkxhevjwy
B7VLermG1KilTSZKJW3/N+P1VCxImLP6B4dBfiDjfG2s0IXafJE9cpw1T4E/T+ByEC6I/UM8aWo+
UgoTU8FBHW5d/ZVg/PJ6M7H/GVNnApLYhTE4eEZ9cdov0IQUNDJmkY7KeLMNwpgDi56uzKXYbuA5
7ywUQFFRAuGMepOMM7fgVMJpjW+MKPwep49BdyEGg2IYja9GzMeQVecLg63uLEr16PRuyMK1LxDT
GQy5jYlcMie2boMMjAsLUGqpeZac54Ry9DIGf87QIJp4iQGc0BkzMsZDsAEZLtbh7DDY+9XvqhWS
z2W2c3d9oB95pLslrSt0lez+AI8ypp/X4SiuhmkyBDjV3pRpfVKUIqRHO4gKd3Ax0CIHpOy4X/lU
hKqaAiKkNSVXhIJEaiGxHNl6enwxsGjZkmvhvhnBXsVh0/KG+eOF2tGyFPeI+eyua/PcB4W9mqtO
yVMrzXOL2zmi5adtO7Y/UH1rcVSVPd0XGnxjWT2WsK+HQVU556fHuLspqscEcf+it9Jzy3jONe/Q
Qb88jviEAV/6uwfPZb035DX1kHRDqfh4yXkvin+26zwULcatrFS9gokFifzBbqs2UNOSd72OktYv
RDrXOqJy9CwgLFqEBlUjgAM9erwuMVcflMwwVL05SzfMbZZiJT6Upq3BUWdpX0CFYvwvmqQvWpZk
hq9eEbguLnemmG6Cr0IjI368sI+OInmhYC0uhxBN/WE0w0k7z1GqlKJG31eJ3XFYIXA/DUHF5hyd
7HazMzmKa17e5k0TQeppkXrCovKztHOUYH/znDNYBOceqG+teo3hcsh1DsfeQJEsv/2YQl63N63B
JVbLooq+wqHUsz5UuJnnNE77DRhJ0D+DAnvLo/pW+/kFI0/wNjSrNOh1YkFb9LvC0ZLlTlhfhRw2
QqBdy55mXGvINW4jeEDHNHREDf4pJGqtxzf1XYOAoJmLaw/dmDT3memF3vh9YR8JcjlyiqB2cvFw
DcZskqrPRDO15ZWJYuILFNDZkqyJZ5k1ZLb7QzXlj+p4vdhMivw9wFxcwIPoy1QMFDut/u3JbQUZ
aqm8gVAESWmrHmpWhZ2g6/yACXwtmezUoHlFWWvbyDD7SwB6RXWPcAIx5ZMO8IdHZshYW1jNnRgz
VrCoa3HRbbirwoaP2Z4hhU+YBud0QkPpLUg8T08GxWg0bc0KlcFrgjA7EdgOnmnjFxuLBO2/wLBU
9m0tGlrOsH795pwwoJ9nKybrBOn5QNGub8AxT5rDmm9EBxbZ++vOC9WTYz5it5Kqh6/ivH+IHmcr
0aTuA5+aSEIPV/Uv3ZTqioXn0WuFgV2NSmOlwPuSOcpGWoRVE3CSKj7A9/L05iYgRuy39sAh+cDy
pLEiNVY/UjgrJsywWsWoLCpna0nhPeKWv7EWMzoUChL88EQeSxhTeki2MG+hOUUYvJ4/piEGaSDo
buPzy9DZFLjHJws9BOnbkEdFbz/Upz53P0DTF+ugezxjg9UHxmW5smAxdGlUeduPazPR78anjbsG
+VeKG5V1VZe588PnY/wzI1diE1Wc2ECpGp9ZG9WHcHRtdHgTS5WreuV5p/w1dqWhBfcHEaDJHPL0
Gg8hNuR3zTiv5bid5VqOtJ+GhAjg9BwiUuoFFCEOTZdkuMzZkcYzdlJ2AY4MZX/ltB3LeGfBRSdQ
FJm1dGM1QNG/jIjw2RKxFvAVFWGnw4MtIne9QlBDUvSL3F57AWX+LJZHkx23PgmXJ3ToVWfJEEZu
TckwfWkyIdPEebAYoWhJzs0R/7lycf/ALUfkdmiI6ob8ojxv8rLiwVb/HalERgxOS4BKsi/z2tOz
jwtJDQGx8yGosAUX2tETGhWnrSanw59Ku2wunyttFHby3Kx1biDXaGLyi4uO1KredlaIiZU0mClb
tgNOSeDqw+6iPCmc6Qm2cOv1+6svnXkNoUJ5o9KMGNgsoo1q6KROqZ0Ya2FH4KgEkGvCTI2G6GPZ
cTkReP1N2UYGhmGPxVpDDKCvPKqA4CLCgFxgAXZ8e7Wx6EGFzq/yzmZmLLn/zLHi1Pds91pd/pJ4
AtTNHMQ3zsKIXr350JlKh2it4OoB1Rgnm/aWLzECjbpcAj9/v2UqNHB79muQhEAaH+W0gu30O4IO
L9rrBYMWfTBPOMitqnD0P/Xxx+/M9B84zUp9DZKI/s4UDxkZnCmGz+yumcd6AnefLHWBREdiNnlj
uZH1ZoP71J+f0h6YEQB0lyQmPo5MLUkhtTZdhkbDlrAqiz1sBDVdPgqBSrTDsz2uQCw4Mf7EPpFc
YkE4xd84IYglerzaWukZhEgEa7WjNtmjh4q8lIJ2MFrOd81g41imFGrHc77tLKsgGgzmUbNwJeGU
5Yn3rM+mG3tBJhYUVMbEH4FPf4qbx0omYXrG5rdkbUzZ4P5+JPyuFPoSr5IKVP2jqcISh5/8JsEo
Y1mFnQsLnEn2hgX+ZO1LcLPNdLsvuJV11hRRLhvRrkGVqtCsuYi1B3mtNahqx/Y753uvRvn99/dJ
2MQ6NJiqOyvvB5FsdKXpWuJADkIV5BFFh5+1SYeOTTlsaHFZg+Z2hpZg4aaol1Uoi9ZAbdzkN3r/
tphbCDsySq6/uY5tZ+S5cXdsWbeEtORarm44xCQXydnyTgvd1ofAyB63Mh4h7RwH57VuMQeptakY
1Sdpbp1LF0KW6gkk1EmK4Krw/FXZpzNa6d8VuQaR/5Py/+HkwL4gJCMVGabayZ39K4fpqdcKeiFL
24nEwGrEWiENpe8KvuGgmQeiV6rNlSGwfIbGtnXg2ccllSOuhQcFtu9Y+r+RckeJVLOGzIfmIP2z
IgwRXoX0wRunrKNu9aBpGS4LSXDYROMktij3faZPeJWgExgJiSSL7esYCwGENye+Sz3ei/9xUUsu
px0b5Su61SBuZwtjuQETTYATsGmceU3gER2wF08yB+k0XGUxlavgMGtBDNIHlJ8E6Om0XtXJE/SV
+ZVZfmSujjRknJKXzYUONESWVprrsoytr0XXIkVWMaIGJidyXdno9PskXAXG96t7BBdyJ0yI1ciK
JHxAr19gBIQI8qkPDM8VOd/L8+T03gbXE0MT6ypmD7sbg0uvxQdnoP67N3ciA31z5C1fZVaXPwkp
J7XrrOEoGFFy+YLW6q8PlKFHzpHbonIiDOVj+VTZuTFQom5+Q3LDAPDwQp8c+GfVMj2+cdS2iz9K
x07Css/IvB/yVqntmsnK+4sDcYrJ92pBi1oEJdt+9OvwqA/JuXIjbSe9Wr9xEAs83vpSUrOPTK65
81LZtr3+bBBDOfAUQKlUE49nv8pd6lqLa3T7SLLPjOzqysQDqn+ilHBK0nik3wwGij8QCbeJoXNl
Ek3YXlT3mFlF6LfJAkbTg9hj8d3ZVplya+5TVlbEBc7DnDsccmWqloQOi1T+FXiL9c2Hnw0sXRvS
/jUt9XIvl9h2fppEsZfsAw2cA9Xfl9LrRRxq8b3rhBqE6YIPDiBKTBJebwhkzJIhaQAm0YM0zykF
T/AfF6isS2rcyEQV30YDqoEauyacDeobsujnOgoFSXwQ56l86/K2UNzMoUx1IhvDPhf2KWd/M0Ow
rtBTWtU3SoE4kV2TiVy0CAwW64sNSIXhaf0SRj6AIKpjwClTlCg4Q0klg9DjxHXGZ4YTEkM67UHK
D6jyv9ihg1Zog+k8oksZ/ExpPbcJqPPRC4q74JPug3LhhcjmY7nHU0wMXP8GDpTmhEo16DEuM5un
3vRCaK6IUxorVSQCAFwOJ3wj5Kg3bd88DkPpIw65bqjO2ItHlq60S6G1RyrCe/L1MNeHnDO7w9Wi
o2yhBCEf6/bGJtAD3rKQUFr2cxvVa3kjINnro8NCbj+fjzhxU7n6XSWLUNFOPf1wxBkUJM39Y+5U
edEBuoCp/P6h9fbqh42epTVJJ54wu+1mf6sBFME93B3T9PK+sC1ggS3y/xdYj3ZIuC6zq+/zwwrH
AfbGozxr56to+HV2BcUZ8qzkO/p01oRUw/hJxJqgiDG44pJ05eSq57EOT7mIXdRmhAT69Tzn0RX8
DSW6F8Zm82QUsMEwNweArj/zYqH43TO9Z6DvRb5VVSV0tCdJ2yE6CBlHQJGZlG3Rpqusys3UyYdD
72RJoHgDfrFoHB2NAx0qvuPP7tBw7/KS5vIE3oCE36t4aRwcb37sW4J28F/Jv+RR6/DdbyLsLONt
iLSZUUt9NXOPF5PR/WC6IUvUXNsLl/m1re+J5Myw3iUVAvMs4HsHLVXKlzyTBhkMCRfM9wmA0GiA
lmp0YwDCpzZwXLD/YDSr0A1CYgjQql3ANlYglfuRwYX2Us+DSLgDIUc6s/rjIhNGGCJ276V128Ya
Vwh72+c1Yux+MMgZ2C/JNr4Iyo3P7bdzZyOCrplJcvWTjW/O/jPNZa3b3PnER24EYLfGkBIvppuT
u+X6Txa4CGSHcH2P+JETP6q5PBNLUYL1fAfUVPJyXjadApxU0l0DZ6C8vTKBi+XOBQGTefiNhMOG
es4v0Deog+oLLagkq3+ipPwak05mBeuj/88HZiPbMLyP471/eWyWGV28E5Cs14q+cWsJGQ96usxU
05dE8h1/tTEiSoMzKepwskjxU4lbiJ6TQr3H/zCAFTOr+iLu+IxO3TJk8Jc3Ao7jvjfduZmU/u1L
NB2z9w7n7d8b0O9hpczgSyQhguOtT1msFpYilZu/aX+Qt6ns0wwyon7c1t+60uNeV7ucgTj9F3cP
vWUFHejkxNqDLaDcZBzey9g4wabGHvdD0qBHMfdK5bzYQOy04yeBk40nIqPiN2t1yO6rKUfyU1JO
4JVpfgOzMPk381yiwxQn6JjPRJ9pUATDN3VkVG3MxyApjDERE2Vme0TY6rO9eSSJfj3ETDFPNiXz
s6iYDOQQ6V4AMSxOEQ1DJvmccfMgZ7i/s3w0MfZMej6siSQVFxZPvYwmYN/3vSRwcg/W3sDRdgqn
mepKxz3MVSoMuaM6/S5TLt9q+CvxbSxxOqaKssxqj9zZSFqhZqODBVymcQ1jiY0v0xLu2bZG68i8
Wkb1gfUTPslRhg0gO02taA2V7EfXVPPaow2ULzCCZjUx7OX8rB65k8UZHy+RpXNawwxiewFePK8y
mxPsrAE39+iWa0FJMV4ZVSQ4F6FvNIdurCbAi9NQEDKeWhXMFCfe3IFP6++Hsnc2k21/LaBhRjNI
VzXhX4sdeIg6p6bW2LiJv5E19NG/zwCZa24WSGF5yw7p03lRdJRMwdZ2zaxIxppriMhFCBLHyUjJ
LfdCAv+U+M56kldBYffCU6YVBsW7VONxxkNZRVfgHSXKlghD23c9dofvGpVDyIt6F0m2J6bwHNi6
ZVLXDqGKLyTnM942zLuCYjlxdFn5hk/bfFVmOLLg0RLsJN8YmpGq0eASz6CiWH0AsR4ds2VvpvD6
8CyrlhEC3zh0tzvVHcL9O9Y5ZHsQr62AaYkq9cE+nWnmYjAq1szzNJQkzVr7VC80vYe32L/OXfq0
MHwLvdGw90AY+CF0SuFWsgcb83pkIwg6/lcSM0Lky0nxQTqmWCxQC6vaLLfJPh+3u3QSeoqEcbMn
t7UNXGxTjxR6uJJs6PN5OYy/DFwec0s5qffBUa6SrM0gkXqRq5GnTn33rb2tsTuhzecDYzF2vKeC
gZt/00oh0+0VPLoIBqbuA2WjziZFdMyGF5qSERVgoobQc8rhY/QcOUg/4YfsK+M+hhQ7olVUFO/4
QED9xOHL8XubULtr8I44NZmZP+nDOeLxIbDcYOOb2IRJ0RxgKNGzRtxcoJJafkS0tQ4kT+tXskMr
mx1TqcLjYiiJkA1fXEeacT9WVN4azZDLFYCmxxuPdyKqlZTYOs2Yt64IKZX+Whp5WL7IWiD+jP08
yDsn8LOFxO1i7vPzdto8KLUthwB+phgKvZMRy2l/Qje8drj259J9Wq5s892YjcnF/ikInglXOR+n
p24y7vFo1q5hi5uwSQksa+fGeFP53Qx+JJUpcFQb2ENiK3coVLFZkjsQG5e8w5fgXsZuCDMKz/h8
yC0N0KvLpaWf0QgURYItgqVu5dqQPDcK2FDMtG60G+iKp8CAnOhJrLO3XjuGWPCB7Y3sNJst/EM/
OhlcJUSCQC2Sky3r4Yg4VBrWOpZWHOf9YOY7oAlhbDzA4oZy2UMXOIztHS565oNc5MgQwKfaBGse
g1wegftnODGQops4f9/lMBdfsiiHf6nehFZQE1PSltt2cYKmld8IcVg2v3/0YVW6+priYe4tT9VL
EAEdrAz+TPARKG1+oVylp54rOjKWjLPTeGwNw3fvdBYomR3hQLXNOedCorOTCPeWf47Jd33xD3CC
R2C6kwnPQCiFvlsBCH6S7TGvKmOlRGfbXE9cNbsyjezblaMYvNrLVdVIYGNqxI5hw9Yu1bgM51tD
S9B4wqNfe/aluys3DEcz8x+mctVqv23GFmO6X7yLCQ2PsbsoDc4vg6Hd8ZJTEZKBATPBAFjPIor2
TQJsTVqUApTPU7X+r/qE4H9eH6KRxm7esNtMkczbbnSzAt1ufkO0lDB9o73AHNvrH04T9VRtj4RM
e3DC8FIF0QVBEOSREK2oj3mBb7y7CytKSoORO+PAbluzKtMR6z8HiaGI4mMj3EpzfD46IXhuTjtI
0NR87rZL+zyplOckrjS1QYyRjf2bKPB3XlIuqR/Q2mnvgsm6nzEfaY2gdSrZCTKtwhp2r/7zQdR1
h7Tp5c64sA317ciHyihHeoczmHlFGml4s1wwKimfGL2RXCWekupVKTeKkPAnaRMhSq4zkb+gB2J6
NK1IOg9U29XDMDDDxBoITwmM7MS+0Ye0tXLGSRuEVHskXfi37zcW0nBitUXC1DmCusD1vcygJzHL
koKhPQjNGAIqgok9WN0KUqYsaiUxC5FaKHfreY4dROaViv+XFkj8kk1Uawl8BP9Liz9vMVWWIZ4q
6jTvd773eVQue5kdzdo65lszXOxhd/gJvuxgexiFCv+31/vt2voygQO6YoCJmBpPZysUnEn7f6Zx
afJPLsSbOseZab394ut7GzlJrw26MmJAgcpuNgUZ9i8GpanIy8I5AsBJxuvt09ISb6z72x4E83Bp
01SiefFZvkb3TidoJFJTRzRh07BLgJEKOJYgIHhcaaX2+FfbyGD/JazCmcsShSJr8iNmBMEyl6Iq
L77L1n91k6yWRg56K0wP2EG6ejYKUv3X3ExsBNG9zeoW47JWFxeHS/tPyn1v5bczsmvlwnVwo9TM
KL6rOFSNamSdozrwsAf9ou006eLQ929M4l6/pkip/a2WQWSi4YNEwykGZp1oPTeUxgi49ic+96Do
c3lC51/pASI66mw978hbsrHTH2iWBp3kbKd/MnySeIgWVYsAbGTgk4uuLbLFAp0ABiN6NytEuYny
c7aSC3teP0WS232K+s5IqpAR5kiZS2jI0ptxQn8EdRCZuUBW1uZ+jMfU39HLX6u0NoYPDedn464J
wsV2azF4DTJXbaBRLFzCOZFTZMa/tAhrfvZvOAJ2WSdYCJi4DaGwubR7T4C9QsVFVEN0VhLmQhvs
LAQaCFbeyHGHeKeROWC4F/MNB9lrfb1GhNAF3Qp+A6lXsg8Tqm0mg/GJTE0CYzTEWAVamIFrz0kP
n8Oikd06ceEXQBJa5rFE9lMGxF2xwgfa3rZbShDjfKNLpNwmIM8KY/aGCNAdHdu3M94C5CW5CFkp
sLo2RIw7j91/iM+Hn1bOyL7ipk/9DThld41wJa3AnuF5FpblACffFNT+CShJiIFoT0jiVXgF+bJd
k4g/xYLZx34VbiAXtU520WhXkun2pOE9UEYhBN9hC+kniKJtjNJKEiksrC6yjtNksUsHEVElSKSd
WTPQMEUTCEaaqxIPpp/AXv2sC1Hfm5jjQacUXJE+83D4XQ6wbCMZGzcRLirw/vSUkkpSj/QY9vr6
NLK5PQ5v9Ce+dYnQZoPRBcLzPpRl8XGXNJrM36X89R6CGmc3PEdC5M5rQB0Rzh/zNVsQ4SMDOErH
QJsRsyYaWbwih3kifxqN8rhDwpalvXzmDbQr3CKyrvhsP27HChjqD9VA6MNshls88QZE0AapRiwb
mgeGPMZtG4r0ESMspx3z9rHxHq2qFYV1eevMqQcCDoydEi6gM9zPg+lgo9FIrPX6fxcHxbQU0Tew
i3r1aH4caJgkdTL39MiwrEfOT2scla6cVXvX5RTEB6DSlCdX4jNzVqOAdgcyP7OOLB8RdepYomhH
Edn5Com2a93YDCMxoCR0MhxRzntJo+pJL/cR1hgzytREId6vm6RVWRUHRpLnivZ6lScTYamDd5L4
L70V1CvnW16qVStJnNWRO1UFegz38Uq3OPy0oMoRZgtb9bL05wq78wzzX/3YgHldB+nZRWp5cIjj
xINeLx38DWDgA+9qh7VTzNs7LECACAPDnHGJL6mrL844XId5UEnMQ8hewd1Vq0vWTb8oeKSPhXnT
ewH7ZwOmQlvprmMc31hyYqLahApBLarN6LCnVF9HyBNrvYbb1veYuRD8TG8Q8kqWVm5uRbsTEwk/
TDuL1oXpPcgZpYGudeYQ0p+tfqLN8HJ9n1ld31n5L6w2VuE3FXMHFXUrcgXNk6dTbSFrExaKBp63
xPio0sa9hCMMo/Y8SW5VKAvjDwFSCKYZ9NYe5vJ5Om6xo1pTafXjiI6+zyysnNXBKoybzfOICEQB
ttGQul27d8lZ4pQh3lnMo2zafpUenXmZwsk+ZtKYQXgdIprmWv7pyW6aeICg0Ao8AthJM7xva4WL
tO2Tkn1NQ5kVoQF0PwOq5FLr+GtVkFiEaG4NILKdl/uUqVoC8tx+JM2tAqfhRH1KDhL3rkOn9EA2
6njVF/mIANcEtH3hGkmeufKXxvsmwxZyKLVsN06oqdfMTeIwHSMS2LjZYRFDQ15ODX9SBLZFhzE3
FNuoHhDFyPTWz2mN/4xThbtNpYpHdkwG4R11FalWkahB96ILid4sciVBH4IK92kBR8RIbJ+6go1n
/0t4RXWRNgA5bLrUF5g9tTJEEDjjmvFDiMKSIRjf8CEALuumBYN3hGMWv6LKWtGvDCTpGpAqrPh0
0T3rdVZ/Adkt3tm4jbYLIgQnwK6bjdOhgzmH9m3+uOhBErj2fmVn7xqpuU5itaOV++LZJ/VBTgdq
8dK3JFQAMssHXv8hSHKIf5ufnQ3VzoAptcaTY5h5WVHnnNncxhMQc/RxQ6oNCLk7hUeFdMnmVl5R
67xcPDvXmKMXjT0NW9WCBIjwPH9WRzA9D7IiA+R+oLK9J9FbXAHSkgxZHGnYAkDOoaRl9lTYM8fJ
6lOmYNUl6k6eSbU7etjzutZorIPlKFETwSdUB5gHpr7rIziTNfso1PxTBGTvlyilHNc3QmMW3Sz/
9KYiTwhU4CfgtJB/2YJ6L38fnzTxtBdkXDX/x3iniZpckMa5GJ+Bw4VYgcBOyXt1sbOEYkJpcJNG
WNQsTcxOnwIuPEMPTrxsEisCO0q6Jff5iKDtKNIU/qolRz7fO3szxdzeC6SLU83yZUe1/jPMWtsz
yVywtRvUHx9pcoG0bzNPwWTJHdl2HKmYU8ckAsVw08jFd2Ix4Nte81nnL84w6js/22ucbLxkGK+i
SNBx70esbEJ7Ax/pe+mbvRQnGUBC23CCTzvCsIHZ3M26igTB3Adz5XMW9hIlBchMuyhEEmjMn8Qp
tL5sziJUCD/bNwxXasaEr+Fm5dqIKDcmPIXK4DrBdm9s6uVFiMGkgOdbjmQUXnJ82ZMWurmUeJ+l
PhAYBsw2lLDM0eRBKIjZ2DIOewPTiEzn9nn7T/BvoERP5n8grR5h6Lc/CBw5bg46yWA/uQgMxvMG
Amko6uYkkDFrg3j/8jB8aq87ijjFbPXltP7aJHwLfUwFkPvwDaVzobKFfE4rnxO+w7MmXsuAHaj9
2aWjwVs6YT9tudR93zg4624ItSf+7wYS9N5PAC9O2DcETQv7IYQB0ltsMP0/vigQdVwXfFarE5hd
kjLDnb3EWFe9AISYuzBGDGk7xlyB/Vffvi9jfSDLnTMnqdj6lHgzIv3Gp5fhm5PYo+npCyQu+cU0
3ot/0ZjvqMN3949vv1wClMlrug2CRAXj4dNMWKrNLsg20TZFIU5xQIXnRfSJzMJPmSWOEpYL9zbf
yUXk2eERpRJzUdE3gsBmo1D5146CsYWwwHukUK+XNsP+OCMjUuQciTtCXsslkx3DhChtYZ6X6qcM
9ld2hTWX237Y4vk19XfiuzatIpxZOhaJlOtzh10eq0w3zl7SM20l+9bROemP0j8Nn3o9CJlzNfLJ
FUjHH+zzimjY8C/rrXkiCUlDhIYENNP4P6A6MRqCllhH2uOYhPzSd3b/TPj9uSvng/SI9VezhfD5
cVYijuz0lTRymyTEeY7TGonCAWtW7GN+s0PXObxFVeNlbhpm6nCZiY8Xp99LFd9a6kKEJQ+JJoGO
Vv4yWqQDnU0Y3pnk2pu/pEQwrijAMoKrzVmDBPeoIXtZPJnYGfaCL7Za4GUjjRHYRSuH5GmMmUls
OMUgnYjLfp6ohXicB5hntITwG8oJh01YM6sYJd0VhgFLdekH9JDL0SX/kKWxcsQdWkCYJ/StypQY
AboYh4IzxktGk5r7OMKJYbxxoUz/LgbeLRss9wHg9VuYHWUUCgbo6DWok/1venaOGyECD9MHJ9h2
yO74LUTGShWPtpVz5Veppxf29/DRJqCfkWjPsPWOYNYt/CWkp2X8bnxtM4n1eGrcENLXOSymIsRd
49gatMMBaKiALz0lLoGksu+XloVf208wdVhEnswieKpM7kHYhzB39qWBEuJHKmm7Fe5I4QTO9Hgq
CjgzRR7Yd9slsXsCFq0Mjoo71QNMQN0tXfEiQxf2zuSy6cVw+y+s5Zug09obZXS1k5C9qns+ccqD
WnIvyqJTtW5N3R+fuaUwn7PwSXAmYoP6kyvFhmFXPzgFF3dYkTlx0gROVXxbGbutdwxRm6mhkqHM
PEgrMtcQx1653ZFd58cBhNDA8VuZki59lYnxVVyM4gdy3b3v3Llf7p/FkxmuwapYK0vmzuY9SFmv
MxLPdN4haJYeNyKiFwM68IiZoQ6XK9X2gpzsM0jRdz/sNAn5IAlEgwEVf8btG1wAYUbdlkIrzYa6
LkILJyFXimDYGugGkZbqPsuPA0TJAd6bHl5wIRqLJXig9wfVUUcHG7OPiQt+Gw5DLc+Qu4xZg3at
7uGH0A3+Eer6vCbvjhDF36YqNbKLLleBG2KLL0aUl27ItnnR+kD5e7sWwlHBByc1SwlqVf7F8ywl
qwEEORBvBJmmlUbQ0FQfqlMiA2XhzpZqqxdLt8BLVcqpbT2+3dIYEmvR5vooDMKv5cV/GAOichRz
Gnz+DJMG+8KItO+JivmF+ic8D4NXbNEHCvS+A00bYxCEgxfq1zg6NdyjKUurIZZZ2o6zfAk38JjI
KkQrgYxH9d6B060SQTxoJ7FA3T1fbdo4l1PJNr9X7sS12Ai+YWElN7jYZ2rp+CEVqfN+QD2eS2Va
5pagVDHxkJ4fUJipvxOmhNVedvUDtS1Ln6vUZ9or6FbyMsx9oUzIm08dvT/LIXnFxTmiIQqH6DD+
tJxGicbxn0NmxdcQ0azQYZ7BN6A+ZGH1baIa25DVWJa6qS34zX4LqSG5qKbTn57wH+3oGcPVk9lW
Pnxd9THuJ7QmKStdtXlV7ppwz8i8di+DRDhjrRi2TSdUovinOYP95Tzt5QWFhvIFSLEtE1IoIoMp
DF2iKOG3BrgPhj//HwQe/LwvPlj5r1ROQMftpVL/K8rPoeXr0Fbpm79RMLKYaKmiPYSLnZurDjUM
zOWCPBzUhxpbUCs4vqzeKXhcbGSDWpuuW/tqyJ/ft8WuwFKDTUcD0XqwbdEFhvK0kufNykWm0+08
TVYrCejWdh7DPkj+vvqQx8k5Qxkp5FRCsVTjJLcs8xaY6aAc1lBdVa+QWgR7q0z6Ya1H5QCRM7Vm
DPf5D6BLbpAwMnphcq9x/ifZn/3LKX9R4QJM7MZEpIidI0BDntoCdK//ug7153Dw3fyFFyspmRtr
LgyELX9OOIJbd3fmqXRuE2vhvUURsF9jlp5+CS4+nCJso/ClUkfgNNkOsdGEdN4MpDJhNJPRSkQs
j89jtXaWcAr7/CR4TidyIveYn2MCWlKTWpSPmfmXUlhddJhfiuKBNSMkz1TLgk3YRIjUbtX4t1OT
rH6EAdZvlCrQlaLiEhhla/ka9XbKnYFrJoej1iuVZcQs2xK8otW5vYfRRE6t2HErTnihoGBEDT3c
EGWiK56tsPBjQ5PM0woUMJbPRjknfSa1V0oSAgBPAGRwj/M6Q9vxEhkh8eEL/T/t7A5FWi/G+3OW
pgZVA4SMhQOAMBIWE8qTuSMM1j6XFu7fUcGw0VGn8wZjSX8mHRDKNLFR/OPgeWz0sPnaCTa707fY
X1lXwVhRhIJRg3sTjuTaWeM9AQhmvqHhsh/g7muDHVzPNjORoHfgGQAkTpp9Ri3ZiHsmmp0aITs2
QoGgeZvvKHD7CJnOovl8hk/48UKzHfqlhY52YaqGdIlWYrBuQB0Qdsk4KMwbhzhrws6jhxjkyT6C
Nx7bsZtifXSoJ68IPVEmDyfqTYjnJzDR9qy0TmIT7obPit34m/JJQf0NPDm4smMS6kCUcEb350I0
SFwYvQBIsket9AYzMyxWathZeFKKVc7AIud6W8OWbYaZzsIuBmM6pYz+s8kbkKOAANEVTN7Xu8kk
/nfcTN/2HfDy8wORXZHgBlNCC317g6EhedT/hcENou5LDaEOasXp2n96kcczDI8SyB1DLNRYyJEt
URPbKA7nXGMvgQ0DZBB4f4aqqoe2CMRSBEgm4HrTlpY4dXUJWaZlUlD2oWUWicPOixPhiiHyrQH9
DkCLInLXXOMyg030++ySDAaTVN18/+w+smLGIg3ShbYA8ADNlgkhVZhfGf3Jagqqrs86wxvIk+GC
KsU13HnwjcLjoHwzci5HFxqDga5Z7ha5WERuHY+Uf4+a4CJsAHXIpKs2jQ0JH44x5Gyq1ZwvYVne
3FSETMxNfeEXMXVcTuwczVCBokU1cnBBkfQ2n7tmxOFNo2R8Sv/+IpO9ecf3qSbOnetA/WXankgC
VG1dz0d55fPxxij1Xwj94/q3bWLrrLBP+mbNSR1SdSVsX7xeFLQXmX5vNReR/VT/VsRtR1Z/HYj7
W9JrXY/Sw8SvnxgJ/b0WkYZene0X0cUa9NSeQi/s5x0bncBjdFgqF9tUKKT6niOYAe3hwemF1gnD
5mXbwQ+8gBleZKg4lWrEU5jjzywtNNi2EEnxLX7t6Rihq1+vipw9lLobdlhnEwBT/XTRAl6SKonz
JrM5W4dSUDbczu1P0gt6B27wqipC9foT5SX621rOlo+cFlFhsJ1diMEI6DRd6U8EI14lxSZPWEBY
W67flnKSE61E9sm6odyDclSjLjywimFwMKXvanm2y5hJk1e6FGIZxnyaYOaErrMJ/WJjlNhpJ8/6
3GJ+4Od7hxMLttRM7HHCvC6GaVehKQv2AGjNiqmoSFfbOW/WYKM0VqzNH6o6t7aahzs56MR2jyHL
/0+tjU3bOudCcdeFQwrNx1lxYqqsgMOH+Qw6p87PdCk13/LHBymoeIk3pTj3d8n1K7dGFHnbekW5
xp0A7lLqOd6mQ+A5bdu9dP5RGuhLsDOOka0zUO00zMG25LS68Fk6UrK8wk0HXlcSdl3uzjL1xBsL
p5+sPMYMKJNVx6kulLZvwy3JQ6N2t0XBlx/OsvNBNzLDg2D9pDg8Wbst1WatCsmrn4TOBzK7YN1d
JiYm6T0kFf4SMHiD1QOgw9HXn/FTT+Rp0bxK94+B/42XPpEJjEPP2+BxC3vpEB7PWSz+DWfqFzqR
lPUXD7ZbVlEfW402n7lhfmo/eB3okKkeEdr/szzUhzywidD77h9wf0so16YGokd6QTWQl/gaCPej
LCdP0UkzJlh8kvN7/FfYhi4PK43mU2zYd4l+PfGNrIqpH0fJTElHrJjKYYE3JbhqWW/J+DB25wec
IJ3bmo+xsKHloWqwKT1ndPJWvUaeC/djrX3VT50DkgiwS8nYwEueIZOmso4k7wmH058rgBkbiCIj
DNutns7OkNHCKYXrn7Tf+cG/RaUylYY+tZu2UCN450XRyrlrxEdY0PPwUE9uvROKUHGgJvLR4rRM
MadVFH7AyPZbp7q123sWgw4tiij2wZNcYV/Tw30X+g57Y49cMh04Y8PSu1nhy2bLdMm8JEqWMy6E
5vAkjBBQkcNZzl2Tv23BvwFD542PCgaN9d5BG+XuyVh/CnAGEMaIkxPNvOcO6SliOuHoe+k/3x9U
DbYFdb57xY9Zi33LXJqFwcCLr3DYy38s8qqmaQged0w6fImg54LFyPJPLq5+fj+5UgHvkOE6i5JM
iH6fvNzsRvlOBnniX1Hnk1uIxrFDAKCtrDz0jrmI9ij6v3R1/vlvoh7QcpJRaFQqPWY2afGPh1Ml
YF/v0eJPxUNvS9PTZUYwzgxX3gR/e9MvnGABYLsVqb9RDDJl1uHkPWDmus44oeAYNnbhgrHmw187
loBUgflBaTIyOBzLhHQtQ7AomoutD+t0ID96/pVvEZ4hy21bt5XtyugkmVIJGgMdf/ftmIG/BW72
92EYSthxdk6Nll41yLo0xK76RSjpDq54PFZEWqiN1qzemLwOQORLl2CSIIplQ2mgMFpOFc2UFVPh
yJ1k/eOnTdX2RmMZfzKp8PevM6thGIwRU4Ujy/1UDQdbxxlNO8u8xGaAE4tTV2lgPd9Pu5z1Il5Y
SAGJXeJum/WSbVEY1VjUtt5/RpGznt9F0LmEmJJiOtc9FuICIvD09vOaYEnkCXEbhuEsi9mi6u2X
UYznn5fWo+yk2Ni/22V6RYUNd1d3kGg2WpZgsQbJBpXBs/bxIoWC3Ew3Qzm0m1rR5rfC3IvBeinC
lg9M0LHBnQZ+Y7x2MPFmH0Z4VDKabnIo+ZQrYfShgGZb2bFBTtZnvlQIksFzrULWGn6TPMq8oSzL
ArLfOt3iS2jxxZ53fQXaHV6+OHFmBiTVsTxKaZiXCjU1ceubkyz1tBtV2LpsbkEtld4eJ5v2+yZ0
RHL8r2ZXgI1jPF65gZyMtzaDLgdFFuqeqpGFILEdDYLMETPF8uqBLJFmxgplLq3kRocuhLTuMOYO
+q3Tr4wB6BYFL5VpqLHMEXa//Kn+IzMs+mOKpCI9QZ9sND5hfLgZ/995HW7Jbg38PtU3QhOhoskW
EHqCXJ61rbmQme1DNshGHr3eBoAegSGD6KTw2FTx0mnCITzjOqmmlU9wyXzfc+izIdbz6xqQYw71
OCxMFehgfpA+olQM/tOmt8VuRMuI5G+Qo0i3hzTvVOtMsGaHZBaQLyO4yBxdSct2Cbrrk9kmyuzI
xGDQheg6/CeeP0xJDLG3SBefeRVdWQSaFBEftC4TJbmqn5QLTFXCq32zlc3VeyHa7SL6t/04RiIi
PvrbszmADCqfu3ZY4faagN7PHCe7XE+CAEyrxMoXDvIdYIO44PrkEV1weHEDaopTbNf7sWvYQJIK
IwkpXTno1mT7KMEFMqt9NQCEJdl0HWpFupM/LvDa6GniJN6w76Z9sJfImzf37B1fBJ/q9Fz+8tZy
KAXvZKSVfaePnXexjHxlXUJVWsgiTiKfx7pIRApQPSmpzo9TnOD0i3d4O4Jrh02wIoxL84oSXQAe
z2wTIvbbU1UvKqmogFnGF/YNfBTKvJqFL2HxMdgcnR6sL0vZe3/5RCr0E3CbNTs2AKDDJOdPhmrZ
bd9SQF5Doep6BV8KddYVJHWNR4dsrmtEe7H9k8K6aKi+mjn06sTOeBHcqZ4UDGLOtnO8Uxm00OHl
sNsfrfQRK/4cMw0Ftf+jYamJQGBdQXRoNfcCrcUnuHF6u7W1BUaP8eL9tDuxqltS5xkayuqcak/y
BFSnF1kGQvFhzPppkEaE5e0hpqJXW46VV7cUFf3W/K2h/5QwfWXGc09u1lBx9au5/mgAybiS2+15
plUtg0dBMWMNlqT0CD8Vi7ny/EZNX0y0FCo1AxZWnTyHPhDTa1/cCriaFMJ/s4pk0H8sa/tu7/bN
Ka03+b8Kyf+smRcYlTG1KqMfCRpQx22PhR366HAQfOIlxWdKh7/lTCUUGhzfycxi0XXC4XLXZeBT
rTJdoHlFlcm62ji66p0g+hALv2bvxzBh7OyoXmGPt0UzwLfS/OpV/To9mhrtiRuyGpn9Ez+EQ17G
OPrIaXqzbD66M8guQ1IhV/p7Pj1BMXfv8qR35NWUIHN4rquGREs+hvMGD9fB9/2nTRM653dY+fG5
NTmgdUqKzkZWrxBB4DrYGpx5paPTLgcQmmENzLb2d8hozH7wCrthhBrY/kDE17O2Kbufsm3TFEPf
5GrTf0JDpZ82yXYMhl/vsyr8gupZMwbMe/7WpUTxZLBLUIUgvZJRdwb7P/A3HZG1AuY3ykSkR6uT
7znqXgFL42ubWEZgJFqS4kIbTSVDBtiGd9FHF68nMRI2jZaMcUTuJk0AIKYDvcmM7vp6D4zr4k4g
kX5TSMKRwFAIWThV7RSzywxahEDMc0jq10VG5YFJ0WxrAJwvme65opI7v8P1yO21GDmo9aWlnxXF
1eIJFDZQg+qBtY/VE1K4p9HylHv647FnESSD8fEpQN5QibfNhmig5xC9fecNMc+RPv2binb/Vgu1
22NUeI1qsbU4kJ80VgRnIPgf23fuZ1lQs0zriVRyL4TUZ611F98EtE7Q1/0Cy9D+gAOt7PNTGQSj
c3rm1LUljlktrqdiAjSKQwaxA4ihAUg6cdes+6YhAoiCop6Xqk8rnWEXNJZ4lT5c4jNWxAhLpI20
OoBJcjgX7MRHbmgL4LH85jsiXoBsyRcEGXmYFKPUzPOkFdhJWyterWp9V+jF/EwBuhL98CocH43P
dEe6G8xwYx50EaihBSJkrSzMqjLNCpRAgdtNb/s8f6g8eVoGZFSIQW6mXMHtKtwoGAhRIXheBFcP
IT307V9lJootuqtcYkQsBDmJhKRb6th5jrDaLaCTH8a8n59tMa85AAzeLFz6SHKizaLIPLtl4BdF
mfn9mL/5OZI43tZgbmvxnLEjnnvDU073wyiUIq76YWnO4kkShcMubk2pROQlX2i25tbIEKFzOorZ
O8bv3RqrPKNTHdrbupXSQqCuR/155/tsdkOYHRpbMWZOQ1gMObNsuOfTubdzCsEN3qy3vw4ECAqp
DHheJo7xe4/a1en2aR44A9/2aZGg3X4XrKC84cLC+WqyW4dXQ7XS6W4VNjRVpY6avIODwTwxKAqw
eHXRQr94H4cqk7FsYpzLb1c4NNpKn2y7tEUM7ZUw9II+ziwgRSdPbku+ZtTzgx0ASx3V6vKfeEIs
nvid6AK/bxpeVQSSjxmlUL5oVYvITSnDfBMlnlcGaeF9MGuGGXJNrA+PvJIItjnRFJ6OHmzgllu0
Eg4CSgDcBxpe9ifRFC8ckdhrEZdbX07CZff5kOC9Ts9Olt01afnMNndP7jGRSk+YqdexgWZq7S8d
HFEtJ5Le4TCy9L6rIj5i8inEHMpzicQM7PUxsIb0hfCMfuID7cjuxZXJA43r7Wwv27z8U8JJ193Z
XyjBzJvuqkkcRRbRw7R04UhDdNJ6C3QwsQTTCXN56/sbiZMoPrJ4VJS3jWrCkSlZUWDq9MNYcE4p
MVgH6PHbAv/8paImeFdxSkyImtoowpDU4N7tjbFN69ovIshP4NZXUhfHhZJl6zcGyGVj/AZCo2IL
rUQG5ZvDKxq5OHBD3T2147cPoxk2FvusLA2HgbZHyMRNXqe6LJYr2a95I/hhTuO7sNpmrQDZhvFC
un4EVei5dBfK3K1dIWty6eQXEa0TdQxQn+X0jGmiCyUrimfsX6Qn5TIurdB7QthlfxXYiCkjCXE+
D9h3WPzTadOVG3Wjcta/FStp/6m6Lb5ULtQcD2mNhbe5sGFJluttB5vMRAeGbrBn79a/3bJZEmBs
dUiqmZdANVVMlYlPjo1GOV1ruQHt3WB5U2rGC31ITkjrH/1IEgZBsIrR92VRLnQwmK+KcjkiYCKe
zAAGy0SqSooFteKPaE6SDOtLfbAOsE+LAmeBQTCaFHAb2jCuWL8/yj+ej+8MkN7rCCG3fLg5XR+D
tdjUJ9FAnhaTH85wjjReL3tAC578142VBQ8Qod0S+PcZNsypLM9+MyKIonJ+YmBw3ZrIORkA3Nbd
6+VVbV764ZHqqo5bZIRKKl239waVthXpIZEvtWzRXpBUz/IZCF0DykRP05tRLN8rpy95gkAPpzlr
VZC/2ip7tN17mbCfWVAFCKsKKCA9j405pGbOdkJMtEUzrO65W0uwKtXIOCpg7oEwJDFVg+ll10wN
KNuSOtl/NS9Xw8Wut+mf037PbA1swI4hqXQGMfMY/QddMaf5fz6JDAq0dRH+cLJAU1kTuB5x0qCh
WangYyOVvFRX3ToEhBLNGDUzP/JDdpRMnrSTfwR6wSyjyfzDXrxE5HR0FAmovgjNTIpTqDVdrBqo
eQKVSbwHnsyNROT7y0ZejGBdeu0/7qXH9Ro1XJDWTdxcrplTHeQeCyoy6G+SdG+jtXxADowKr+PJ
8AzGqD3YZ35bEVtz+5oougRoFG0dPBXKHJTVf0yxP+rmJ+uSrt4jfXnU1HWSQXZ9IQLhebB81uXO
Xm6iKSlv4zIqMmsfdFdWFiuKzsTO0wWU6pq5e3N1wT1VcTLiZq8iJQpupVMHWqyy959AO13gGxJ5
5Z0/Hfi0gPTNUQXHRKlQzxM3yaFfUH1CTpaOFW2MRhvFDwkYOCDbx7Zg/tp/upKgZVPZgBaKf121
jbFMzUoEp2ZLoQNiz2fh4MyN7324n22F+s3ektpY4DJhALIm2/MQH4ju3j4RQbZ5HFf+FzlOTtam
4LMJBSSynRekN6+XZD22AzcZR0BnvF3WUuJQBuAmSbXcUR+rZp8GuZC9p7PJnMkXW5IEQ89UJMyO
eIPDyBKQbr3Ddj8aFFJc1zPNHRNGrYkLB32urFheSpvT/MA9qi9u/jXa29612hDmYwdjoy3LskWW
5ijSukHTQXFWN11XGX1OzJe2cwtDFDeKfBtmlGt4fBiu1imfIsmBK5b03OduwAn9cLpsGVRuIZm9
ydDKizfWwr/mmiSzM516Xr0JHDtJPuemNOYTBsWD27vJIqdSPaGTkDb7psh85HZSN4fzbJcNBx/L
oNW4T+if9Ok5iuw5yPJWqS9jDfbITHLwFkja2Yf7iMqbE+QXLqyXYw3AZpFpXglXcOr1oTXjF0OY
H4vTxad6nGsa5h7GOYaCNy9bR5QTijoiZg/mvIIJ/Gnye6t7qW1Xq9KMdIFps7Tff8uYS4bJrQ9W
7NzIiD/sQqutOXEmyxFNJAvbhg1/JZuGnshx6ffVY5GlBiay+kvgtM//hF7TAjpoGumrWu5n16T/
pBE3mbSt5/PRQlwfdV6n49q/iEcJUn/FLZ2tAIlb4vu5a8Ge0JDvdocnT1NJk8RMOQWqjqYsq0wL
Wu4Ysr/G9y1juLRhKiy74+2AY2OSuophsx/qPxuX3IzErOjmsNNfXM1yLCdpvFxPg4BFvCzUvZkn
bzmaafWZsjykhWqmCZcwjahJdn5UmcxAzUAi8RHakynz0hGDFPfltQ05R2dT1a++SfQg6+7eFpic
2V5dMXSecF+bBGZ719u0TwwrPkz2XTRuGdXOzvFDg7Oh/4YnrqiU8WC4Bw24ZHetCRQKqXV/6I4I
lEtZdeFkB4ef3/G567i+bDa8Jnw3xMbkMp4yR0iOi/wSgLtLEaeS3iEcyaEsvRRFRZhekw+ctRk7
U5o+IgOAa1JJynSnM3KIHccUU71D/Lq4s3IyC0hwtHe5OOHEw8IzOiDOxJeZtkFsMB5qcx92SG/1
30S5NZ6JBx7xXiBhHg1kk2tFfBhOiE2XoiGTVPxtSOqDw9uS6Bk3vY8ASPLASkC1ZoG1byMPGibK
p+oJEhZTZxctUPzRF0K8tL+B/yu8r4pLlWG93kpcGoJfbOgFrC2ivHGxhUrHyOD3CtgqlshtqoGF
p8hMq3uHp2rFJtu60YtiqN2ehnDvN7jaCtmXjQ32wU224WUtIbBxEVAwlYLhRW2vwimaA79VW5c8
+otgKahoYtpBy+TdJiV71SCIpEnm7tkLZHsq03v7v1n7DkVITV78Py6ImuEccx63/uxXG4o4VNdL
QcTppqak3XwP6QtR6vlNBOhy5nlPvS4baJxoBzYPsd9PpqB6LqLhyslaBXpuCYV4lFxWMVeQsyY+
5+JCUGSss0tYYteXdo8q5ZeFjlfFZjnFUE0+1t/9KNsvD5ebVaRUvCJ9eJypCMBk2zEdWong3c/K
y4xhTw/NFGJucJlxBMsoZNYg7W3aK5vGobpKZeiGdFKTE2lH/BOT+It5rvRq7ZwyyRAQCz4JG+VJ
7J7H8rnVHR8Htj+OFzxmpsZNOzWjTBh5CDL8XrL9wOZWvnUROHahd3AhCSDlFeytXXNilmEQupBX
2o322DHddGR0bZe26MwlbyCtzqh9Bh08MXFuiG70b5L3mP3t9A73rGOHgpjLN7dGySjOgDxVfChU
vho0xwf5HCUBU3GSv9ztS3GhQGG30JKhpR6kI3JTkJj/xOvpCHs7ptv/NIuLgEcuGLWiuwk8ifPq
iu8hxzNfxzFqP6jIXwxNEtAeAoQEWLFfTLCChIlcWC+vDL0IshFcR3FM8qRsSC4eketoCu4VRdty
rMSMOl1BS2GshFoUVyp7xDxBHDUNVVGHlF8KFiWVnDGjsbrXOrdrc/XQmZ6o1ZRRINjEf+EqAAud
F6FQ6rANM4QfoSyvWJjvbzVJOdixnQNMvVHHec6SMTzugo2QXmnwA3IQAZDzbzbvpsn3Ypv3a0hw
eXW9sJeNaTNHNw3zNyCT+N3hUNc1BtUAPN/VC8bZFaSvfWVLeh+RVRLoE5Va04lrBqEpG0lMl3IR
qDdf5x9crExm9XCcFgtI7h/Fijtb2oUiCYAevBMBDaPkDOj1fcwD7kVC0F5ErtAb7gifGM8UUF+f
oWB/ZGQdGCXTkqgk/G+4jY6iaMjX16F3wTKNyI5BuvLDP7lUeT067FiBH5gKZSV+vyJrBKaQHu9w
l/IThEjo/Id0cStLvvLh8bXlenqDQhtjtvx+fZFe+FiFpBkL3WCoB5SAQ6bOBrdtz5RDnPc6klpJ
XiS9rOFPYm/GWkSU6vb2ZjaIJAJy72nkxHRxG9Cd8ML970UUFxoAqB8PTTXc7Lk3EeoHTuv810kG
c0aXg+Ir4wXyWCvXKXZwfoifizLH9NB/O/oRd4A4Jn6QJIhBtKLHgpea7NOgSlxd/5+V09+AM+YM
gMR961Gw6ui00t5CxbRkjMYcj3fUVbNd3h15cxND4LtvcModc7sQJIvZGmmO2ebbGP6Q46OJZphk
burCMQiyZMXsmy3gJ79sx/sfi7dkamdCJP5OUCuDDJZeM4yDPWdXRUwm0wl8O7fMPVo1Y6pPnBk6
rBWT/fnes/m88gHzKwkJHhJ3dBUgXI54bq2Z+pksLQXUyXSP/iKpUa61agYAsMBZe4RgaNjobsaz
HURm54KQ4P20aTjaxl6zynezozX68RMtOEsFgLYvi42pu3Ka5Dg/l66UWkWFPnLFdv+IUpXbM2N9
WL5G2O/7d6rhT0YyLefElK71R0jzR3XD4ahkan/tKGimmzOr2E5sKWgzVuam73FZsTqVlTlG1S53
BINdYEF9iqOzyEpBxWxD+sK/CnNn5MViuj6I/ZP01THlltWzyoA+2cmCTCq9BYaUC+DcBWHlUxMk
Bsg/S6AqOtmrHkfgIWix8l+pYFUQ9foNhMqBQuvbcH4PGHSuGPifl97OYU/QB38tfXvPrqyoSaS2
cjVpbZWIWGcejyY5nxSwM8JFsI0xN6jNwTfYbmWcouqosVOkslBNqQmHYepA6juJuTk2ckheJP6y
zGaoCpX/ZmlN7sK5VIPFOx/rVBmUAWCd/jX3pQgAYxZDu5K0dlhRX/N/qGEvTTq+x80oCbebxIo/
/AxYLQhidDCM/Z/DtySyPDv3fYpx+pF+atr2knw5BFMG4Z+zyVh2XpRg9/Zk2/uc8SRZUuTGhld2
cI+UMNX5ReaTATmOkWzOKPx1CrM/u05dYK06d9qpbWb7C2WD0hWVMz9k5Krf25ErI1QZkUw7mAl1
+HtMvq10icRW/sEAeXhS1TdEmcYSA2rSNkVMijL3hSsfcs/tUXnByuO7YvUScnwIaZ5R0TImTlmK
tBaSgUqW2N0YPL6m6JbrFWp0FkoCi22Rd3/SXvqax2PvDFsIUWmrBZkvrR32lP5WuCAJ2JbDg/lC
nojfvztrnohLwEmHGL1Z7GgLNCgTb6hb8znz9CGjg1ByLHRfzeDtXjbdAHzNy+cHHHuQhx9FFec3
pHSGvU7j6lDte+ZJ/jgieBfNg3wb+cLnLM1MTv05CXCwUtc+tYel2ArDUzjgqqetqnECggqnoJFg
Ovz/hZIGI5XrqZlBtRJvDJGyA7zukJZ1VVcPYtfePgzjumuvhEjQN3Al57KXWmjpJYjwfrLo8IjC
dQdDkQ5fYHc8I6zBrBvvtRy9FtWySMd6osQurZsb8QU18vwd04mmcN/0jKrKzpRJHS6CH9J6Cffm
4p2M5jyCRC42rXFLzVIdGYmczmkY/roizsi+zjnsJD+DTX4m7UJTUZ8GHUioD3iTxpcD6AZdcWC2
F+0I4uorYqOe+G1YQZ0kFD6gLomuYw+LmrWzFwJZ3cmP5JhtXE4bzEYgDceDxALDGPpUz++YBXZz
PbGaiKk+FytOmRw4QMepJF66Y+SN98wq+rwu7REFK4rsLqk+fniwVaDa0j4RsIQ7jX5e6eUVCkBp
QvW+tK09tx4OaZkGqZSXtTEB6RfNgf03XBJs6tbw+QyA00HLV3j7viSHVUtG4NTa6lpNA1BmzHm1
4nBKjXxs6TMcbf4h2mWJm4QT4ecMfLWNjhUkAQLOrytFyWo9oeW64/x98WtnpmHfqh7ooDziRS0x
F2giaki7VpysvjX7TRsOUl/ujUGZ9v/7lU4SFnkVQ/xT9Bnx6iQM/lXPr8T18OR0vedAQY48Q7vI
AcQpctZ5Anve3LgL2AJcY2rkzYZSNCnV089Cwd9dvPNWiD2HEN/a8Asa5fFBhXO5kdsXxg41zE9w
3AU/LnJwofbXNbLpY+N5QOINqJC9Vmp2Itv0AxRcEo3yXqHwkb6igLLBjhxXtet+NnccYYoKsLpb
DIaEMh6dBNmYq73I30hnTM7rE1s1MmHYQVsKi3ikaXzQAUCO/fqRTousuydhkChiGsY8CCNwnx2d
ek+P4MVmhzjalslcAsASJ3blo6UNZwkx7OAGjeS2mlv32RBs9G0SNUqhzXgB/gla5h0rsljs1tWB
/OpcqSDckheYfxiTrAqVl+7LbkUnYbxeo7CzWvutgRfBZt9CkulPdM92+g/NnrP7PnbAXRpXgDz0
AHifXy/o8AFuqGqloxOn6ekdh8N5cBMdFhc8iI6CrAKKWRlY+76hJoTuZKQvIb/Hqe72uYFJsL+6
7RdTqBNu1LfTG+yfuxyPbbukigF2hHNnTjcQ72Qyj0wTMMHaQZ+k/iy+yHxE4aZd4PxEZ5Pd5Cgl
zPk0ghcwmWvTpjPNbUYuYUydc5C2Ny1GXQWULH9Ia3RDRv5pPt0/ge3smbpcARa4PZEPYHgHyRQP
UG/bo2FARjupsrNgjOw+7SiauxDp4JFqBnBhE7b9RuYMdJ5GYXP2ItjsY/ymnejIkJPVjbB4APQj
mno4iJsSze5rALS9MrK3IdkvjAvIa18EaiWpz1jTpFJ866StnD7PuZZ+8hu54TSujQm3XDq5pTMB
l2UcrxjlRIH/KfRYtTM1upd8YhV0nanaXvTeBFPrnfVEqAKLvBYvbiACMzkcTdipHF8TAmJfpl2k
ElCgGh04uyM+PU6dEJ4AY79PN9/cLbgKI/AEJVY8ll/AVUYAVQmYzGMpDZltFcRAMwk921lTw+DH
hckKbBxDAkKrwGgoPXduLhi4TqOBBCTnvIsCt2H9/JuKgi0ao3t+KJTqqY7Ivd/LwRsnNC1BclH7
dYPTXNmv4gUrJ6AWp3JEJ4Bo72AL6sU8zYYISiVKawHXjMDmIHUzrgED7zvQmbrd5sCdZm3SzoBf
BF4TrejmMx7YMHkDHTo8uXjwS/jQJ/fEavZIUDd+O7zxDKkitZyIeWep2r8vvB6wU3eiYz3yoV66
Fw/FMeY8/A8m/pF5ug28iD4U+0A3owjrfvkcpXv/HWSKPGIKjFNF7syrakOmH0ZncMQUsLiWEqFR
Wd4XHqgQ7WqN+AWim2I1cBfoWOfBkwe1e2WL/kXKTheucmNOnvz1zg7rkuQhMfz42/z5ANX6iqq7
uDiJnM7aX6zmH9LXAI9UGicYcVoihOrXNMbqEOSp98lrJekWnzgOObkpB80dknChMAwJZYmgimU5
7d5KdPIo3s0BEnqI/wL8e2lWWomspPkH7Z2tEcoQYOCqiZzUY0kM9VfacqVfHrQ8vlo3WroNDcTv
CJVYn4Cv6cjJ5MBaaHI8AzDpVKmg2EWczYMow/xPEPU/Z+VWbHW8zV9qL3YWoViUkmVZTUOgj/OG
FLfn9UNH/WQSfwDRRivHqIL2W4vhL1qj7KftCz5bOKB1WXoZbyyof+geK+wraymCU1p4PCHDzSGa
G6e1bU16Vv5NLScOFhykPjTJeo4wHPcHW+WtCVbpYsh2qgKcckRwVIZVJNmVaanlxUAGI7q0i5+s
BmkEWhNw33XU7pT40ejXmdcTxkAwqPoNjQlODZ43rxxfv9Q47XzKz3YKtmbMZ4cLetQ4NZrPB8Lr
OgCDDnsAklr+LZ5LUiD2jI3hh8mCKBoy/iqsxRjoAMfWD14Ov1DE9gKqrZC4oHQZLcaskbhjPFq/
Z88XrqUfDrC84yt8xverkYJx9QxBM+1KjlJbcI7gyfN3iMwUgb8QzRcVVZMiLMJsyqpZkJTQdLrt
HuLfOIDnGH6hrWliNkTipjEI5gdx/wQyXZo0BiSqIHoIKbQBKLMLpGsT4BbQrOJW7cfRoOyadieG
a76F55QwuckKPfX0pO3Fl90mERFGc3pekLxk1WiCMMabtLFZ0sHla2oNy8ZCHS2pSrsVpc4rU4vQ
sLvTeuZoPR5F6tp9Rgyjap7oRjyZiX3P/MMe3QjJaROS+M2CMGBY29yoeJNwNZE2g982cd/fyaPz
SYrsEPQ37u0zIH0MozdMuXQ1H2JZklHRHdTOpoKqkFFgSqEY5YCjgGYUqENpQ9NY2U6Zw7tvYf7J
lCeyI8oGZj/uv8tptWdG5n4s3aXfl5yYBvxi1Q73lO3X++jq+0f50AXnXbGr9mtybaV+M2QfQr3j
tkbeoBoaw5oSyqx6Zvj9VAGh87aliOH5+wZ+h1m1PfUovxfpAh8tMHpLbifXAjWYqXmuZtxEnOtC
H6rzwSrDyTy8ycdF7/B9aYeDAC7/tun6tJA3lQRVwTa1w2zBhSr9rQqe1Fky/TtxFLh/CuxFpYND
2n4P65ZWpRQiwRlgB3AbfzJBj/t9OJpSzJ3oolT4nVVns4fGObtulUI4GkfQU45PRqp9YOWmjTi7
inB8Ve3wushrZ4KhOcxK3g8ScAxpPYokTpLmZJop9yfBJ1njSOiTKau3SYJZi3YiFMDo6rItZAS2
CDB7MPvaKzrDrxNklYVfMcwalG8/QwJjpQ1bJLkD7SBkZd3cmYHnnv/axuIuZDy3vfaqJMr0WTCL
xFcxbFGuNUT62aj/r6B8FOws+QqO9WK7UpZd+qP/Ma3uOBfxS12DAkRnfK0R0R1Ty2BRJzeew/aA
kaQ+gOtnha0HkUz3124HEgBRNi24JA9qCOGMfC862kAPkftzZ1H6bbbdDjeSVhsR+oduy5LW9w/t
y67WUPDiPY27o0NEENKB2ukUe2QXIpyYRBhwJESxyIeJUXNqWzTi4eFLwjHujBRwOVdbLhnyLd6q
+UIa/MeBC8RpFxOfpCDD2vWI0Yhm8N0l5yiVaEGOo0UeEAN1TAoYYfc+Faoa2lBIai7rDMPv+Vaw
JWd0dHZzmPpKJjtjyz/hw4am/IcF0m2tWu1o1bAe7SCNj8fZ6LIOgLLPk0T1nwkalxoRf2UKKORq
4qIXCEykmIMijMbsU0B52m2al9Bg1tZbpx8rW3tk8BoatBMjanNzwLWwyXGu6iO8W5kAnKLkFRXA
ldk6GrKhhpzUQ4yhsovl6k/6YYNwtBNcbHbOWjtnd7ML4MFO2JrT/3praJzOpX7MLLNrM68GwDvt
4J7nC7uhh27kp6OwX2T8JzXI6AmZyj5O9ujdvBqxHqmQ3IL+VFjxl/L576tg7UB3i7xaQBVzCtH5
ekJOZ40zFoY1lnxKmKsPdGZbqZUZFgTZEwdnKFyrUEUAG/a3Pk0VRQt/oLggQ9H7A3BPrxrufEer
dEmzwbhHl3GZXSKA2SOpOVzRzOjYyYat12JzCvDVzNCZojdjp8JFuv6HmEIEek5Zx7XjeVDaA/yl
nAuhmJ/ex7n5f4jzl0CMgEyfgHaAV9+OhyqKIFOS28Ej73jhrpxGoW5Z5IQHMOGb3YkzvIwTtNZW
YzgKPLeXzTsGFpaW1F4Plafu1qyaAGTefdJ3QefgdEcMgdSbkJ5UFZveAXf+KsMDTTXuKJ685QuB
swpBZx5Rt/he3h36yrzImVbsMx1V3bYwB6bCwRtiIVAmRu5QkjiHZbrNBzxJJb2F/RVWyLgLrxyu
iBC3m3bjko145eQMlFBuijFx5wwWlGzDT35ppkfk5G/uOiVrHUNFKSB/4i6rViHoZCTWHrGdvWfT
3fcQrue67JdHFmvku7EqQ7csuJHf2IjPkM5LqTXJPX0EhAIEeHiW3UbKEf0dthBlNDHrDvuCA1xp
7oBITnwgaxADlKp5JxeBSNEq4rzA/cls/z3w+lhj5hJiNXxI1LdoTbuQVRQtwaKrr7ED/AWL1diQ
2j5Y7fBR8NvC0DSm5yJw2i1LeKWuLrL1iLoF5FF+2UesoQsx+TzZPTZPRlHQuivBsgViSOHetQGa
UddzM2RjiZxdNUVIBTAOvpx6QfWCZlpSjOL9pom+SZvQPyLBXkr/FKQWyL5DXG5cHwUcjStosbG6
mI9mFBUvEHeBGkPnCmWCvUm43wmAUpz5FXKVwnq4NbneKBk4G7PKvbvVmwi/aQsWBA2tUi7MbJor
bz/aslrDg62Yg8lUfdYXTIDj1x7DjxiP0TTCDHc6h07jT1Ad5dqBq9IKXzJ1XKTIkr/P+G3wkAMx
zv1ct5p/pZn4IYJ4KZAHfVm/LcLHX2zHFqjWnmeeY2rgqyclAa3mk/FFtin1uyGsr7Ahu0GGxaGT
uxSoc7BYAtsvp3Wpq9wGMK7yVFsspG5MbTJhPH7gJHkIKIPodU21nilPHwbw469uCtsjtB5pwtPb
Ga/ae47ptuLk0vTRFcfX4/bfuXdRN1QIVf4AWOVLzIz2vfU9AXE2RewBL1XSUdYrqUazXyJqVGrs
1YUNoW+pOBD8y8eM8mvzpmTldjdYJgem6ePOYSK5aO9TOxJ16jFNyR/kG/h2pKCWtpvFJxnffJyE
W6DzwNPUCHmGTrJ7D7YxK7eXlqcCz8jQBzW/5iFKD+w2UPaXM+GKN8ufISu0wWQIwVFtXgW8Zz7b
jh0K7lYYrOf1XMuE0eBxUeiLyew1WBKYVCR5R7J+1H2/lPJaQUmAREsXeC4a8KuSuGpGS2lOAsfR
FSZbUJrMDfdhNAnRidDNuQrXloZptXu6INLgEkPE/ucnyfv40+42j9S5CvMWN5E3cz1H26ipBs2j
CfUxwANKjuEixctLmyqejR3ya0dIXLVt1O1u7wPwppm4qQtHRy3J7uAetxKRj3jxzMrE/kjrf1n2
8v/d4QGS6wDsEgXKbfLGby2UEt7U1wF+copVCotxX0XGEnir5W2cZ9bZWAcxkWxVQbDgiyGVFKPe
+jSXqfFs8vf1gnPSp4J+fqESUdPfoGRc0F89VmHlRHeILfrRvjnchClt9sEof9WWoUhxahvGl4uX
vk8fOvLIzWzK7umACPN8M+wv//SG6AxdMeIDrrcMY8CQqR43+aw0aGIxidS+Pofw0rcY1AJd6alY
/mw3CLa29zZ7ihZV2IkmksczeoYdDj4LgnqdjtVlM+gMC29cmUbHlw+/N50mXlBVM7eNKpsyfjuQ
n5aKJHw3rAM0Khb5okxO2RmLfgPDzin5kUezDe6do3KsMuTQmMgk3zm+lCuRW248GPZcUuuxJl/s
dKuS9dWtFZNQxDAE2M8fNfPUoEeJAmIeWlfmEm8jzctJmITDxdsnmO0HVA015czFr1TvmNNSfn0M
gJ4xvmhMzKAzIAn1lAD7TfUlPRBQ9gA2R9a4iQvKh7QcY5m2Slg7WSvzS4fD1R3AMHVjSzzoQSI3
bnXcMTTn6m39P04ni7TltmDPuxpEraEQg6gLEpwTEjtaJ9V/+Zu3tDPjD3MHS7ZjWINu3cDFd3wO
UX3HUYFT2z/MMXKjEMUK2JHG/P5miQTFWE84OblMWlUyYT+1dtcRgbWRfxG7HRFuG9wYIClwXB1J
Zv6MlYxbgruvydn1fo0dWt0eSmWtNRfTqxJbBRP5BqHxeeE8OZ7uB45O5dwuvR0PIiFYwSzDwfBP
J77tJfLAqoa9guSo9gsn1eHloQorb3xoFFFwYEJITS88Xx0dAIXs7huThnPTdOQt29UIcVqSLx99
1zi3oPUisXYF+VSoKnTx9G7m0F5PnA3e3+WxgmnWJ6zVk3yerph4sS/K81xOFjiah5EohIagXSzZ
fH9FZ+r39/Xk6H9SOZ9Xl9gxdSbEgg1GGEXVPHCG81tApMvsQvg7WmoIE1u2f1ErKRxUEKlGtinR
y13TAJ5+vd3eR15++grtcpyFOthW5mZhYB2CU3637j1hQDnuBLSwXMUrV8SnYjesCJgx0qPTS357
zgvDthYNUt6iWFSgOSdt5jiKyTsTCYzVYhy8P75hfR21Iwd/t2J3ZnclpxCiwRT3fJuWlBypfX0L
nDzBtrZtxgmkyKJ3aKgFNzPIZesHm5Oyi0JII+53NmtyB4tN4fKnGLFfESRruJH2VnTcGOd4wpG8
EICtVgH1xBMESLG77bxa5vkHvwqThCvEuoN0gSfW1V/n3TdGN/W9CsOATVPeOfokDrs63aCsVxB9
NHOHRkoUHnR4gny/Y/M9kGZz3XXJ6iPGhmHdD8nzrIIrwXG2CocyGkEmIAiDolcC6GCeliDvQ1ho
3GP6ULjYekWLNgy/cUtpUzWwbHVBodypIPzoewmmn/eqIF6MbqMInLMaOEhT58oNjxFrRuroBQAx
i0OZcXD3K5gpYJS2wvrWBCwZZ0+HvJMqKs3rQmBucRGov8APilHWtHvL5gWR0cNxBthI4N8p8Cfx
JhiqTcCN1L87LYete9l5+CZzT/YcNyuM9oEys3MmOEw1kYLxFh2mPw0WXdg0Jh63IHzDB3YWitb2
TR+PjPq1rKV8kPQaX9f/sUMJ0BVBCtXC0e8HE3IfulsumbO3blWEnMm6UEiOEZdAAFiBz53AwyxL
0d9jNYiMSai1rMG68rRAK35n31LWwHT13hfTuLTGSVyKFbTL9Nz2dWXOLGXgI+7CZKiDlJ09Te8X
2FvibBYHm9rGAYsEebHxSFWUwvTYeyMg3K2/X6AsosCv79rHF0qty/aJpdpSMbZ8nA6vaWbvvc4A
GH5fMxQUS8kxi1RmCSlYHzmd31fZNKlmPFFLvDUOz60D1xsXJ4+ImHX/vQUgz6mycG9+BA6Zljck
TCV7J1gShPW2x7/Ye2HEl3xHdmZ1e6KqwLGH5fBxNKDEL+XEIgdsn44/SpcK089HUVBXJs53m3xf
96N2bjztPLgpAiMmuSmOYKAKPqsm87kfdWA9MdFSLx20cybMgMkdXE/MojgQDT/P2xdcKDR5xKze
erBE6OGnIU/5kiT6+5DEdthJbNoDe9IPBxN0QsVbQVc0SZcSJSQap+Jd51eXsCzpbPzMMWfGl51z
rGt9Gxax4T0xHTl8C4KLApWEKLk11i2HbN6Ts3uPzQbxEOtlaZJQBBvdabkXKTrj9OlVa0LkXcay
cXYAOpyRwuYQ3WytzUenKMAt+Tlk6QBKTpRbnJ8bIsFh1e+QAvToZ6Np8Qi2/XRGFL8K3lrNcCz6
1Vb2TJyCfka6gXzaSSa94sc1qpmjt9MxLJdb2tDCOmazkO0vXEjVi/aueXbABQCKqhEtHyK4Fqp6
EPHIv+fn8Sxeoq0U9TCLTQ3TK+2S9J9cPzKqM6r82dE5aWKgSV9hgcSQBLQnoBwaafnQmPxuHvr2
RlBfwA0l7UnGZUazf5bpThu0HDicr1I3z42Au/O9G4HD6OG8Jicxempn1Lc7GEc/bGfNK+RE2e5J
DCXgjT61wsZxe+j/r6aQM6E18TutyDFx68RKAl7MbPh3SdwR9TVn6gTFs/bCkNcf+q5V9UOXFmEx
Ye61OdQBE6kiTviOlRd1QtHQBwUA9PX2D+yV8KcBujw3uCvFMtZCjJlt2nUcMibSwHEbnSLiXMI1
bwvqM5qZ82FiPZ6NpzpuUflDTNMt02cc/gv6OREEsDDiKpWmum+8uoNTLdygiEjhv6tzZYNIt6Xr
DyI3FwXN7BgaQHsNzGqk5gbF1w+YI309Js3VYxtPgYcuRiyEgiAFeZBb1PCZyk71bmxHEaf4bZZb
4Ar/Nf5ev37MYvrCwZqlMqVhOxSobpQ+1GG2df5aCDJcvdWT+LysYQZ9o4sfugiBdI6+SGrqOr05
23ncCodtbhAMB/59TI3iRh5eBwu0U5MgTdyU7wNbDZibh+1I222n5Wg0B7URCTAT87BUFahcC/zW
jp/1xdJuA0g2V2TO1CGAp/Q5zvr7mkqmh/uir3ul6Et6ypSWNdi3SNzk/v/J8/1mvbIAz0UClNcj
1I5CchS0uMlBlR9H8VC7PQJfjAAKTdM/ND4/WDnw6PUaT8e5xuuOPhA2rBQbYPjhyxTrRehK6hzq
aX7/lJeXjDg1sL5iV+1TfddxSwF6sM5ZnUkwsdIqOf04DrH0qyezVUIlieZi/5KgkXl3Ow3FMPY4
wnxgOOL0fP9pNzi6foz6yR0yvFDfvpB29VgpEG5zMcweKK6ik6UoNSY7KDJbz5Sc6NOg1ujE1u1G
50wuyl7qpgUq+m3JWAYWNXlINZbDDm6PQwSnlSTke6+IXL8P+gxY0taHu8jEtMP4QRDAyzjmOUns
RCUsO495zd1BjyZldZnKBxBwhR2ODw5rC3zzDV7idGgHJMA8c8yMq0N4Pv/Qnr0Z4979kgf+w4bV
yBFPOLl1qozKy7s37c5zYa1iJAtOxVbZFgJg90Nsi/xVjEBxY8v3PQeG41rZXqCeAHZF2Ej4eOtn
HQ0PU60mgrupZjOp2rV1zknYuVPrldvqxPRwtsShx3t2pUSqBT8pesEmud62Xgffahs4DyT37wAG
+SccgwmsLu+PIfbqUuzrIIDj3Je6EvIplN0XEpPu5bVAUP+us/DNXuFq5CC9ITRUQQDsYAT5DVzV
Ni7WYsrNLNnQPiN4nnzqPs2rhLkrzcbLtOONOJ4kHGvYIXIl511yDGSrMa33tkUCrqYpbdI+WRum
wEtaky5pUNqO4dUiWHjQab+wpDTcidOyZ3gfaTvnFqlcaMQ/y1mo3rDCnRWMB78LkFbvvRyK4Vid
0dAt07R9uMZkipIkJ2x5pYWAnqgcvPwbtU9yTYpXIUfJu1U1ZtNuWrWAb6QMoLGwUQMoAyqGYh/A
ioN1MfTtFIvZH9N3k5KUPEz4gSGnHKaL8GRTU0UbpePavP0Ol9GPAj9GvyovlADXEinIelI6tolw
lJY+7esBLeOy5+IoJz7ncA0mkvmFowSfDumwudiQNl4jBZcvdOdkkMxR+tYBDd7g+lFFrXSdbJa8
iFc3DgHkR45We4hR7fXgaP3jLqpHhq4tKBI6ik8TyitV8GqB9xjD+bpA05OgDskpw1b5MrHcXf8L
oO6ZCrLM9GzJIeRFZcgROFacMGyW+GBQ3fh6AYluWcbLC8s+Ptl20VJ45VINvqPxC02wnQdb45xG
OD1bRx3dyzjKqwRKYwBjAkjHpuqPNQLEc55IOuN7J2m57Ibt8MDnQWHZUVYnyVNlZ2Lf44yWIiVL
orEsrVWVsVlGN9TzBqMRoyw8+jEhUOnaY81XG3B3ldCY1UzAS1xLudPmmpZpJxPdZDqpheaRo8kk
DLdJoc9A4v43ulfo1C0uCw2841LpnE7mKJZeaf+sjDYl4nYlezwvehmsL8ggWJaaofplc1ry+HZY
b1563TML0JXkzI6PFfVy+1dYpAR6HlYiM5XF8ja5jsQj4WPQ4MSrA2TSyUa9Cn/IuuGEieXMRdLW
M8HRq/dEf5DNhVuTwTbwcTWAb6ZXlXmFmYNDDChsT3DYViITBIcP8jrlq5eGxfrcrTHdt5bIAaxq
aj6vXdMyeNwfjetNOFC5fa5TbEX85UGdvzMKMKHFm7q2/eJ8QhS/IL4PNK+houmt6S6ZYkh0Rj5x
gKS6vwnjfcq0MF0CZyq1czLWWPkNGuwwG7lcC538Dz3sNyq8x2na2zj8z4CVmmferb01InsufS6B
+vMQYXH4/n+fENpAWVCykDWNvGU3SiLEQAEH4G9OBUzB2vYw/m9wjs5V49NrNKLL0VpffmJ5yTRR
ofQrrV/VdfHoLZaDfAR46kC880azWCkHWI1mg0XH9wOL9nijMqUCTP/W3lPDfC9iQurHhGbCxbKL
7HbKyGNS17jzSGx/2kL2jp4JKp6JCtCVIwrZPQy8SiEXS0gliFavmhSSSLzLfEMVCvNqBjxvNgvI
HAg3lfZNhh6ytmKMif/nlF0fvsinOHFNMH4zLL4z5e3vS2WvyGDYyejepYD4jFQBKIb024omTZWn
hUvJkOY1AOShQpJ6EnrHohvP/A0/v5YusqbZg+L3svGw6l00I8fuYZdhmEu35IiqZvw5mZsIzwMs
Nlfgsfc8FawkyvmeQxVlSmYpJFKDJxHxtgcxRz4iZ7ktJrVykOjaGG48QiGVwqBJxoYVDv21qryv
H0dIZrzNZiV6rJribBQw1RCODECQWV0qD+zNeqmdlBo8hCBfSBPcPuY/ujBoVobjq2z48iYdcpV+
oZF2DoHCNqugb3GTLxtnS4shGtDx4b29+SrXJkdtQnVLBUjw0LVZpSfIeD6myeOnodvLY5rhW+3A
UgekZrKrUvg7clwhHwDDDbkFLhT5HNpazVxQIp5Qfq0MknKrOOb7ICz0Y5w3KJQBF/2kcXEpoGE7
9hgwtV8vzPu/Jb311Q0mA+z+5wkrljMwceWDG7RgExqv3wuaP/3XaBuGwkyq3atUG6Fb1C97gHfW
TH1+dbznDx/hz1mIQLXbAndi0FYkCE2VDOMlzZ+FpsiE8Yahxy1V6iFnXBiiqmGOWpzCYCXCWb1K
y0smbQ257O3XkA2KpDLBn6gtI6xxPgik0MZXAfKRc12TNPt0NeJG1vF14c20lOngKOLsfQbv3e1h
MguXC87XLBvx5JRPeowseJfNZtOINFboFrlgjBGNF/QSkrFMl/3B+gdCoe50HE9/Ehg6KwwsR1/j
yvbOeQlRZz8xMSYnFQ2kVf4Dg5Ps8Vcik/Nuc224lsTeFiW7meoB/lVVEl38B/6T1cDenHAlsDAZ
LLPKFlZXvbK+tbLa5Ai8cb5f/J7ajQ/RG8UJfYItGc33j4XnxrRdSSO6uS/F+XmUmrOsHRzbaZln
RTSH9bBxJDhP3zSgwidVJ00h9AtWN8b9AcdzrQfEcxrsragDIAZStg9I2Xc+bz4jLL8fVSHwK/kW
HOUAaA8DWveeMZGHKluLB3+EIE1H4GCclTO7XIF26BWJV3cBdBsrCWsiW09+WxQnneqY8xQaa09/
b+II58SVCCQoaoYMf+3bMJMgKhRtm8PrQ5hp+qX5OD2Es681hNbenpvK4kMpALYaMXx4YX1eLUFM
iM78/ovCMdpkf3DabouTMMfC9eajr8hF6KiChKU0Voab18LAn7Q4V1eOamB1MN5UpT9WbnTWVdK9
a/oTnSBHVYhKVTaUn8y3R2TPkfHK/9A0KlzfltbR91Pgyv+vppNkLSPH9aFp2ejiranr3fzo1pJT
9VYFOeayMqgeZjnJEh4irkcNULhG9qdVGLywYhCcc2PaiSumMDgxzUCGS2XYh2XXSqmq66Gb/fFa
HRJtuoLTiRGkkDV1mAXKVyW5PeFcl7a8FZfbll8Hm+20MSIA6hLqPeUiAvVh4VRmjrl7W7eWpYpv
52tXXc9x3Ypgg4ajotHhouhwCDWK558RLkTvRxfWYsTzGfO9wq7Od9aX/gebnldQKfndzAVzwum2
z19RTHxGC3XjYYD5ZX7a+OKXblNzmr0MA4dQkfRhPqL/Imis+opoxpRIwpeHl17/QN1Ngm051CRO
vi3dnO9UJbzTO4NdUEktRyVPAWfdPfj59M41sEOvXEsotTPVWdO5hku6mC1ER+xhllJnJOqCHCW7
776s03CLAtyLB7OZVDU9zVxyCDSeSYpTUNPrMSpf3xumGWTju/NZ9Ie4PKOyCsvpjjf4lmGoAoQC
3UaEG8nfagggAisdJV5tOKBbnj6VMTmAPPmXRKLUjKtbd3KEeX2QXZKCbiaTN3F4kJm8gLvPQDSt
zvY4ex4hNI2mdQsLH/i5UzYd9yvbwzylaQ3piTTnWyzOEBgytpfqDrZ8E0azGxiGR8/n6JBiHrRh
sq65+xv2/nZYEJDo7TR6ivDO3GZrEHXFXoklJj+tbGX3bW8zRV78UfS8lM7o+4QM1eT3M0MCqGY1
Ozu0+iYuOW4GBCJNdzy0FrfkYAhnh6O3IpDZ6rdG5NA4wdhzyQAwK3ACtt5Y4KXT84uKPJaO/gdi
x5Ls0+Jt34aGeBCkAXCii1bY01eaQkrQqfuEpMaEkd2PQJDDQ7rX4P71ICMhLbipbiKxKjI0g8hq
yKHcD+57DHeSlNBETUhZF1OXwz4UZWRhxtBKyFmSIiRK7yDnleGvKZkMR64+hW0m/wBbA/wagSkA
JRshhdeDdmMM/Zd+zhVQFyH54qkhslnaVdVBR2fq9Ad6YSJEaQvielxjgJtpPyXyogtHt4lGAz+W
k8FKqGMwDkIzVX6T+fofYtq4csoSq5sqq3yvs8lxN9IfQkFrX/e+HfDVIyYHH5yV/GnMywvRZIpA
DFEBfTa52iExg05N4XzfT2vwE5r86IJ9X9cmV1+UjCBn6ugjDJcj49j5YI8WXZTqk/kMZrz4DMN0
LP4b1n8KfH4uCQkn3A8o7z/B7LEw94tM3Exl+SvTBdqu1K7Oo5mM5/T4HaKW5Qp3Yh0G2A/Wukwb
6qSPXckCdzkd+eBW4/FyyEmkKVcf1SzYpTsIUiVLwknNOkA5ZtB2kufpaz54Fa4MU9Kno5XOAq6L
+lju/sHGOp9luOSmDcjGALtlN/+SCrCwLMrEyk3cLTXYJZA9Es8RQliij0v8KAoNf5fCoQofgtTt
XQasiVMGRyBtFZGGuaj+pSz1JjUzQ9EowmBjd1nGCncF+jK3UdcTjJdsbGpKBQY/oB/09Zr8e4Fk
OQaZFbs8U5F0kpfKD4+uH2EGXsrqhsJq5K8nOD5nOcQafLK31h8HmrwcfkKuZCKqSEYuvbVMm2QK
W7mjs+TZTj1NT20UlMBu31KoQcqBJPJ0qm10AHZHLaK2n50fgIL+fBdqVKksfMvjBBZyGhp8Kr+w
ZdFbj+9VN4q3dTjLA/PPUfTZn3eABW0hDfkReEuXxDWiziFOngikJgMtuPMCzP45NO2Tj8wribmf
933l3EV61qBHyigVwFecLICDyxukeX6EN3Bdqt+XdSebbq/s4td/nj3wYiwwHWk5ExKNMGQrGN+T
mLqF8ivIBVyTuqfDsFERAwdsBAl7zUgDzKuxGQKbAeE/YA6MiZXIo8kwl9rPUn9TtNdX6Ikj4TZ3
ubNMGO97KdVkpLOlNJU6oQWHZRC2VKABoWFqj8aLrV0qAOhShRJy6FmS7OqQQYSZGFJnxAeK88R7
zns+eo4YP7nUwlv7aM21ohNjZMqMbaZbhccyvOtCp/RBIoS5t+4+XymOJny0PvPmErJp7l75Szg4
qNLiIaMFHFDMfUj2XqGwB8uExzv+XYBaCAbzPd1Lgg4mUeRSYeEZNv5J2B1pbhd8V8oJ+kh7bT7F
9LwllEpRvfFOxv8QNi1kAN9fF5gqu/9I7gE1HGAb9QtM/qZB0w0n7zLDwLs32c+1gDz1/qCL8w7b
x6r0b1u1toJdm1S3Wma3ybm1gRqoaJN+Ll24Z5wsysytPKcjl4iR6VQe8DCAfJ1iujdY4ix3Oz0R
1vnjxunQIesnfa2cc55VSc6dvahdPJnoWgUVuvIczX5u7ntp9ICMHsngs2sjt1MHnyQHk96UMajQ
VSI/J5ueF3D/S9twSXjqlS8321UW+NH2X1bUezDh8W0P7O4LxsFzuQWheCQdXqNY1M/4Drsbq8vQ
Tr8Sas3y0NXF8zUZkbsRDGOTT1aVle/2oKNMvAd4oeBVSUmEvp4VhimY7jHZk6TjIzocc2DgeE83
f+2DE2b8F5mc5c1u+uJcrvk3rN2hPxs2156i7vPoaOIcmTm43iZHMk8SBBwvSeNoZ1lEs+V0HYhq
5mJuVcvhqJWoLLOTIbfGSjq9+tGLGZjsVQYLA/+TVfTkWqsOoaHbPFaAZGCn5E4DSoKngwFbZacr
ZmICIKRgai/jXKAcf40vcLbrPbvtgYWR4bmT39l1dGjJfh4fKR/64WqApgB/3VP72DVkWWnry7cS
N+h32okCpt7ed5gvZ9PS0TZrp19BH0Mr5/r9yn5fX0qoSWiA/13pCXt3GRLZNANnUcyLEO0BCQ1Q
/ptHQZRBZpHD8Y8rpj+Wp85X5ay9rZ2SonfLVzeAPr9nUgM0ror6+7Q6LV/j019ZRo9/DJVbsdhr
gjbAwK1Tfl3LmLqhP1KE+vh2xjUB41wTluxZ0DjxuLXZnIEwWbhqszkmvuqujtxn0ocy/QeHKZA/
TOdBPcwF2DLHgLOwt7NEYDQhhZD03Sw6NRywDyk4BYXYA5WbdB38aZER8CWKV08B/bs+cKVr0TTi
ulnsdtieD82e6ZNvHC1Enw1t7/4x5dD6Tjp+BnhnfGRhOmTPJi6J3hU/ZgVKYSR4Ga5Zj6zRo+mk
guEHHZoz8olRDh+XagBye+SV1Hs/eSnSmdaCA5KttkA9LNkXshDUT6mjppxDhkbPE5P9oCbGQcQs
I4iorfpTL+uGsHjX38NerGGmBsN0pqA8FohEZ5KXzSwkG6KGeNr5LnHVZgzwRvHs/wKt+rLcif/o
BvBmZIe3EWfQDhpqEvtVAEHmd9Vb4X6/tCGLxPemtCUgZ0IkRgyQcikaVpcXY/4RbhW+m6QgMAeY
g8MmlNRS/ZIQIgnyc1ArbtDM0fP7h/juSRBEg2MiZW0dzD35Nwv27IxPhRbAb7h9fjGvHmdLzUHr
Q3Cmf87B8CmL3QLEoVQqCwsPIdp6f2A0JeoRSK1PYkbSajyZk2g5OW1h0SM97Yezh7yOtK0KKcnK
pHcTLgy6bhh+Ao+SDJdTO49VDfRLvU1AybAwZ12lbK3A5ENGhbUcW8OWrEoihj7u2e2G9SUWaxGd
BnJUbtV5mVOIRA9Xr9aMwc6r1H6U9sXy9xgkmxyFkfQSHDsnhiqDe0XR4mr8Ck7604ZiKBV5glfR
B7kEMZnQR3IiaFbuIUUZoJah0bqEk9/GlaOs6aRA19unALIgsO6+B7HIHzvb1yor7FxT0TJYwt4E
U+e3dxYTic23+MS5yJoK1vET48DnLL/MG7rGG8E87mC1nbh2fAyBR9lIvNM9/JQ7K1YC3AiIXJjH
fTnqnkgoV6381sv8VPX0Joko+X+BdMA9CN8Vxj5+J+Nqz6+IbGVNPIjefn7dbAmZT48pVvVMVUPQ
1j8RpqcKaeeBZVLtFTpfKN4qPZWTWm6ikXkwZB3T3TcPaFSTmOXhFefg4a9ItkGKxtraGVHy+7qB
nyW6dhp0Hf1iW74bAhT6817h0iYK8vowNIgwA9goBOdkOgwzZMO0lfg3kJgaiaYle3CE2lRqP7ei
ZTvXQVH38Yh1D++cSSI8D1LHgkifCkK6Kkg38XlxpmeWjQzyhJ7mNmnPx+XrWitMjUfLO4x+17eV
YX7EcsI1yP4EoqFJ6rIrEilvtMrpSq/ZUOy1UD2mxESdyFAwpodH8+RCKQ7l2k1olYEtNfuHp/fC
p4N9kjQJtPWPbHeeRHVm0wHyLK2y8rXvtPU6zoLbgAUYsVBKx/hYMP2PwwrHL1Qqy+NoPJNxp0ay
2yQ13Y5QnPEF+AHGMwY336bUktpCgqXiZqWUwZJFn4gLtBqS+LFhBYjTgxaeBb4sFcOa6qyL4jTx
103uRAiFLBZdK5FSQjdbTRfDMxRDU50qIsQYJ/jblbTA6eyid19f6j73jluE3zbxH9b6L+gFfPNc
5wnsHldP/GjBVVIEAK4EhbLeB3MalKu43pG/Dik/9dzoBPMdutntDft3+W5NpdKUeIW/VrvBK78Z
/T1/1KKy5KuxV6rzrQfcdUNLEx70SiDERKDFaCvY6JjVEQsU+8WM9WgvWMB1EIQ27u9ye2/MkZkG
QOHyUhGu0jpXGr9ajQNdCGUBgKLwBOFUPMUAWlnA1/uKWdQYmJ67ZXAg2fBiXrcTOJIVTiOWD3OX
ppzvLt2DDy/7OOnwqMGWgE5CMBBT9D8wDfGIlBl5bkspp5vE1+tMdJxqsP3nPpLW69qx+t0QNYcx
suk8Qc+d5E5qMiDKzbTJA9TeM+y8bKSXzXrmJ7qVjOdIe6/HCXW/PM0f1DjnK5mj94O/RKPctG8l
YMXNxmTxLvXmHZvu7LO8ZRj/+HcRyw4F//4WU04mdbcNuBqzsrGOsT+w2wGEjMgmFI2l3oASMdjp
7W9QdzVxF+WDfyAYjBCUMam11GjC/RZlmtaPpIibgiYaA4C5aO3okkAtJNs8c0OkdJM32FjFS+Hc
06fFLio8ZrSObgJyqPQO+OMt76NVSAOuwnc8ybcfENeNWT2CIhUN19rUDLoa0I/QXhoz1Ek5pSCK
BGdK2OJPo8oqPgE2+GNyBxVYvkL+IfxotX4LJNoGY/+Y8ffiACDZEK0gMEyofXy60lKOlw0ND0b2
rHYOLelLSE7ThKUBdoz7dR+Ksc/+apRp7q6xcnuq01CwplevcuTxmbH4vYG+k7ycWE0jV2cLklUa
vRe4bd/KsPcHtfFtG9jcCLKfRTOPwhqx3KAmizHDmQvqr9+Gr7jf7Y08lJcM659hm8g2u2bnos/b
X7Zhl1OA+DhAg4zfZTSI0y9IpGSpLHiV9r/EdiwvpXEaQcpb6mlehApQrIUKD0GNEFjR8LJGfPqS
251GA4FQOLLQfLw3QQlzhlHumEIofJgcEBLfFdc0l4jI2ZU2XJIZniXgd0UE/0MX602on8CPCvpv
3duV/QYS+AoLsSlM++8Q4GHSe7j4WE+E6OYvvRWt8iVh09Xr1CdjOqj5XRiidrvwJ5Um6MepJQw/
fnE7Bz3t20ZU4w+h5yKrgpVHqcUIjHtoZO1xCo7AfrWxpolk3tU/KBApesOmPxomKqECfaTTOWWQ
+fbu6vtg/SAp8qYeKWX8bKDyV/BpA1d4KD6iuL0UJodFF8lB6QD8J/7WaWN/aTb636GqXQuYJaDp
+4aonTeXJbuHVQUiU0RO/Jx4q5LCopFG8Mkz8tf9i7OS2L6R7ihAvTBoioxJiJjHKm8S7L29Giel
8uOCwfQRxINNUUnkNu0pD7q0It0kUAcl+RdcLaCpbnR6fzzNICEwkX6+nsbord7QWbUOvUiWXoYN
M0KJQ6LvFUktdCJ0tJjulA0G1evPxvE967PsNrImB3nazjJjZvkmQgJoTWC3dNJjv6NLx+Hpyc9T
D8SFuh68UXPa2ln6kR/BNHtz+MPcTOzqAUgnArWS0y62DbpA5ynq8gE3tLnaose8QFPr6HCD95qr
g4L3OLiT4VQ590SqaTwFnSICVHD3LbgRZmnV5kNw/P4EpOm8u9ghihj6NmGaSnm5ZmeVOUodnzN0
RbMlnEXkcCaIC9wqtl3hQDfdV4S9T22470grTUGg60dt2pD/G+uRZ9gVPDaMApzplQFGFWeJD1Xv
N+kZRcsVe75tbw1oR5/vUOKS4UdYkEr3PE7KHr5GZtA8/y6ErtxLHcbc1LtcbqdRq4sE0bzpFvC3
LFZNcNG5MKSsVwvPRKGknPuJ0DKo/n9mEk4o557J4Dib+OAUY4l0TAWn5AIduSaQKp9l4cDSWlLh
+4Xd1r1IFYq0K/ziwtSign8Pxm4XpK9eB42qPyNH7cucH3BjIcAUiqfapK9oIXsBnU/1KfkkxJxp
m+iLvl1IDgCRHhSy0QyhBqZTF95lox2ocNtUE9vIrb4X3a6rbGZqB0vssUaoO5YPY34/p1lHGM3S
hYB930CIzmfXxyasDRvely8OJ28Vm7iMZWyo2P15IIOgVTeM11xThy06R8LVZVOoEfmDc1JeDfer
xLFkAmdwpSuAxOI0s4L6PphkajEVONGe1J7xExElkao+cCg2QGPgfnGPYRkEQwdFHQLcNiH76vTp
hsrieQTgP56CDqCodkC5dLycyd/2DUHN4evvOk4fr3DjB4OmvzaLo51IaWt7onES3a1+3LgIgBN0
3MBrljz3E6jYiNn+j2ONu4JR8G9kghOePEjRA9hWjZOzN63WmMabMVFiFVoqF7zJHmvTw4PE/n1m
yWFrG+3grLAQX+A4AqEV5VenIJGNaiEus9SPvto4E57E8bmUWsP2KDe1Xdwie0oIqJ3r0J5Ewq97
IIKVQ9S2qEMOlvwAFulxcxP/p9bAluV81WhqQe3bLRQPUJUEWXYH77/8n2EarKOJTVepJkC2PACO
KN4a1ONGKh5lOCsIfWev6p8BpHlsA/bYRwS9xBdg0zOJzvohmInOqgW6+UoI5N98K4OdXOV2Dtr2
mTxa9guN/1ugNLUSNTDoq23DfCt+l6aF7BUHydBk0YECs5WHREYik1N4Dw8DdeXmpF1cL3OlPt9h
h5ytq7ToPObaDzLBr5uUVo5s5JdyWDES7odFdVWuk+hkF5dxv2x4JjzfsWfF0AlR/TDeh95eQUr5
Gz+AYoMvMbzHRbro7EGA7Nh9iwj9lHaCFU0igSO0sSG5p9PjauV8rshG2Jl1/xPE/hMKA3b6e5uM
rRKxuUH99rlZxlpWPPm1quERr9XbG0lZiKov01UULrrzU1F5VPpj6kPcxzJIQfbdlhJ8HbnCmWEc
Ex2x51jtWj0UwmKLnPG2/+EFM+CFMcJ3toc5lRQNtVC+XnQXe9uSaamqmF95kMsu2aEneBXVaG6q
r8dh3eqxBVF7lhAlrZGH1maQTDw3WPtNewNL08DrYSbT/BTWYQi7JBHb+QL/a47UpAmygimEs8gO
Ag4J/Ly9ejUwFslWRDZ2ZuK7o29h4HMbuWoOnyGVmCqqXPiyPmmIDezCtJXLGdJ8sKIjOjV2D7a4
opZ5fPbINZmY+wbKJeHyUniPEQPO3hRQXHdJsOqbwuOouZcLPxvboFiTUG7dd45ctfCIeOqDczdO
su025wvpireSKWZdRVwC/H+RuGHGH1O+BvqglRjJWCAFeVzxt2FLnvm9z4NNdB48xZafvAdCyrcm
Rnrw9qBraTFSoBQ1D2jxqwWlWe444RnpGOoHzTA4gy5I29kxZhKstudkQeA6yOyLAal/HB1xrZ3P
k20vrR+rOErKBN3vwzcmv5ydN+4Z5lpK8W5nFjfrSgEFNW8wI0TIutk+TUSbJorYDPpHn2jTF5z4
Gtnp3jchiwkCy6onWTQXhIUPk4GSzgQe7hpHHafAygLL43t6v8ZDr4S4vjoHy3mfkwcr7flxg3Ig
DhTxkSKYdmApyXwtalWF8tHCz9b+cPu4f14ChTrbacneURWz/fNsYIQn9gq4AXrYTPNfuvUnVbpS
kq3/zdDcI4ujNcUDc5gqw4oeMg2N0two899qjWvo4WHLq3Bg9Jl7zWuq6VXrajC47VrAKNMq0XhH
vHxV4tt5V603uRkMIu6TwuYR5mtyYLANOxq8f0kZ6zZ5S/SwqWx6oCGDBDfy3XiDaYs4sHI2VU0R
zCQvXxJU1gyA5WGIEJvuxP84Kt0YxXFoiAnsIVtYowLegmWn1O68C7RW5fPpoZAJ9o8DDgsjHvHp
0E4kqjzWhrvGPTsjlzAbOmR5GSr8Td3ek+upxzjWV4fJc1Ss3JmSXtPcfkPdVFz5e8fB6Lcbn7iP
dJ0UgbF1lRfip1yvpdY9YCtB5MpCVbSDHc1exYJag0XEmklTiNLqMiHNAxqosETx01SR2Damfyey
NMfC6qa00bd3HCqTvqywPXIUiWMUrUS9PQZjL2KHo0SFA/MAI6eM072Ibl5DI6Um9o1db91eDBED
yUqO9vN03H05Bny+5kcPG748XSEaa+QTvhzCMi3XxQyuARG2Dl3gTYG1ZcvAURmcGVYXjA1/NVNu
vX0vsnln69Ot0bQ4unNs0dwhDjIaNWNevJgHmzdQeNJlC2tCVhAyeF+luOmY9TP9GZfRQreM+TkC
0mIcN5Iq4vlrhjhvh6O+sZ6hcmytWzT85VAhkYHkk1Cjx66sYS27bguBSz8/ewY8GIQydD8ujP32
LcU4lQIOZXrf+Y58Kv/EkIgQM5onqhB1DTy112T6uTD4PKNKvCCVvf7BozjNXpoRLWSM3iJmWjqH
5+BiNN3VPkIkd2whvJh0JoMbsRxMXkVlctUqt5AxaMnakrv6hHpGY6VeUcKRVHj2QUB9cm1VxfJW
TE4ddmo3AT/BKhXNinOHs7lHPkQ4MdiE380piValUFVwO35pRaJbI+UFiK2AfrcZSF714cgNXDQv
WZNqghasdAvalFT5Mw6b7v8s2UbLjRQ3WwYsIHzpOBl5xLh/DEW2JRpsg70MHDhC8Pq67+d+GEDv
SQJDC06bpxQi57hdnwR+6FLF67gfg952g6aXTm0w8kiR95dFAwrBhLf6ZVqIR/45Skx6SaTdU8s9
VE9MpLzb5F0M2aq8J/yFiN3Cj4nTNm9wpP7+ye2wAs4fMzuCqst+zby27W8hXWSjEiKaCGBBvJTV
gUD4JB0Vk8Jna89pB9B2q3JqI2xV2SpH21cBpzYbXm/qSZ2E36jy+79YsiHP2ze476Lyq9DspuEc
i5g54M44/Z1DlL4ffFYaoPDzylVERPKtJS6PJB5cU+2B68UWm8i8sH18LSM79n1HE+cnU+t/qdiF
NgicpFlQC8wY2CqI7V9jzWsaqSjU1zbqBuNZMo+dqcHjrYHXpVjpjyXzJf529PExz0XKRpx+v3mK
U5YBGXkUCEn+yFcCsMJ9+uB9I9ve5xszA/a8HFkxmIUqYRTjG8zMvxM72uqFH2mE/3OR7PfFCu3O
8FIwg/kXGx2VpkJfoDSs/ElZlvsMKAPGyCJZt3kO9y8fBBtdNltpFnoo071xBjHs9YyKwcCYK+lj
BdkQMKYG4OrmBhJAxglWgklDmyEwQg6C0tK6f4xXrQ0dCp+AFFEvJEQHzmfcTrhKkoKpxc3zkTZx
KDE6kbkj3pBBluWURFckAfU73bo7F66uESJqLocQC1/zXfv1RFnJ/Gj0ZK+XbjuTXIoqVVxkylLM
79TDXitipageL5Zt5Br0MP5A+0NzAAJgPxQ1Hq9itor4wAkGQpsUMgs9+3UV24YfoL8mo9e9QdQ7
1Mv1Avix5OoogjuuOqnPF1VieLJ8glK9UfgMYFGAXq7EUjSidO3NxUDROfyvcXmJGtz3XjiMic4u
3a95H+E+QE47dCpnamEbn7hGB0S8EshZRC3GiuN6fztnDUJfGbpa+TcuYBpPWmEjF8ddKpFMJEgd
UXjt+P8hzPfjo6SrsYTamjKxYqtU6Yd8syekxGcnc3YNJY6nZp65lc48hU2YvilgB9Qh6LKlwEqg
kxbcgwS5to7aYYR0crCmcK5v4KdAkpn1ecmW/OpB+IsVr9cthogpcOT3P/jgp3a2705Mhny3HrGr
eiE1u8dHmfyztomWeUNerUttYkD743Mz/ctGfrKOL0cc/9WUXXo1zQ7Cwc/KcTCifdstePEC3rmF
dI7LsX1uAsx0jT0bnXZixURc+Ab5H3BnUqhzv+j8YHY9DpZw6eahBSjxsUrxygfbQ81se72l0T4j
SHI1iEt29iQZ7vTrLtNvjmr4YhtobHXyKw4qci+bn5YOAgXRHC7nRQea1GNM2uxDrWV/E5iYpqDj
Cl5n7+lXK2/pSL6LfVDL+vd4HVzeIrt7kVWksqoJZYJuR97V43oRTRGqucB0MCWThBoTav65YtL+
Vvz9/U739SXvZmkU6pZ/loCwOK/bZIDcjvUqxErkN9jC17COg7Ol1Svi684UBCz+9JOl0EcbRde3
Ji6vJXcgeKdM9W5WYkHKg1tn097NDirggwOYaJYeM7fyiVuqHhB7gA2JvtDI0GJzRgKGYeEW8wdU
wrhV6c+2PUfTsw7A1uu9QhAizSrc+9ODWeaeH//VJ1+29uxQP9jsXQrOHd5EyLp3S/qQjzvoHhuC
JJd29UOdsfmJ1r3/j7uuxLicd08jwofkKLVsEbE8P8mNdgXdDHbLEM9hXh6DPp28yncZRz6s45QP
ZBcLzf6rzZa/ZD3bm9OwLsWtR5u2aiMu5cfDGj1RJ2ngvrYPN2rYgnDr2isrIvyDEPLH5AQqoP3v
TzoqaOLu7uBeKDdCrb+Lh+xJ8ntOgfTZKgWjzbR25ql+mPnjcWvkdr3TCsqOwGnGAjzQxPhTU8yH
O5mR6fDKkvzfBLjsXtZ5lMW7VnQ0EREwMYJhgNIhuFgNInBfCkhP7O6BgeYBZJhZqC+cnRBYqRhq
yWi8TXsPSrnHqA1W5JbUnViGSRYxN4nODGVvxR5ptYWGEUV2MiEKqfMNXDIrtS9ywDz+L9JviojX
36h7a0llCK/6+v2xiyt8xpUJT/BLm27Gzdi/MLZpTBk6w6PU9J9qfw2O6Q03pdNvEmYczw+64DHp
k+PnQBuD+BrfFVmpEBszvzQjUrWKjXaxGvcqZ4nMOrk8xuGPBFamH9n87XFvC5G8Jv0Jhoflqi+y
XpyqF6YGKH6wRsFUyGTbR7f2+baFcYYLCMT2fYrpSkP23lgValKOvxxexLyxXAC5LH/+h2iWg5TP
preK4asUQe68dVT8vcY2ZCbjHYb02lXUFTyXSCRkTcPRZ9nSkHFcM7cVxDJn/kHcIUJB5+BbG80f
CFdiSrWRyvxTYZv2r1zE1wf5ss+R6sWmFYqszThtifM2eI02Uwp405wvjtl0r3P7q8yVWVcEpAPF
jF61ORyuVyAum2LdSGflhnmXzarvVoTuHPtjxSTirR/NaQWzHAVFi6wndnFdQmyEHFgCPzqoLLk8
fToTYnAp8sdKULv6IXLe3knfi2qVdVB1scoi9j3il048mB/6bQ5hEJqn4Az6OEoznczseBJYwd81
1EgTel2SSESirnwxhp5uTaHhHLxNx8tLNhM1+ejurW/AxtzXeIcANQc1tZqVA4S2qZtZ163/cxhf
mJ7wD1kjfhRU31hTHPatmrWALSCOLwh/dgPqBRi7gAK4MpdbgsT0aqdqSSgqAbETEdrJJjTv0z9D
HMEw0RqEnuh42ZoACRM0rZ6gy7wkbOSIcnPXgR+2FvDxmaHmZLUljGHAacYulX1KVKngiMHFY0RT
Sa+C7T89BGWv4zim8bEehArHDubBfcndlkd2yx7LbaYqQRDRDZ2vMCcVNkHJL+TfFRmTLZQFVNRS
ZxpHHxf/1oCi7XinBVE1PT2nRBbkiaUGdUrucT8HTL7NfNBNwumem0k9mU9sbQjTghCc2y/wAwb/
fgl8EIJr1VfIMTEFSg3uHsoKztxenf0RELrGRJQrdVpljk/AMGpsc9dogsvDJIhBF3hy3dLN+Z9e
NTILYbxRhWGuM29Qz39MbOnOIoCbSQ42rrtNPaGv6wvWEBvHrj8c24tAFLA7/Scc61bOBpiLCWGR
W1MdARtuhQf5OU+qVx0N3F6j0GjjH7PLzkoIc1aupS898qFq4f9pY92tS1q6YOKDLaQkwViXwaXZ
z86lj7ojcaPRZhFXUoVPiP2n56KyXLqH9MsatlBAen6ZxSgfp/JYcVSBiDiZCRWs65EC7kTC3eJj
4JxaOrLfVJfa45UT1lOQetcF953o4GafplfRmXCbc/qXXMLpYmtodDtSdmk0eQOjqb8QvkAG0xjD
WmgZYVP32RvzmC93o9mTuhWthu1f6J2DLo4KJUx5HNeDRQQgJ82vs8J6pYUjlAau5xInpHlsAedx
QUPdlFY/xnbjItuj6xkgXZ2rtS8WjHRM9zt24WqVXFZNgJNEdAnXZbLvMfkhKQ4lpjlo13UIPQUw
wg4D4mWZL0C0ouhKXxQedJdGPxsLIbiG9zYaYq15chrpBZmJqadxNM5JGw7FLP+pDz8O9GY/1jIg
1MCuM4Tbch+BRfiQx9BNANVk+YhUQV/e/JbJQC1RQXtVyEDcGbDnwlz2J5nGtaQ8vychp6R/Gf5S
vvkrKTUfygCC1KGZ5BPG4kodih6X+fOZw2l7L4pGIBQLFttZRA4+050Ff17cxB5My6R2S+K98P1T
xgX7MVyM5SDeT+pPjShOIq+iYfbgyjfqX80Z0Z//8GW8D4vHNSl0pIH80OOKKfJNJguregIe9OJw
6VBJfW1cR5Hi5y9Zyb2PM7LVdCW3cfn6gHk4xDFBRIZzCPfHAhJvwk42Z10/KNOXE9JG2vozXDiZ
xk38mflxyclLkwNwOxopWKiAjJFP0tOMrwqCQRjUbFNTNmiv73lLhf3Wyglxu15tH7ny4Tfg2qIu
PvRtwcTFPDlna8owfiKt43/XVeQdyeJ3FVv6e6oDpvXc72EFRL7clWKgLsbDqo8wqvfBKPIX6utR
72un6wCzaNGnWyk4IX/ZFbKlyV7c9KuvjBqVfIZLbLRhdAqDTM4VrT6c6/XkqMyxLbLLDCNtUCfP
xVdLHXlgJMN9z+yqMUVmNRUuYLG5vMx42MZdzNCZ1GewBpHtXjsojxaUPkeczHqj5sgrj2RjCuEr
JjwHwIz3b80eyjn9MB9Odmt3zw3L7vNdkfV5TGGaXwWR7NJ2IxavqqdueAaLC6DGc4wWuXvacByh
x2nLsMsT+eL622jPgxqS/pA5G4Vjxd21Uz9sjBLR9qkEuof0oE4PgHfP/kq7Ktw3CdMkXRMDaNLe
bTcmXiBNWqbabd0vvIN6pMv5YqWaM8w82H9bLz0vX8Qdlkr4DvqyTl4aMvKajgVf6wY1CJ8yBEDh
YMo91QvHz980lSYWUdCEqmT0xB1w49EsYlZ9RMudH2yc6DNijjs4KTtaFMYxtvbdcSRNOLawFVdr
gJUCJ1IcUztK56vcc+pW5DKL2DqL73B4MCnoKVzAQsW2+APo8wHV7NL55DG4BQU++4hLjzQM5Lmg
T221KFc3N9/LS0ld/596AD8naMNDDUH5dSXANBt12QRKLJzTy6I62oiwWS1OLJYnK9KfwI0nlxAx
2l5mdXwC+RnAe1o66ZbSzAHM6RlxJ/w5WsCzlQIbdxs+tPEBGEupIfwEh061+aulW+X7jCXRniPc
uaMtkXs1MY4IRP5cwXLhKv9Vcd5fMSOyRlghxXONx6YB7aHd2a0n1bfMBccX7rnbSmxaIZhXwxXb
EKl1gWig+ddXmelDhuWoaEZGs43y0OVt4wpZrnvlDIdH80vX5e5IHyJ+YKd2ka6Pc5Hs9CeWlYQu
z2Zr/2tFWAv+7WFWYa0plGGg5WWH0DsktSIfqSq0YxGKzzfe0++ila0aOn0EB1nySEt66IQ5M8UD
moylQZduWwdOlfQJgIiikWOl2q6PvMOdoVCHMuOn+qhO3BANeJc4oc0tpE5VQLmbbeyj1jZA4X5e
er/z/hwMP9tVWWl7Hebe3NCLLMScfO6DZ4myiUnSkushCZ9lL72Q7lgC3U6ur4AWTnp+dJJelQWn
TMeEs0uXIbXmqHgj6BhKzawjJ2iR7sXVdgBR31SOVsKMr4t39tAHarS/EiGEWeU7TYVKyU/pefdu
bcvyaBcGsLS+rGiFmQF9GnsRIjPGQoqkhze7Pq+AgPSHH3IMuRJhZ/yyva9iq21IUNkIM7Dw9VO7
9JY9c6mSwzYs+UpYoI98ylaGO3kvHrc98V01aiogfNYj2zAYzZmkF9D1nToLuST1grdIWAoxTxvS
2NjRP/oUXsM63Iu61I+l0sOyqDxfS66PzyrIuVN66Y8De3LfOcUAQY1nW6GtxSQswe19SvkPxWlj
m9uQpEcEXwUvUZElUFJsfK4Oo+j04qYjILeKuyFn/HQvLTazUbXpxFX+QA5k/s9nYhiZA2pSxUgw
m6pFvigd+x2es0InNQ2lcK6Sq2RICQQUxbt0tAvdCDywdsMZouiUkkn5oZAuD3XutfxKf9Es6YZm
0KX6zfVeHq+aindnDLAoUEuco1+aa3qEoRr0AMIk1JTuwVbuIBc5dIcZM+fEgMHWMtyir1E3Efc6
gSVZbzax/bfqEOslFq5wV3UdzmGtY+GBZDQx0dpman2vjuLb6SiYF7kc0OzLNyQd27QPJfdIIcnR
7SY5XUR9Pqh6CBZAc2ZZQjWDYHriRyewcS080fVazY6sLM0PqX05GuFi81R69fmgaFHEGngnKYZe
YavZ+ybVVSY25bJinBYr50IsJjxhpL8i5GaBrgBpTc+2PbNicubSVznJJ9r5dB6RMNL7Brx9LZUg
WrVhzdL5/rz8VKbC4NQycxTP8gaU5prIwkXJnoVjRxs+5NhWoVsPGHf+UQLFtDSz8UEWly6ydX8M
p6E6lZPwICCQBtYy/38ur2BSZLD98PrJXdhB67bsfDCr0JCdFm/g/oDeouJaAdY5rWUcCH8MiFmM
+CmBDTIs+MWd+wMrrgGj2NSZj2N2X2Y2dItzsF1crzvQt+dMGs00P4AYAy5QWIsKAwye1y5wDrVD
EsVW9CCdnGTOHjGaRfvXqgcf63VY2RtlQ9bvMuvAzmi1Du2hemu14/febHJaNjvrdAg/9gT5LmVV
MVIkmuCND6F8cPsCI0jiumNOorR40nsVWNdpf7zBj0ZvzKq1EjIYGbnpN03V5+C9Zu2j0nihCSB2
/Vx8Q36532LjC+9UiHcPMtzeHW7YElFWOn4VrZyuX404t394rRdxKuwC3JUgZp2PL6pqRBpgDCuV
JUFuypZ9TtnbRNAePEwtQxsDl39LqYfm79m4Q2dDR92/PLHa6Y9BeUVH4xjhGkIqu/tAx86JPix8
x+YQ0Pa5nc+woNVI+jH8KddO00wz2lR0nz/U2/w3SrbPWwzciHNoMdxZMHu7xs/f0K2rwyHtfyGQ
BYh/hl438VU9jrHS+/HbWursuAccRxGFYogrCeduhMJY+RyV/YOjeZ56lQm1uYeBvpaDZo98fWmW
tPf67Nn0H2nq6oUckWgAQtmk9ZSjTWGtubTNkduGWIPN8Jl9lRvAkpWxk4g+gjtJDddz2gk8vo6s
1bgWX7mpRdGYUWt+sm9+9JRiRQaGwQ4w/DMPK2TqvaHM2VOqX/M4bvgzQa5Sj0Z6fXTMutYVUVxH
8Bvd0MQugFIv3+jszGolXgUzN6jPaL0OGF6lrQShhM0S4qcKLKZTW1zzDYwaB7kGAXpPEAUA21wx
s622F5EdXZYPnwrQWKk75N89XQVDWsVygKXfnl09DOOfIWmIMzH0BFDNB6WwxrjN73hW210id2Wr
sdvF5rzjUtc1l3NvICTOeUv8OEU8IDC5W8/yuHPJQ9+VOl4o8Lite0N7/n6hPUu8KG8aueWSgq7Y
lDekbsC9WsqUanoQ43row6GFkkBR3K4FxrkZ5hcnpBCgtlxPhOGqqRVLPFGpo1Dlvyvw5SKk4xW8
3tuiR1o4rHjvZC8a2FbnG+glpThor4gMThw9Shl30n5dQ+9KZ7waD0CZEoJYuKhpYz5ge1hs993c
patPcjthpVz8UfgjINx37JLTzyrNUemthjalTAWQcBhiLvG4Neiy66P2dLCExCXR9689uvBC1rsr
Zz/epILJ0CAbNRqC0vAfTxS7pai0zmZnSt6IV8R7zR7ujb8qKugchMyYmmf+YHR30vE3H9XG7952
BCm8bXdCeeY/IJMPeMOXGx8mmQElLYZsPssSDM30jCQHohk/2DUtBQ5243WKywZzWqmVcs7nwHEq
e36jypiSbvCo4Lv3wIoT6W8Vz1dqs3tDuEOQcxfDexWNKGZCRzrEbpThCkvknMCjENLY6pupsAO1
QkCbC2yzwEFVx0jMqJGtpu0UBqI8bvdj4FhcMsNVbql2BbK5kUM8gVYrkhlwoMMTf6na4D7Yg6uO
816nN92OlomfBCJwEGx6qsHVwxEUOnfDjTTCrDBk0Kqhp9FSfJxWwFLoUeMGcQQWhoqejxcWUEXy
fmznK2em0u4YsofWNXMLt7RZdSmoxqYevQEBLHycpi6ePFd2jw2E8QNm/8GosEaQMP6HSdtdvotc
/mDleXmkSredCMr7ypo9DJ3CuiRkhApeMaOM8j/pBLXgOqqCneK6AtMjpHsEox5kXjjKz0xIyw5a
ufSkUi/xmwvJ/VjDbfBKOF6BUZU4xVCgXHsnmHKtEPYHtB5vFWZwGmSlOWHTgiX0cqAQYwyxFGdX
bQfKnSAlnbv3+O0J8zN5lgy5TuMwDgNxDr5UODg/nWCEp8cM1v4vUt/E1A2YxrQLmfzSwvHxn2lp
tle2lfxMM1zXgiAVUukECrfXbG4W/f1DJ4KRR7llDYNi8bL46B/GawpQ8HFWI1fonZy8X4Q9QJK9
0G6DjP3xy6MxY1Bq44gP1j7bZti0Z7Q1TJPKk+XpzTqpYXZcEq8kNktERdT6benzi4sb6y2+mfIJ
SMeAzxrrRMlWnZFnOm/rL4xaFxlW0PALs17UER+AcyxyjZFswPmQEubTbxbNka0q16FhozYdNC6l
eQFWesoyunZ+3GKVIS6v0jXP75OBewLS/SXyUOjn1PnC1rK0aJQTW9Mqfkr+xtDR4Ehdas70xENp
KuZQkR0lPJHmcwvqL3A8/veTLENV2wla8+gkPbsnC8Y0f4peKqRKKRFuFBB8FbZEJG8KBO+Zisf3
3a7zHVvAgf9gEeuFPhA5w5GVL2hFG/jmjNwH2EJnk+kwYgj7ZwzhheQPOcAg8rHQXMpSrkNlzvdW
OGMFL+BCeT6zWOSm1jAAINw/GXpjNAPXK4vF0QjZ4Fv1JhyE5P2LzmPUuOmYRTRTvwcfWyub6RmM
4H2xk7wwBAbD9BL4QAVZl18jASSk8X444+2TWC9Lscc3Oui5PMU0hEbYqpRO6ERMZrIaYEyET9qc
sXuUAv2XRDe94eUQePaG0DoDEIoAvLAVvQbwxby9WuQnFUHTgzZ9zhqAaSX+ml0hMSw/vEBJprwR
GP+3prX62Gp1sggRDQ8XBAdj8mAxXVIc1UQ1c8JqCnFi/9SPafrf0EzWdf2pmMuFnryA7KZiqmKl
yErq7D+bo83VwWuJKDPqtdXTgJwMu4LRVq9fevbLWdQndluUUw+puEB5qrljRCzWaDRJ5o5F4Hx9
ZD9DYpEW1JMtBprSUgp0PGKq5gjDP+zu2qudWZSoUhaZA1n8Zjn58ufOAL8kLr0c+f2oz4+oUch/
xFVnmomWxIx/ejPZwOiTwh0VH1BZBK9OALAFt6iB2SB5uymmRKxeGuNk59k/RCFoZriig3LmucJT
Ji+oGBDfXa2AaYMBIuIFzvTcYkyr5IKKP4WMIcs+Z+Y0Ii9fXt4Kfcuv4JCXB3eZnZfsH6AXzS2G
wzD3BqEsieLzjKohHzLrC1C2RjL7NXoMcj4uOJis6eCtU4SVTvnN8vQ1AqFCIOMCanKB5I77f66q
TERGNAUan+CZ1hs3pzGG9CWmrK8CkiLDpPDRtPSqFjzrXlYf2bcnWeLVJ3VLRDJ7IwZAzU54H5Yy
dmuHNzeq0Kbh9Lj5eDKQ/W9YIk2LSAH6Bk+wnimJRmWQOFB4p6aZi9r9IWgOdDPjzU0/fcqVldVJ
1YPY6CcUjJrOpV6Xy43uK0Kj3KrgKvXx8Ds4V6Nr4LknS8MU3HUMby9jQdIjZVkzWw55KRRRA60V
xyqvPlSuqrhjFm0yxDCdNmQxAYaHxVs5iP7zb1evEnBxIGG8fscQBJmyMNPbNfCfcxbY2ToJtsfg
N1J0z6J+FZbaZKpQkJiDN7FWuHKMlq8PgdfcuWus2TCn/S3leEBHZFovEL23UAq/vQ1bknAcuFKG
CzBL1Ja4RI6b+ZB+Ex2R99SyPnOajCsUieEx3XV2mISdYNwNA7IrG/vr1nf85dxSgINUeyFlEy0w
b0j3oFlE0Hbz+uGq3TjOZs2a+g0vKjNPEXJn4qGV7N2T+pCTvevG5yUmMq8gext+Mmqr8TaDVd5p
kQxAeSQJuUzG8sM0cvpZyEW/I0/8Xd/emY2oyJZjTQs7gWxtQFbzGkBarKYDGWcQ2ojcuzr6qCiC
Rs94xIZ7QAJCD03sO/bF1EnERlfa2FHL/dYv0D/z90jL/vRg04/jGvmgytCdtQGhXyI5PKyBHE9l
7ajPqWZXpEleIZa7+8zUgVGfXOJU/rlxlYCzCRACXdWil/kuULqHO+F/6BQkbd7dLiZ2TbxCCn1y
tBnbwMYp1LB24nK9MlBK7KUcWbb3cYls185ueMHi1smvNuRtL0yZ1Rc7hZOd5drdtakrKePUtC6W
AUJudROyHzESIpGZVuSzJLYPvwQYm3604WLqRKVkTR3ct2P4BmPY0/5FoFfPCDv/KkTFlXpQHzP6
9ga0yUE2xNIpAN5c6tiQnxtEESeaZ/sVQnHBIHD7i8frMtJdMD/uXSCed5FIv7f9whyJslqrq3yP
sKXWoCwVbQSVRjDg4gTrzLzAbO9gFgvjiTWFlz2bCR5TRCcdfigTfV7fV+9mx5p9nvjFUY7MxZE3
mMTv4Y0/rctgYgnDPpz57ktBSulrNl7Wq3Kw36t2v+f024JfwaPqzxmITbnMeDITTZReWmupU7Tq
eKeLzrPDm28k+9EZsXZVyXbF5m/ukItK+OGg4gjPQ0dO8fuLKQaBFFyIEDIX/P0mGEQkqv8aXyU4
NaVNi9oo1FIxzXNYcoxe5eZh9h7R3Wt9xobyxPN8TeJO7eHdd1mmOdIPPLZyEEGkAxkTqEiQUsEP
CNjUvNgop5XemPff5gCM+N0UDwuBBK4Ahl60BZ7nQCTy2XGB2T8DIjnhOI58bDvIpP4T57FfElgc
kSB6BJBQnSxgWFPOBxsTFWoickDosBpQ1sgaHRm9TahFNzoxyzaZ9j+49qB8tPOmuFM5BrK/iJ17
WUX+nFuOZL0LPiCXq09P29W8isrpX44rvvvcyDDNEwC2Qfb0IhmVCFlVRLGNbXyQurB5/a5R7na7
fRjKpP0mJyB0cAvZBi81DXsl+dpiB10z7lX5Q3HfyX3U2igQ80AcWVDBVet4kbNlf07lG+uVYxSU
KoOVBx9AVAjzN/LnbRnTzOfxbehBv4qCDvhe4XenxQEkXdDpY9cNO7iRvtZan/lohnor3nDTRRbE
7Eslv/Xt+zMP6EbX3+n7PkHvyxFTox6g6BSlB2rfGOfnyF2nG0EMVespTzO3y6mLPLirYI5WWdqK
KIn+43C4ewga08Pxu8szput9sWZbxK+2EA3AT3Lzd7iMMaOE8Z8kux4H8gTynrieZ5Je17IbuD56
R44vh+xAoI1d1AxF3PUmzKrZeuEWiADb7CtBp08O6EpAglVB1XfRE+aPeqmad5G5pmLQrUtiqDxz
1lM/wOCgGOvt3O+bbeMa+oZFR//+VBNWRAWvXWKrpBeF1DSucC7cvWN7ypq7/W3jPAK4JrHnnff6
Vn4DqXo5UcV4Sp3u8wypsmC8GqSPvwX9+VGyzu1l609yZuMUc/v7UlGOqLVjQjqYfojlz31HjxI+
8IG7sGJsWbBOlqIhwiTxE7/QzFYoeeaK4A8gN/jNXTpFQy4BwHfiGKdYeAfsC0T6Cp1Iw9piQ3gV
YDJP9tuxM6kMR1mwFRBdyHUmjNUtFDulI+HeKZ2s00vF4qs+dv0SKG3Dq3JkscZ0LBmuoy35W5Kv
FHisUck95dDvaIZptu7w89akqkBizHaR3xUpwMPghOkq57cDcDsFnEFFu3DR3/OJf1HCEaBRM2/u
W8vmkQKSJKQYtc09/ILNoylt3qsQyWiXRDNEyyyrcPL60dZYLHAJaX/GkiGMSv7y322Kls/HSWWl
nQ+UGk/SFFwniGRcInLrHVN/Iu3UzVBZBreQKnbA0KP9wc0Pb7e60ateLKV1ah1NyZcTZ6nKw4TD
wezpJJeSSIbWcat/cfVkdlOkP29ao8AYjzygSsbf4NimWzXS5kOBhWwIctrVXG2tTphfXqaZD4DQ
LJmhPhpFsdA85zMx+rHTVu9m/QHpysfYL1cDnCAiEYHm4sUDgI5eC8JAeNiAWgOMayJW/g+7uxAH
StkwNSOcbG8IQywOUDQg/nNIOFX+XHs/p0DmMYvn5TU7vIbQOQuyKYpa0J3DEHXpvu11gaDkuy1g
6u3WGlETolHhGRI025MvoRzBwZuO/RN55JtR6kegAWsArEQykDyRHC7vbILYQykrK27gb5MI5waA
iuYz/K06DHJlFJQHD6NhU0NOlRq5eenP6j0qREPZ1RoyYDctuU+yBX8Vz+BT6ihxrHjUJ24wcvhe
sXHra/wc8EWg1aREaTwW5l3E8nq0gaRDVAckiS41vZ04y1BsPiCfGAQtYoG6Qp2qlYL7i6qt4kaR
wWRoOqBKqYVESpu56hfGqM6cj5B7u5435xrVbsxpsycDWi/uJBCwEUg3+Scudzur040gtFWLESMK
B2WY6BYzbNAFbVQ2nI/X9fmvk95QJ8lPDDjk8kNnoIJVaP+V9E+pnNHr3FICsvdy6eDeLu2i8Tby
NTueM0yXii9MwbQ4Hw4vsOjE8Oy1fp5Qckvw6pIoW5R1EAhSJgtNvQQ3uktEI5fE9A4wyRgHC43w
BM4Un8AH52aT0I2OqvTN86gw6QPi4roHVGBZ9+u32UcOX9XXWPObHnDVMiR42oK5DdyGS0ESPa2S
+h7mj6o8Rxbx4iNZqf8ONsn+Arp92tmxqtXxv0lHLrErpBJAr8YOkCZkbzyHn6EixYvzjjlXvzat
BTVi9umdEAsASMO5axIf8WLNIVCfP7pyufiHH6a2dlrbVpXTILKmuQNqAaxBiTvci/45bTiNhUPz
5HfYKUIzCUSM7zYYFrZJ+Ppvd9y+aqA2Ird2einRxbuganH98W1FnHIJpbTbqHRdO78TO11YjVPO
whduTe19GzCqPR3eqaw/SYFFYfpPLgomO0f9q7Ug+mTESmTkTLnmhfA4rVZrRQa2LkfbWKzceD36
3EXOk4Gw5RH/BYLhhKq/BC8g0EuNpDnonUa8eq0o8d9wv0VJ7pxowY6WDFs9l4Rx6rWZ0rmj4KOs
eOzTeFrB5yudkIf6IHlMosscaF9M9fRJaGCW4n30ec7N7hXp4D+X1xDOB0oZ6hi8YhI3otIaw8cr
h88I5JzHFz9LjWHNYoPdzmPpXGvh0nMWDZhTY+suWGFksqw6eumhHxAMLS7jlpg2lse3I+ABGQ3c
OLd1sb8QPJP2Rg+sJCttYUSf9ZWVi0XfpWHhHUCU7LvimnF7zlVXhA0lQQDW03J4X/U/mfL6phd/
pbTe6jkVC/El8ikCmrNfp4CNAuRteqymxAC14g3Cz1TkRxnUOXPUfBQlkvy3oakIB7sebfRZ9gwD
Axh6K4CW4fIg95ta3JMHaCUjSmIq2PRAggqcEge5vRNLCJfFe3ZohMSQuTpyT4YG211BQSzvev8S
D4FQowenpcrfwDH0D+acfMJ6kRVG+hwGLU8cjpDTaIbxvKQ0NbF4CpaDL0YQnhOICQiUencIrWB0
ZLwmvA28xQN9FwP0zVGpzD9QHvew+K9zFE3cUyaOFse2b0agQH6ssw98mGFGpfoIMQosOgsf6vxl
1UdX/WapnUwCwsIPtpkVDaN5Qbup76yHbvi+kSzpr90+thXK2kTps8o6fgOfio5XMUNwRPd+vyag
1ov2tZlQw+0NhcIDTe73v6BsWMsY67eFGoxwRpUti9ppMXlmE4rNySfMcBuENIrU4a+weLYffJGv
lkBZn7ShnoY+MA1uUxYvBPz6lBW0/LJ9lfs5HrK5EoUKmCypkddPuVlYfWZ/F1MZzzQIR7m9UlCi
h25QCEr+D2ViRjD1Wg0xJPVfBOM8XiHZI+hDjOBcVEllIYvpZC3r7ZjyCnhzYi8508ww3XOeh+BQ
/1YPDXabAu6XU6ovuQsghMr/6PD6z/muFme0OmDnNcORMRzT5ZXasErE2GYnsgCMQ9X5cdFmpgRZ
QX+dKW8co3rn2Nxkva/VtOWL4amX00tVzUH0zapIvswmaQDGntg1mD22CsOhmjIgL0EOMtQeF6Xg
vvtKUnd1Wf+aS38jb/wYM5zHUuZqoiy5/xakvY000M8fim5x/YB8oEexQk0sG19+fBNgSshyd14F
F44Olazbx3S/DoeKwWTCKHWz0HkhS43PrrVj6CBeLzyY5LvPl+RWOgCA2EexIxybdiSvZU503ou6
O4N+pzQbEU4OTpD8Wb9zFMZAO6T6wMtV8KbdFCZmIHPgKDHO9UbWpH3XHyrzn1CjLudodazDT8e2
oNWnFsAyYN7cgZ0mxpAVe/MFXYPv+51Qeu27zWiEpb44CleDRlb8ochEeTkuHbHhALFpNHF8F2YE
MUdehZiiFHTEoApUhKLwXhKBCIywMauCllgzsX8yZdqFOIinFsqMX0NZNLEm3FsmjEEyPVvwCtIZ
Dk6iOQNfYklGYzx5hxPrvdE4rMkDHZ4jvY23xjKgUZB1KeLfv9KsZHNgagTUAdpnhXC0731VVLpF
ElBlgcGWMsVqer+MXt0GA/y1G8OzGeeouILP6RekYrUBXvNDE3SVdhXeKlOOF4d+sdONX5mwCn8t
u1iOj58bUdBXaXDGMKtVk9DXFpi/Jstp/Puk55k0CZEzzGLb0hRtBUmMiJARs6uRUan83VrOEivX
hD5tCfGJIN1av3UEAVYeB4xwsVwDIVaIi+oQsEx7uLFt2VqKWRlH2Ie+mvxRfS6a0+HGKMspcv3H
sIkc90GtoWO8mC+JjKzIYeLD+XLkmYs8qFyrpF5kKOh5h9GNbrcd3ZtYvKfYRdqivC4ka+8lClis
v2rXfttqOyfoFc7iXYhYOWR3SQrMwGYGy1mDzf4v2RyBQWa40Zrmy0ZnKBM3813pwrfz8LofgXcC
sDDv5WL1yZPlWAfS4y+q8VVIoAHD3BDDhKKa5nh/X31xUXQ/ykqO8JOzf1VRCxrIE5gwZIOOF2jx
uOcdug7jT6wlJXQ1PM9Kb9dMUikvkvJIxL8SOo6MqGeXziN3Ihh+0m2OBDcLTsVFFsClEWppFUAi
XXtzxJNnStUDE6irrhx0JTEqteDXXg4Iz93WV0LCT8HtZQBQUtLyx6KjObN8RvD+VshU5dEG5KXT
CuMsa7g0mwnMAOD2W67bPkc5w1HMQtSe2HjnAe35uZRERpcRxIys2gu/oecxHAGj21e6taQLOWs7
wo0N5wK2u4k62QILB3I0sw3R/PBRSsksOmukAR5XJYAwIrhF6HfVO/U0xd8wdlyS/Qz4AVsXMwkD
VJ/bsdwK+rwAP69QVVdVTHA0GLDG1J4S171iStVLd1e+nZHZOTKq31NAptwt8R+8KZxFxv8YoUy2
TiQJXpRACCizw90KLSRRBNNpBK+elkfR7INtTJq8Hbeq5L3uXKeN5N01GCYDE2fvWmnh8WU7+OyQ
nZv7GfxQID1Bz33I3zjDBmfkF8H1ZjM888n4SyzS1wB02tah844Wka6gc6Nqf4vhEgzkg1fDm9lX
Bdtdf5cs3jERLrYWQCRsYLoMSTnStllP9LAyTvgOYoqGkwq5CGhUkGhS5xpzgFSkykVCyZd3NoV9
t9Wv5RetE0iuFskox03fvs9DTKt0nPsGD77UPWsLKbpyACEn195IAT0WZMzaWr5waAppAd/i6E6y
l7+KMNtjV1U6IamrCc81A09WAZK2M5kI0xPJJq/QKcZFw1vzYg7o9mbExBa+eAcnlWwWIHyFOx5i
VH31pBOT41R4Sqm0qTxt5HOSHFRdK9OGOB8YFUtpLXNTKnXxid6QcElkwzU/8Zi+qksWR4DHEpgK
s8ON5kXZ1HFYI/npYLRslLQBMPtJojKI7Gg1BO/Ijt+9h5TknXvhvCuUmmp/36kp/vDe4NbMi74D
/RseNAfg66NH85L3qgZBUDGHsVObyrwOqjQsKSkjhogXsi26xuSTAaJbIEy5nbEbJo0ijG1rVChf
ZVoLH6Yyw5QSGwRdg9VyCcpNTajhPY3B6TOm9mIsgKFzqKkBb2sU448JQ97k2/b18k/SNcf5WI5Y
39DfrIMszob6N5lYfGrocWy46ySsCCOfPGT+x0MZ67DCw8Jizg3Y2SZ+E3co5JppjklioSRCwyul
F9+K7E4qO+j+sqgRFpmXKgDA6KddeLTkOAgBdVNKUI499sys/qf6GwqlESxFYOD43XfEUqNijTYQ
1HZvRwTpaZXP8b9lv/CeJBRAtVHb3nUqSoK6d33kdmUQ0p4GSngzgUHiRDAef3Zan89bN5FmT9K+
tjXMJXQt24r8WeVX5Orwoh4MVWHHCCv70BXAohSQCmum8slixe3BFZvcW3tW5TwFmoXAYzqZFm4+
sloX75s8Lhkj7/OC5jjOXNsagMUPiQd10t9niQg2SEEvwLz6Ev2Moxz0L8Q5Y7MFnNi9O2y/lJqc
1D4NzEinzoDVpaSgTAqYSGWyd0mZlrC33NuoIqA2il7IxhhXienjGGmhHUreBx30j7XcUfg8Li7I
uIpE59N+uQLyT6np8dW5/ZR4ChTjRvOVD5s2/z1P0/ME7lwZGAdaDZ86ST1jjTVU2EcemHkvmtpP
AerJfTyeD6dV02wqT6qiQebtTGGq486UmpovEbOQxPJm7QKiDORsZypWvtWd35LL//ufMDmzJUWR
de8rau0i43HvOd3yxE3+OAY1KyBelbs52SOxOvm+k3WYsoe3H3Wpp05sM2vx2Bxqjt0Oh0nzqr+d
W6A6cutXmPHvmeZITjSvshdzmj+Cv9mBaoaOgQ90G8m/JVx2YHd3ZkdTHlW7k3k26pd8Y+unw7W6
d4CNv6ySCPvqTItjZOYh+wJVbsYB6J9OPcYwi3N8AdeIw3YIvBFr8PEzFTh+sMLLM0fsoJEreXuq
wz9SJst1u44rDn6Y8sJluL6Jr41RPv56LkAQzE1W4WVul4WnhP+3/b8hXsHo21fxt2+2OhQze7cC
NK/WgRVzCeYVNSQw6igoCieC3RcSRRUHF8jPevReWSFSRojlOPp6clneKEq2pew3fhzp95Sh0IKz
XbTsUsNWnLLnUfs1s5sRtb6ryWuQexcKZpx3EYC/HnnSnrOgsobUkvzKeaYboLHLXn1EOj8RsigC
Gu7EcPKlmSTSF3wmmXgzOHbCNXuyQtVgk6Wu7y3HUEnJEWrXYGz6/ueMMI0vHrwhbafu7X3eNYrd
Vkvh7QKXM1LbyQjALWfGpfphPrBV7l8qj7PMMLGaiN2CScy5dN/9HStBZtKnt03swnb/zODv+t0X
IHUPG6PZH3jzpzzQw8ycKFjgQoEZXcOMVh5p2Coe5+7Zy1SK05WJnx+gurnhPWTZU+O4/8DBfw6m
rzJnEJWqNRhB9VuyT3JZT3PoRxDfM6L0iiRLKMP5FOmJNgElZcFZeKLWds5e7J1EGpVOlpmAdoD0
rj/oLP4IF3BfpUc0TncjXklTIzeHAMUhnjShtvxXV1XmeT1jBHf5KNQp39jR/BgvoVxqUpX/QcPK
ijhbWpPtb2JKhEWJ2+xnwtH4aKwiP3Kzd/jReX1ePVnqGXX3y07yXfKmGXV7lQrwypRAvtS6QLyG
EyC60+NTJsFe1C4PA5nu+uH35hTguZqSv8GAgDdp9RqbX4FjJJasQYE8o84AwlurGtmKBK0U9FhL
i9GbmRzwgfKqkMsWb9tVngihLTw5+zobgK5GRoEo4qDeQfnpulxuf3fxSXOqk46w2tiAK9hmn1s4
Jrld8WQera/TG4rpk0fyOCKE5z9N5IJxnA2NYwB41B3rkAxyy96LTGmHMlFwBleYOnkzRN1Ku2aQ
A6JlonXu2CHlXhTK3sEL9PSUMAKOClgkHCFd8Z61sBcyKpw4G324q93fPP5ujnEjgxkSrO3KEzNc
Ox6aGexIw+uLX64FZlMx7igS7dIBPaPrR8BEp9h5htZCk0UOHtMhwQjZiv63MdDJtzIuF6duOJ6L
Lye2Oaw8srs3AvS3aCqBu3AC9Skjzf3Irfjk18N8I5d5dbXDR22oOmKh1MHegWFW8YOmM/039J8l
iOciI279hUrLLBkMTx7aiUjzeAn6qrz8z/XmoRDaFsLc7ke10qiz5XkdK59CDv5I1XW5jAtCGkZb
3YIZGTj0oKi9LWgQqtEpfp4QFB0TqKx5syHNyApUJubrMGHLL9c35w/1cJ6+f7e33+iVbvuUzWMG
qMaG9jSE2sDfkHUgocBn86F25he1fNxbHc1ZtV72lUAZJO0Zpieot5em7VB8+q/3QE9N8vQ9Y8VC
/u4fFaSTaIpqZpNYy5kdtF8pAVIOqDfr/PT3jhbx1NWS8MvRWnn+r1JRYJJXKbk/Eksc9pTIONHr
5P+n1hpPC+rTOgXCg3iHJSPNwtHPIoBNrD+/7NgiPjFDHwRA9+dhdyGFBjZeTZ3vqvxfthf3rl9q
u1xEOkz/77Esg0FkNQy+7aNjWFYL3fVGXil3w7ke+xZS23hcvlRoPR50d/rJ6NG7GNcSr5rDYr/i
H3wxPo2Qmkx/H64WGsC4XQH05ZhzE5L5i8pRfhz8O/6PZDr3Hgy2r1PR47wGAaWnuKv3gi9zLzqu
GOyTzWjth8pTOcQy8AXZKm+nZMNkT8zAHQGZDPHDv66N5VCt4vLmQM96sCxy1WlfCMrVplqrgFmc
vNQJOyGE6yDDhOTZfpVCt/Y1dYhigRDLZO5CmJBm9Ixh9YQouiBJ9lZWjcFawQNbSTrCSEPpz8ln
35A5OEFEf/vhZ4SGwDeAuB0m1afHa/ydBzWBQa6JLTvpJMnyg9Y1IuxrpPz7xD3ZIP9TQJxkURR9
A3IQ3CCrW752w9+A1ylpOi4zDxKwstOPqu9cclUxDiaMq3R59wiqZWKeVh4H9RZvgGlDTN9mmJV2
PclzIhwBnM5xryjWy/8w0vagj2SCoXGxBuYd8wZxXoYUV4jzZDz9/8r+waXYxlqGktp4JZ9KA67H
pzFmE9g9qmRQt+Mn1Y45K0XL6kg/1VC6X8T2UrELcMHfBnT+m3mpY4d/LhMaxM0qj3SB31Gf0Hfg
df7U5QMm306dzUV9dudpdzG11jnzJ1XXXDpK18cMaRTueF4/fXmhxdKT+/ESdiHC67FAjZEzNg+f
2vzFho2579mgnrscZHM2RVrOCCJDjXrzGcufGs7bJomc79aq95kJoWmmr6bk2zszFNqg550BIo/P
8NhsMh4BWQWyYAs2KTNPp8S1tmsahCXX4aFJkD4mwzTUsr5JhpiWpy+xlgJ623jOF+k4TeqRlD28
FoJ7SJ8XQz/t/sVTYyBq5BJo4Hw5nEpAiIQF2vzbH7MZ6dYbOywdSWeSOTCkNyiLFjrYBVPEMQmo
/3mxj5ThkJMGp3NIxjRDdtc9L0Djh9DBqposOF9FPd/KT7mQ4+PcZsBZbMxPh7ol5aX519VyzSnu
d300W+ahYGPScQjVcviAXpxt36oqVYnCtK3/CQi+R4ihcrsKejVCPQmJfGhSHsV+pe6XwEKFoq8+
s5c6g35CEJ+l6DBcq3gQBNHXHh5SyOKGwvbxoXmKa8ZH7bgYrjEYUh27fTFCS8iK95qpqG+YifoU
6WLg8UOE7cSWb4F9upusS9PcJFBbxLNAuXrZc7/LQe5NEz5OD7HvIUipJdFeibbJrHXu4rJvLOch
t9e5eTPy4GDqI1IaihdEhngxlhdvPDu/jPD0rZuvAuX06tkXtHS7CaAPcRqX8WndgoMhVvrDdKen
hWduoX1k167ux2CdyT/WstAivWFtw9AdL6mOaCROqdvCekdNYXdEg+ocpGfm5r4S59x9OXQdvKAr
erKMfEh5QmoOe6axjTnQuG2LaAyT4bBZWFJgGQFWUcA9wgWtu7t0s+B2fdrJPij9h8y5nifUrybd
i0gm5mGrg7dUzkt/vyrjcggeui1GJmVrRDdy85ZmIdjJKmWpdcUwAUSM/6Kkk3Fp+uLXWac/YSf5
a1ZvbJlb9TziwlDdySmd1nYOA76qz3XM2Ma/rFrN47kfVNy+JCWdWgDFtYKBMCE/Z3/pm/4NCoUx
OXocp+BGc+r48NbTv8QrgtJ1BfSVE0NHknhyOtdTtFVpk3qY00MY3/RkhHIS/RokK/sItZ4cwq50
dcrCdEbw33Hom7wJy/YUD87F5pFcZucSUL9yaMEVQlg55pv9q1G5wJEmdTW8saMqqVcwYZxRPt8p
YqodYEYTNISN62mDvBE2cM6/MK/PZ0qkCf/psLYjtoxWSoXH7BuWQ0adsLUEsgQ3qCOWcKMFTV6a
nfm6a4hL1+uEU879NdVr83S+92vRhfB1eF4y3VFVc459lHQq3Js0ErYWWiHihEEjfbIB2a+SMOvD
aEkRYzf5Z44Mg6vs5/GZxt4WcHkcuV7n5XWH29DkwcNk6y5z1c5oJ3Rnx+CoZkc3eMQFdWvPV0w0
+ArbPaG18d72SiyKmxC4iyY6ggCkT2CIcrytp2lAJXBreTMfLJ45++sxH9zw1lz9qRItFVrVccr6
UrHzrZooqk187J7xpSRfA/+fxKe0OATzJYLJGDPpj8nIDnQGDF+8zEvbTdEZkFm92C8PU9VuBc3z
lhJ/oCSJ0pQ06uX/VWVe4pC/8p1jiwIEoS5qP+bYGBa6gC5Zam4/2bzWsgaEh9R1tdjmnH29n3bH
0lDMQnglpOUf0BW4rypAjAvEaKT06xObKnyGNE6Jv53WZzpMh2gCLG2XMDLMJHn1LP4SPfUkAKhr
JUZVrYDmVQ8avfX+W/NFJGpHwWIPK8osrCxBKVuvBHJmLQmmZAz+dI1UG4etPnNn4bvqgajskOU7
R8bz2BJRxZGjwys52Qpb9r/UcOZqfyL9ZYO+jun8ECYq0h4gQN5hgocm8kWBE1zjTqGgZwm8xozO
5EPFK3qQIz/VrrrP1b0V4kopQQZOeO9yKPonyj9M1Ff0kDrb5AB1XSrr9TEFw00gLly++m7Lo0XK
zJfYjhD1DpuFGKpgZiClngCAXZ+QbWzexVDGElrIRPstlVWwW24it6SWK6WlBeKZvdlQ/a0u4BwF
eH7d1C9S6fXI8RHdfcFoHAlGYTLDdyVAeJi7+I5Srx9AMkozmh5+8I+K+Q1lZlzG3xOVHLTa5hEP
AYd2BywAxjkKDRvP99Fg9GmeMyvUCRtg2nE9spKxab2yJOIDjZNV8T2cisAEu5ICprzzg2soDDtg
lXzPb9kBUUsrGAyON2DptNPbgrPzkv7crtKOt0oriTy0bQAepGHmP44EW6K7Ot4Z1w01Uvmeer63
cvaXscyLpDiiOBFCDhL0a10LFFFodY3R4az9wbwc1/fpsRzK0xpPNHSI3wP8cC0gCXAQxXtRvPRM
2k5rqumR5JE+szQUkt2VUNAOuQKdldgCffG8MVBWVgik04Cu5v/jTnqHJegIk9pa6CEnKSItDCkv
0xwkvfLX0kJLpI23UJdw73EIrQ5rG9sso9j5BjSjtIjzD0HXToKq0JTx7j+xKMuHWbc1ALRbPQlF
KrG3ZJXtO31Wa5xuV2st+v6NAm1dx5NHtxsFwgEZPE4durtlpoy5QN9/v/zXmy/t3m+lI9eN2otX
N1Pa2fCeakcCKpI7K2xg1kL/T71ebco8wyRNeuc1Mu3nUUWdB0sMk9Pzi3zCbVWQCa2VdzYkEuNz
lAOZrQr08I1gcszWTKnjjBp6NBI4yOqiadxMW3Teb1jb3YolmtgcYyIF2ekh+u/g6j9+lvD6aQ4V
Pr5Oy84fr6L0dJPziMMyFvrd/ax7yM/kzk+SwgNtqmCPNIHN5Mmp/t4lpQQ6xxdIsvCwRnPySmFv
RFWUmFZzxbQ+gVFKdCWsCpSzywBA3EhDgDxVTBdh7ijR/smeu8ma/XPz+RNHlWscXMDZ6EmQFRkN
Do0lhRts3EwAjNzMyuPxS5HMNShPv2HmbquBT2UQvXGgQd3UfIfO4K1jO0oTdi7xDpt1nCTb+Ytv
bUvGKezdTisPjbOsmhW0cHn6jw62xIWolk6ep78KUONzgcy0+NGtXzxQ1IXV0HnpXLFGX62tvZ7+
oomWvqOpYRAi9vBM8tnexuYczCoB6OTZpPLg+IA8ws2Ypv0k4FT7aBo67ndeHf+LJK2GDpHV5Cc6
UXBGI6uyOdmT/LZv2rzszygbhdKyMDrLZBAPtjib7ou+1+oV7CoJ1af/KeJ4N0S8DLyTD5pH2A5M
ZWFmQ65HxxUxsMP2CX7skOGPqmVZTWWzoCekCLooOFP5zaviog++5Alh5aDhGTh7JgwamAZ3B5iC
SXbRrKXjaluyB45PaUhlo11TljnkxOKB4hv/IIGwM8rmrPnNwV0ZMeNKDhgzlDAXEskxveEe4OC6
B44vThB+29gKCBKmBetBLSH+drhzQHMs56XjFESe13Jp2OFJeK54sWQdg1Zab7x/9jUkidJPeXLr
akzaeXKh6xOr9AKwtUtgryPa+v39aXMdCZs+1OvG/a8aFESMKc6LOfrGiu3MZ9pLPXB3edGsIoRQ
qq3QoD5UyHr0hJuPP7V3FSNNw8aAQVRpOs6Akco+YmxU2zwBtenIKLqrSfxyG2Hcmw+/hgrPDoN/
wnuGjJvBuw84DKLp2vuMApZMc2KvV7VJRp8ETiFpFCYzR7YGPUhGswe8NXd5Fc028DfDu8uixEgm
xV/1hZH5IZt0ioTMhbPV9jeVMBeIf3C++be7rA9dvlVlkupf90yRPOTvWvPv141qygBtZnV5A/mu
AsH26AvKA2gIla3eDST/PFBxeU5B3dOM7sUyUJX2MHcVV2b85ihwXyLb4vI2GLXIgWWixWazZ6wx
KvKKHPtsjktpWCTiqANMxokl/jWfvQdJWnx6qgw2epO4ci3gR1PDIT2bjAI/bWm6uAv3p3HqFDRj
JhHxZ2VBq/g8lhcpgaC7zmXdP9fTYfPAct/kCrWSwLdSx2PeE/mRXV5WsAOKes/bXdSsWWUtsSby
IGn+gbvR2cdHbFygsfxwv15lg4kuYI8dF0jM2nTvEJhdBw3HZYRWCGn1NCxh2siiuJ1cC6ViLnZP
+w3HYUvRQSA0xdBp+06QCj51Bb1JvFLT8uZ8mqUlE20Zx6FBoVQjiZ0CNg7n9mk03jDEYxciSjWh
SsoSn1ZnQEByM2BVWUz0EhIal3Gd8osOWdu6PcIGXJc8VdL6aVnDLDFeSuoJpeCVoKS1c0u4CW/Y
JAgUy+seDRBP/jqv9HAgv76veZbBiNvPFigVdL9L9+TaeUCKSEV51jNhJfRb/5go/iU+s0o6maHq
HoJOPq3sraCjgOZXICDmNyHQfbfgR9HoyZ2nQNvvJYZZNrGLon9CwGhu0EpEvampEjReeuOW0ZIq
ta7dLrQCyEwe3zfovlYgsHYfgOzS10EdqvcFfNBYpYJ6TTU2PjwQzRMFujrdql4GuE/4JVxYwSrv
aG/bjvoXGbTs3jfuT4E9opu1B03GZ5RkUrPqZ3+lxaERyCiPl1QM1Zjfr17Bou4k8PAc6kxDNEwT
D2YGEMyrziuDy0VTjSbxKGpggsp63NFc6dN5ZlkO525gr8HGB8fMD7aXPXD76WBYTWFQfCkXgKW+
fE4nPFWmzvjaXODl/eMC/LyzQDBP5ka46x0sPkZrFeN0asAPle3adTLjzWryB/llosP3vqKlLZ1/
3rF1aXQodkuXi9n+XVsTCEI1oKMn0uSHE/Kflnmfs2vjKaRn5IGF18M4ff07h+wY5YIQ4uq7dQpm
nZwhxU4vPEBG++RsSm6uUg/8f6obFzwV9MZJ1fRz4V7or19kFcpOo6ZU5KxhKqKgDxZMuxS0GhaL
gsEgj9z++63E8FgrvmXOLEnw6XzJIgeufw+LV+fk7HcDz9JXQpigx66W5g40J7mdBFFWl6l55E4m
E5NdmFGZinuUhWJbO8iaGeD2ceQbFZjDwkUEH7zNK4A07lhv3T0uKnsFiS9lvEOBTnYfHolD0zTK
E8HOLAGIHqXcJwv36uMKs9otshhSRgjqJWG24h8iQMzjZMol8H8YXHUQyugx5nsl/ofq6m/rUr13
GWVuwvSdt0xHt37pi5ldiummAsqhURfuW6/WwPMO1pJN0KPSoG8+tbonPxvgwGAONsPAyJ0pSXY7
2cFNETArgU0vPqZmiBRULNKuWzfkeqladJvkOOWmGB09lmHWzWnHRUOVqc9Te/abzutAEImV8PHQ
hW/dX75Volhr50IkXl4/ptIxhDovgdmT3XMAdFMUTF/AhvLTZwbmk/rujHWLVtWgxSttqy6io2o/
Mwi04NSHpRVbupD/u4o+EKP4HBT9XlODmwdGlnG6+zo7f7rCrkbfvG343/yQ7ZuJ/EsHYV+B8wBj
qYUG1NOvzlAr6AIH6ZWMGTfAy5Y14GSi2E9RLOtm0kpPJ/OhpIh8cbZbhm0rZhCiK9yyCaTy4UDG
Og6akxAc+IOnpmLYvLkaoEj5Z5EqANcmKf/S+sPR3qJZf5oZOYmJlH8oTRa1GQtinyl0cMlss+om
5+s0I3XGnH9KwvRcTEZ4QkFxwI7vRhPpVv/sFU4FFOIxtE2Fg7drH9QwWSdzIy07WudaqAWmTPt5
/4zY/iQqW31Wb6b+EVY5tsJvf8UHI4TWcismcvhtaM1A3yWBbkPMRXe1Un8TMYgGRlvah6yTI5IA
5zG7XxjxydzN/okXcJbv6iqKAiivziO/d4r03OarQjR4nF35NRx3aeL4rxxpU2mauf88jSxhyN/U
9VOl7U3PPehJhv7UxdMWdqaVAGHwf7qc0bOV2my3p1aJRp70U4On5FnToSBmXyHG8HG8FUJ7B9mP
qnM1VcTtnieIIDqe0qa0CmSXMGGfxqnuDi+BtqOEEpPUvIrmvZEQAJ7eWh42iJIzGvq6+NUXaGkc
bnqNArlBLg8QV5qI5/wRXnudnaDnTVptPT6KOo6NoC3pkilpqNoQWelJQz1dqHW3HcmjdBYdwEtA
wH5PAkFKxzgcKtwakOzWm5jRyNNZeLBU2/U8TJsSU8Ai1eKIG1x7bHRShFw3FSiUpKEKnINbTx2k
bTYj1Iv2Sw3jvOJX5SaeAYB7skzRlhCmkJI9crpkNmerpWBHymlqGH6X/cDlFMIM2FFC91JD0szD
JLrV05aXlkHHj9Qwv+Qr9+9uJZlQAcSSEmUfmdfITQ7W2bpA39/SQfWcnyiqldTKmDbTGknH2pmb
xaYowzYJSYAzSJ5ZbAmYHe1q6s4H9zw/gpArj8c7ESYTG8Yxjv5wQUZDCPfK/u89e7kYteqJSZkX
SDSP4TNmKqq5SRYk5/HRt2NXy1howUhcem8cYWATKsOP5iTIg5zYwfhw3Pia14XNGdur8NC2huoM
gHNAjE/o2Pa38zm3mleORet7pU+qyl+gzE2mUSo1hfq9YufMuPOr5jnqDEyGJnhqD5YjnFqhTZ+B
AFLj2EAbM8SDPoW8tmAl7AgwCbEresx4MWPRy+gOiu6+A/JfbRJhfEekckTyoaVvD3js1DZ7D5RB
PuVLa50MAjqxjLXx5kH8R0XrF3MH9D0PY+2OrILEN91S1M2QhSjypqgMuCoU1Sc88pE7NKaABCM5
mNgCKgNba8BlB7u6vIJA14Vh23ikNvxNVfyE+rvUWVrCSa8o10pnhLcNEqDTHT3SuyfGtOxe902K
V3JLVad7r+s477EzGtDuFzPTJxoOZJMpWWK3pX2Z3Hnkn7ubmhAv9QA6VPvTXCbSh7pT+o7Y9uwe
zkKkZ1aeW6OmEkRgbiJ2AiUuM0QTy1qTOyyUzSi3sR3VK4VEM7NYeiJN0umeesX5G8Ndynk8O0PD
iw4DamCYOoIUetNGweU0SKF1pogO/kVThI4GU8JGBadAeFZkLDthvuWdZeRWNnGoqyf26MFSAmpl
PUEE/kdhfBnkV/TJ49WU4jWGJdkKUBplSHSarm5FquLzBdrg9g5lYhxkxKDqIzJav0S9jIKiO5EN
oyaiLFcU0kajF7hbeDyC2apxxTImPV35MWATsqDfBaEdKDWRIxWgzzv+U91S9zD9cuxbkH0m8AOl
+INFP98xNjgofbZFy0c5zHcBO8EYfe0EIYR+wxxSdX/ckEV3ZRR2L+ztzTFph+vI13XBAPfPAbCS
Qw3nTlHuoImDjyviaiEoPUIzAdvQYS8shKwe+VmCxND3Ao6zN84Nqo8h/jGSWtNkTTeiVBFTLdMA
8MpC6g75eHKAUr06ivENHPiI0rthexbVdR6gVB00Q5wyDecIz47z9/mexgPygno7gaWXALfVE1lU
yuMl0QWFdSq4mfTOE8H1hAR4h6HvTULOOJv+8ryPloZPeh98KVrfOrmbgc+kbcfobqvgCgl9vIbU
Drv8ROP9Nf6fE4yd9IHN//ibQBmRwttvlcJUFSNrQIdt05zrqTa/2o60acQiPEQybjQj0GC2U09r
FJ9mGYHXVQn1ccwHI2AWnHSL5G4oIV193MKerb7SQQbGafc/sCZd3GcpOzeR5YWIquS8qHVWG7iZ
kITnpHuoC9urU6Y0WoHuKkkk/mIiyCOZjIu3UpAP9iDsT2Jrfk1pOG6wyCq/4pWR+WEgDS1QkbNw
I2zgCZwz1Iff9lNCYQ4MGaDyncqs6E29+/brR+SKaGFEbyJtLamRCl3qss68HLLHJvAtXlv1/Y13
awH0lArYL+0IQU2kGGndj2wAyHWYPZvuaf4BLQj1tTUltGtDDgiETDBGBNgzGLnIGilwLYUt9pPy
eVANyqTODZ5f7AX7TRS9oiEayW0q0qQYRL2rmNhbxKMr+gt1A1402EmhH8Vt4qk5mVJ47f6hN2Jp
YZ558FSGyZ794JPUBCXiw698OyknMXqSQxrTyF229umGog4SrzW9TL8T5PMBzo+7/QxreqscOVNu
77POX+gavNBj3Ndrq6EozJdvMtaRAfrQN/cBLX8yWR8CuSHNmeIyMhY/slvr1Yz6JxfLNFujKIjs
i5jaiZ7bsq3ldlGwHZHbqhVkmx3Py+ZS3jMyIFh4Or9LAkuTK0nYUoArDpIXDRtkpYdb5jUz9VFm
EezT42a9DeQdYsJTL3pzCc5inRTcwn8dk7tRzyGTKugTQKl6a1X/Ycd/6J008ig9JMOp4qVTboCy
HTkRIYpwSIuzxnSrFY3pYJS2WWVQC+UKnNpOy5h564OrQlaKOg3wNqpoT2MFoqVCFrt3p0Beltig
0DVBaIPz2eVyJKRjZ8NroA9OQ49AkYz9fpcRi3BYmMq8Gf6Lqtsr3zkosSZjFOjDh0v5eYBneLA9
GiOuCQAh0pSRWSn8N7K/+g+NyL6sIoi41MRu9LlynAuVrTkx6Dax/tizQbqAAkkbPsp6L4VTq26Z
0zr4HNkqwNntve8vRJeJy4jMQWlM+g3yZDBgVlrg6VaOUFZzJQVMW/yAyeh/tiKT+31rhgi9qerv
rvjvyYJmpHsURFj1t1ce4EAI5SSa2fzQPR3xEV2m0OYgSW54xWAAMcKclon9H1/dtn7QMK4W6kd6
UOZyuOKOi71aaw/5mlac62gm3F+vlC+yPIAycpD/aJM6fKID5oOMUOq0jFkfjuQdDeXkzIQwxcbG
5PszS0J1eorUe3FlL9gNaKaB4ETxkkSI3tCdB3Jl+Qt2PHwbCDPs/2Kuv3xCKy+ilryjLpFza/k0
g7CIDTdLB7tpsrGX8BZ5jKHVrRI8VRJTFWnWRU6v6v7mcqOEglfDVyKnnm8JbaWMWGQpI1vJc3BM
aiTDyFKWWJNIWD0hM9yeWcPuMB7TaRgRytU5cBEKPGAGD8LbWHthfdI6v/PnKNpwK0zO+pcXWlDO
dEBFFmHThlUHfQvR75ESTrUzNcL295RX5PlRK5j0d2mgNygGDWGiTnGfScHNzYZZnDI67E3+D3k/
pAPcHr0Kp2uYAKYcVbiObwrZ2Q8hu9AFKnDBZvDvAxhYjBuN9Gi7VxXzk8wzv7r40P3ZqbdUdYzD
GBO/+E1mgY4cRBKkwvILlbwTvjy/KAGgsaF1TnVuiKld6rLXC2gU+mxrruAcg89DdzpivkecbYwB
jUXY9hoYRaPLQduhhpaMMkpCvV2ibh9k4AnG7vW0b7h1xHIrRk1vQk5pkGTaZc8qj3IFhvz/KJqV
WK0PRD2uVCRZKLNPpR+B3+7MyGlJTMi931Mq1ErlXreSBK3kB8rOKboHfkMnLunSXnzOLqlpeU0i
0J/N8Hn+CeoPRyL1iXnkIgARYPnJ8cDZr6ufLxBFOclI4AHGrM4LAFlukoVE+0B08rG4zLdxA0Lu
u+OE8ZuhjOu+dLnO4PyukLaU6XoSqdCONTzd0hg4theju7241ut/sV8sV63+81DNHYLOF70RiO9l
0C/9rbIXaI8E4W99r71FmCIZGeCY1T8oKqmMbAMScpOtI3QaEKTIrHWxXNvw3d4ibcB1/SaFJFFN
f+I5da1dEdXWZuUnUtZYQ1nmj00MDUdjA+MUqAOmMmzxYtydG3qZbIDeIRc/WzszU9yVrOzTZQe3
psLQHbKpNQAPSo2+7Io5NJdv7uvu4RfdHc9SBQzF2KQUnUviGWvtmHaQ1zXAk6G/EVU6Qmr9KPeG
95JZQGhjbGL/9R4AJIKZp48Rr8F499WgpAvlxvq0LMP0PVlbtZQV3F7MLzOP+rtXB33hUuNSMEQN
KjcQhHKDw7EdqKEoER+EWINKhgIdRAjo6zwZH027htEe7kwj4FGWnC/vPRkPctBNzsB0Q6U0loBi
l9lpI++I7HJW+ucfpFdXgFfCLtguB/GCYtvgq9K0mUgfc2UsW3yoHaduQEsMxy4qhXl/rgfQDPw+
aekuh2dfRNH8t04tQsOSbixE1G43lCCfGmQAyYA13H2Z50NXBSIoe6zxlrZYkqhJxw3uR9554mDg
H27KnX3FYcQf/UNf5fOqUyY3kjpVY9caOf6fqyCjX1AIEQGoFFFWOlhXryspKbD7FeqxnB6uRCvS
lUVM9T3ysFR6zx0OH5F/BRBGKmsBdJbrgjjiJWtA3EU/WdxNV4rC8Wl2Jjd1WeL22wGfffBRwX5q
VPe2gbyYNKQPnuONtVQ5t/Xqm5Q+ED4Axq3WnRkyfgOM9vM15rQYywX9pXmg2bEraZoV6mZjvkYy
41wHA/K7f7g4LZu1sgcZrUFYKzPZ0PPr0lgE0qom3fqV1qSls/rqdF26HUfLMsqIT7L+esWsQ+QJ
DR9oFlvKWk2M3qefa9LioOGqiIAJw6tdTRgb/CiJ3NFYxe6npTCmJ3/4+88WIDk5kIAeTHsVmuZ9
ZcDlpin6pV1Gl136PK+6AoHMNyeSElcNsrUMsynQkol8b6Fk+0K8jm1I6Q/cLOif09aLqnsyaPWk
bZ1qmP5W5iDbm13Jq/rp+UNp2B6o8Se62B9wClk3mCLRSeFRxozEmrKTkfDNWz/Q9QJ2oAPFXeRF
BXndjepvj0OM96oNFkpW8SVrjItbtRiriUL+GMeNMvdjSHh2LS6jM+BpdtEPpVcfrMBrKzbnSXZM
WEtawDnS2XMhaWpi6fRmNhO0RunQtENxsJliunstzJMZSlwumjSg3B19DkQfqOWwH3r7CLkKTnkY
pn45bf0OymmshGjMOVlOaWZUWRbfz7lnk+rOb7uOdJoCwoNKi5YBIN5EcSx+CnGbieoeZgl/4wEf
3ZnYY07aLu9NeITPJfPjdORyfFNP/9eZ5AJPdaI+1IdLaChAtntoUj1JoeI/S6YGG4GM9EFu0150
iIGvf4gni6jKOH5MW4FYZrXQdtoFGs6O20alI30gk++JPyw3WMo/0eJyCZF1te9v/HOw/d2LzRDS
wmjYWHRJDSk+Juq75IEIRJ0PwP+abUnT1rTz5lfexesEGBN1vjdTaK0gIDAVpMUG/mk2ptLXN0nQ
2cJVifYkL7W6ZBq5HKsCdhgBpgzTqLvpM0CU+gDYqb1iJQJLZw5/xrIabh5DJwpOpoEDdmPcZ5Bs
1IKP3PpIkwJt8yU9KetVBheobgCyjfsZHrxP5Ahbel/tWCbwHvqbp09u5tc9ia9ugaNfrxzhjqCw
kLal6Am+XMIQLHQMFtLeXCqDJLKBMJMEDTr4v2UjPP3LGSV0ykXNeodH+tAWOtKmg3moIy3JW45o
0RT1j0AX7Kcpn1LMASzVt97BqGDV8xEg5t48e0Ypd0bLlTdpL3dtVxIjais/myjXWNO+UkJT+0pE
VrteVszSwU7Mn2BgA066FjsTxhh60/XvE2N0gKDn4AHNXRtepQsbPS2/7OFWUro62+uV3HjPgI/R
sAVzzjHHhDS3oTMa107aZTGdAo70zT39u3Du/gOvb7VvWlwgagKChrjw+2WlVT4r5I9EzGE4yQNQ
T5bGN4VQWkdZx3Qrp0BAI2j9p+8tED2jffwWbQnwZadrLsc1kWeEME5yuavJIVcxLf/F0UDZ9R23
c1Rx3i7hu0pPnpPKc1I+0RSa1LQlxtbpIGPcyQDZm9ScdHA9R6rHcxgAotZr2Wv1UosQYXBd5iJu
yObmq3j7MJE2mwRF/KBj/OTR1ea4KtGl8T/MhFS184rG8PGkcpPBpN0lXQNdkVdmBmrdg3R0ztLD
URKteayEcMfslOAum9HI3Hu2e53gEWOx+hlSB45KZ/uubTbUqh6S9419wETKSTJ8/xsR7z8hywm5
plLuYqU9yaovlln9NeDtbSeYKF9d0/YBEbaNcA2RX4kInU8cEEWjhO5miw1q4jMavmNXtS/tciKt
1X9eoT7cKGDVqIE24HP5JvGcupplVj243+niInDWYLnUVLggka2WlsgbHsiquVj3eTLvRD1GbUIC
S3muUMQGd1L6dyHvT/lszfdHzts0xKe5/O6lYv1Q4GlWMpXkpdsaf0vPGqUFSj2qJVh9uDhqxz2t
u8ah/rg865W2vyAr6gbPzk4owPAumiiewlq4qi5F5PEOx4qQltufTzsGkhHU85kdkym6dpXknFTj
DQvxB3Tu9O/n8b0gt6ytEqG5Nioh+7v+z+N7rpNltBY1R8jqDfEhhZsONTYL0cCSykTJKEMetOqw
KfkxtEsS+W031MqXoH4H+kO/eGSWrsgrASwhxCOU9tx27siWuk9uWauq5YWUfUZzIb0IHTDZ61O4
qsMKDGX05sOuaoNEdVLwdUMA4SR96CG5a/3nTHxRKGXCwUtu1tvoHS8fN2Aoa2oCYu76peXqTJKz
m7pJoTe56PR00Me7EU1CBHGqKb4yRlgayLPPegtpuS6KPsr6TVz3aG0e2/B629a60iUBIa5B2YbK
RH5VvfejzdbQSci3WhMqytQ37VBce6ZUyH4Cr3ag4Ac6wX0Ru0PBc+RA+RmmXRYle3xwmvNd3vLF
WTfcrIeAwgIUeUE1a5XS+U5/+FGGvXR0X4OA+XeQ9hBhWzS+FR8QRfks3Khs2luRluAIV3PAw++L
FFXutXgTyPXCdbaTjV5fKskgjmvFFHODJ0vpTWfoCA13fXc9ua+mgnorOn72bykO7zdDJGQb2tDK
DdMm0ffb7BMouIwgEmeYNPgtg3pY2p6X3FJy7kolb8SIxDGAtrSwJ6aaJdu1kDWYcry2HGnsyAA6
GtLSb3qIkbbljZluDkJJ1QCTBAEvhzQL4V/R+tqQhdQg9DEUvdAcd8oS5YqXIJcK1iSpqI7Tng7b
sr800S+HoWeDUcqU3faVrCDdJFqrK7YJN7w0p1etWymogdEvJoKtyV1g18d95rMpe05cHFfPrjZY
GqZ/fKaD/mTtLDVkPgMIh4L9zx9bjHyKMqoXCF/QfPJQ8WzON6tdMmmJatPJFH+tssrzNe5fDpqV
f4ou4ch39pWoCaZOig9gLPL6jrrNpg9ADcaYzamMIHpatoyGCbjwslnNmTNx+hADGuwAtHwmElzh
0DjIWYlUWRf0B5eJtwQlN/12Hjr34fCN0s09EqakJ3BRTf+LR4SsPFbarkQlsmhg0YwxT6hDQ4qC
BtY2+F/t+coYe8xhaKJKwIwOexMATgdYosk6Xekko43rtRRP0ymVBX/CrNJv7/6Oez9Vfp5NOTAa
OvVwi4HipxZgJrvBBG3K0SHDS2CHloxgGyl9XYU7hsEverxTKcD+CHcKY8iBqkctfrduNbkilx+T
R+I3UPtFM+F1XuqGrYkvByiutBplNeyOKnZ+4J5vGFzBFlmnBXcM0jxOgpV2c7l7Jfrm0CGhy/IQ
xhEiuXb/UMYUBwrTWQ3OqOFcP8ovYGx8b+HU5QVaWAcTZTFhkaH+39iZBvB3Ujin54gZyjZcxB21
cU/lKpULqv8e5GkcU995u+V7VBrFm3hvnzvEKVRfXQ9dJTCnajEplPQ9jWkf0js86UcaiYulvQ/5
HF29vAdBGwTBJRVa7OCtjItiBmc6qclgcEV16vPZIwJedf1CxSKmY9kPdwwbZSRh2gXz8dWEQ0QC
4oUdwvSGloadAF/ECi15UQ3LZSQfboMXBtF3L8vb3AC2ik5LaLvDSNJdJ9DQsNDvskN6ZOSQPnZc
AH9l0vfZca6G/QNktly5Q8HJTQB29Q4EFM1QZLUfVLuRDH4DFQeB0L4yq4yeRHHfLZ7w7F6WVx7C
IjQ38vdQ10Wn/FhMPFPgJ2zeu+I7qVuJ6l+GYKqgcePTuToX/iG/tujYcrvYMraHsMDnIuob/eYo
UyBKY0Tv+9TBgfOeN7qH6d32PfaKz8x16pPUqhMyCWJyKdM2cBg/CExYrteY6yJtY3RlHpXkFHzB
Aq1OoOkTIFM2BqZIrQkMTrqTbMExJVRbZqSrsQNGaC9DfRx/LvUq6FV13RvXkFSZFSHINHXAfq5q
NwEXSq9T+5hhDSlxn5TYDrTfxmJxQnMFsiL4ZLVR/1ZIxkHCvwmMAqCaM6fUqM7nXQ/j8lwOipId
zmSNY5SFfY05I/3245qg7uY13IUzhs1FvYzagFdR8Sl9/MItnIGynFejhiO5haCgFhcoREzfdkil
ibzqrhgx+E4twrTcF10OI8TRVuTJC79uujD4E4WePSsMoLyF639sHQuKkEeSmbtj/dsexJZ95xya
58lELkdx0ac99WatQockY/FQBkYnftzZk3irrN71BVP3COPnl4SGQP0gbipUkIiMPt19UE+LmAP0
G6ZTNEwPrlvBKhnpgknf40pYxCV0SoDibvkpI4q1uGoROf9DD3a71okvX93PRC+fyIXcanbGCknT
iEJJc6bu3zLytsdEubzMGw/XvJH/9KPPMstNxszBckxPEZ7e7MrxY0taGMcNXS+tAK17CAyLpI5g
wEEIvr13WwOFSMz+8agejQQIoEJFCQ5xLKHgRYiHRSYl+wrnvNWpqccFqwyYHuPIdmPfEhbS1MvR
z0Zc3aTW6uFfWAHbiHX1oY8BAQ+prserWtq1d74eONysRb+xD3qvQqmNhzcqW/337wx2NblTVfRG
iqd300TSSS8nWAj1pxRIzgFuTcvBHfeFALP5MjhzjMooeGGjJtp5KEDfzuAM8pTZctAfgaXtvIdz
LXkKQc9uB/zA4LGwW4VEHaSVcG1/Dk9YmE6CjM221NlRxHL3ccOKr/mR2PxwJ+vC9tEiKUAb3q6j
LCjHcw8QAWYp7XqLhaxNgsALPYnj4zIFSWGbSsLkFRuEtITYSdvwss+4fcz03phRZ9kX70hgXP78
pZPUQx7+sqcfrrvO/TT+Y1V/Pw2E9MoGqfPC+z6+n0h8V9mQeI3Uw/VdveuEDIjZQPQrgjyw3lgu
BIZLq+j6AooC3mUmmzSOkzBWy+hSwKINzV56jb+r54Op8Dh6H21/uvqC+UeoUitEsEVmGrdkEKmP
hOeIcIg3LaI1k1ObP3TdXbOUyy/2uVPfY2wv3ZESQx9pnqpgAls17lUwoYjkQiLPJwBd3HiH8c/1
Osh+Lcs5iFT0Qu+eBCVOoQZU4WC/DgpF5V6uQRWznf2hyG6snvh2Iaj87X8VocrhX85hhALJCOi5
eR/LjFFC++kSjwMNyfpuWArFmuD7RKdkWcTZ6Ysl+PQaN2n4FhAtBiykWOliGvBr6GL2Waof7+Ln
5N5Kduf8PCNACd9a7jrZu13fT7j72zHhzDI33gdMOIBG37kcG/Q2B42mqMKTK/P4GlGxlv3CpVoL
H0zxu+qlfG8oEGytzIEwr6qkhFpsA2kJgTL2FiIqXtuknIkDvHvCPRcgDQfEkxeTFAcONfz+C+0E
lWA3NEnwkbGZS2qgOc0BIgfpIk4QeacOL0YdGcYLhIufEbtUL5PPyQCprroyYQP/7T8Tekpfl9DG
sG53fP7+tpgj2vqTxMyFhPgXs3+Px3PYR9QZRrabJ/82hj7sbVCRVx6f6M74LD0RmSNATitHpAkn
EfCjvxbHVf2v36jmdB72OI3ZNeFMZUWr4hUoEXynR8vm7ybhIFNdq8OJTXo33v0oI92GGHyCCcM3
SGRl2tV8Ue/qNsOy0XR2GaF+72X7FT1jx39S5O82IyFOIWJSfP1L1YF0QzR1fhC0LCE1vjVBL8NH
6Fe2+SXYXdKHUnBI59cAeLXkkqkRYIoq7CMH722b9AkopZUtFMFL1IL52F8fI2ps+1O39jKndUCz
4dNgmyguaJpHZQP/RSpomwHiaZNgVTWdu0hmldKLqS+S4GJdApGX9vPxVu++YL+zhgF/0g+a7W52
IYrb2Ba9wDZorF/SDCdY0tbXngvoKmw1Z0elWObpagFitb+ILHzgaJEOSsHoVoobsRqg7JiBXBjE
jYGBQNfP8VrUBHdy5p+LH59eNgQ9hNcNPGIrnOC5xxWlR4yPoR379kYj2YjDivYFDb25yFALciqX
wM/3EijzrEV4/uzlDpHvfJeljCowkvFBI3kHfan5vUvMWARs6mX/Ip1eDqGhbPMSo+cggUFKyKx0
gj03674X+A3Nv27pAmT4eux8vcHuo1y7LABBdYzlrjul1WtaxVhVFMkhCkrlINk41cRBDbXh4Ac2
LkJSM/Ei6YAAE1oVBgFqhwpNNZIKdqsyL6/PdvX53htoyPA9P2heAJYf6vAUJiHEf0dBWkEXxBPA
u4Xow6K68EbV0Qd+LNSG8jjuM7kmHvX18rnKGFWB2xhJJIsSMzmd+imYalHRqSLojqBfFOqc5gmj
JvPiDvLfRUedIoGUuocvZJuor8ypLE888KCPzN69ni95AgGhy9HOZKJ04A4YQrh89sNELmxVKQLb
gE3E5Wc+kjwPm42K7G8LZ0Ya9HDvFuArMR1ACxvWQANd9SrCoDlYOozmS5UV9iNncS66n0+4FqKx
OccSAz8qcV5L3FxeMgvU3za3JY56t3nNfd0uFYNh3LX2F/UWwqb2rNxVRNrQSEhGO4EUcYrIs8dg
6E9eQoUyGPDbWK1lRM/5nZg7XNy5F5gpF2JOUd35Tr1ihMDluJjMdrQMNN2jc/+G7lbkNf/QlEN+
p9uRf+e/I4+AnX1nL/Paw3kixVT6mCoHHM73pJgJafN6h3RHek4VM/0UCt1bryEG/P9ZbQQYXQ1t
/pX+/lodUF9KBrRD0NNRDA6Lal2pTHEIqNVeyFO0OWTr/JQ2szac2cLonm45yCM1u1FIqu3oZcIb
LJjt3u2xORSYEvXgGEbZVTjrKfpPTyuFRavi5jnb8TA23P9IzctF0rdx+8Dyh/I11z+7OHcavmby
6X0Z26Q91BrYPpDbHMrP5Ibvb/UwT0G6NNcOE/6IJ0uhmf4YdS26xp9QawUK1ZeO1NeSBGdgHqXj
c7SRUATMVZKBSSZ/LKRPAkgujH323OEicZeliF4btV7uS61TioZIx2D763ufAkWt2ZH1GAltPFov
DiYcFMPBBQUe7GgVF45NkMObF/NqbOBMa0wv5Ex23lRkdBa6P3cA6aK0NhyV7GbewGE5pA+48vwn
jPkEw7ZjzScXnjqQFBOa198zyQTNWjSDWMpKemRJpVgYyX8QomMgHmwunaN8pJ5ZcII4AmLx7EME
5K9nnXMUf/YAprswhUbgC3Czez/nsqvFp04VWwRsLByXPZDTCU7emV+Hf54UzvgNdQ6BHz39/ZiV
KgqPkJ3vIGwL5Lb2TFxN0upjfyhjXeyVGSUSiNAcoId3L5VXV/MpJnKoKLr7QvYahrYOL/3oeMSV
UfdLkCF3CrqVO/c6JgtBVHy02a4wXvloH0dnPFelJjOwSyTCYqYa3oVf0oh5rADBHv2xHITqYdct
jmHdypjVnIl3CVxvE9VNkT9wngIBCOmRcVeSmhqc9n5aVJ6dn7/dOZ2sVigUmZlhs3dDPgSQh2/P
gn+jv4jJynX6lYuM8rddNVlrJURhaY1VVHdxtG5+GHGpPajEWKMtBSWlvjss5+SKqCxhxHOpHZpZ
zv027ypfACv5mChQ8+5HR6PTRHLOw2npPUerdWA/NjoPg/hBOX6MgN7uLv+qyKq1Oc3rATtl6Ne6
HawyQdI8VXUtBkvrdaWweP9ysLgvgfxasCKWPUc+cBU4QiD6yzS+y+EfGc75uCOBIt202JoN+UyG
Qwks9CRE9fkH64/cVY8I9FBapJ7I1sveBNkP51wOekEGsx/8ry7Qdnp7OpJoWBvKFRJNs6ooZcXw
pWqHGGPlWPT/iHUrVl8XRP+NlJ2lgqUUm7Nvgpy9cNtngRwWeycf4ADeDmoNEFtCrh6oHCo0s8gQ
3VBp2qLvzXU1APSCqibRgmC9fYhDT3sHjU/oflb6hM0fjLO2M72MnzBTw6fGrbN5TFhlYZdatetR
aGRsr9tqWP/gClSWPuQePBerL+xFXbICk/wknUISRsoVOXIPgMUixJVaR9lYKE2D9YJQRcndszW3
kdD8WSsZPQNGnWXIulCAas56CDvZc8WzVjtQlJqbKlHvtqd+bZ0FzjaRg+CmC9PInxABk4qlOp9y
cX7W3WZRDXMn+rKjhP0easIIPnmltE8JonWtDNtrB83TquPQvbPjLSu5f4+bqo69IVwCSEYe/MB6
p4+68jIfg/8JI0xpa/zmDc3K9XiZ+tdyBUtltS/apnsw9IKmwdJ6u3X1G7E9ktd7F7BCjjpsHkqn
54Qa4fmrfww0AeL3Rn8vFZSbAvZBzRHzJJuiUIe9S3QpjD5kZQZWiaELslMxWWf+tRDA4TLTaLE8
d2FUS5qtOuEHpjouVnIRWwaWDCbYj3TyPD8h2yngbYfQ7IEPr1Bpef7ViQd3MOs+UXDO7OmSeSrk
6L+smHHOGbzOJo5NxushKxgYvYahzbl0Spw/IYJVAtvlAVN29Eph3OVq2BU9kgpRJ6CaGhTAS2gz
iR/DGK44hA2sfLdsRO+RR01t5aiQQrGX8SruIOrJUMC4im/Xek+k1D/9JjTkLpng97EDhVtqtuLA
eK0ZknUt2dG3ZcmfTaQEwgqYcXJkCQOZcgPdJmP3XkFxvOT9iJv174e4+L+htk0SivD9h/1DE2NC
JM5NnHuQGlOCBmweKFKp+YOdLyrqGxcAlZAUD1BIMUfb3tj0lrNwMxyFrlvDyta7m/iGoGgPscSF
c3uhlgT4HyEngsO3foZR/OwHywiXvIyv3MnTpQvQBi5HhgC9Md9zpNmPYsow5aXmXTd79DicwMUy
b3E5+yHuPn5LhkSSdW46GS+MClC4wwOd59ildHQHkNuytk7ctAXmNJ6yMcy+7ufz9hZfmexlwJ4S
Lw1exfqauz+ZBETVwB5W/ceQP5u89x8Rtm42ri+BzXCnUFv+y/kPXI0Zuco5WTItxnMjW1K6Yucj
XtvSUXODykfz81a5Kd+K7DKFICCee2tZjNu9i0UIO/BZuJOKC31gIVY5N4ZC6r154VzHeqqww9ge
8FLhfvDHntgPUf0yyRQ/exFd2PgyZsfMardulQt5r5sxfjmR8T7BZdow7z9Zg8AYSwED9V1fFLXb
V5PtK+L0uODCJhdW4r6sfELLMlkmzo6Tg6nGcUTrHTOXWuALnbezetUmP3sKf54Irx+EHfo/9Lmw
z0ws8b1FR0N0YEB7mTHikZRqVYx+lPqkCElU5oCx130x/AwZFOdmjmERTWYZlHUCnAfYfnhNFbdO
thcAyWMw2kCfcrR/67b9j9HRYp2yg8nfxrAGCLapovUx8w3ChesBrVzPpEuFaAtL2Wy/iEL9EqSu
HZqnZK9aS6ABlalLfohhwUP/2v8kFcAsskRSZwM4Ojar5bDmhcO2bgugTrk4RKld2VUA5WpmMWsW
5RKHRD179P7/W9NX/KlIn5a0bvqdakP98tOn4GKUIQwj8jxCbLmXLjBzDAjivDuP679aOiQY1s+u
mA4FMXLa0XOR3uuMZb7tNmHEfV/gr7bToM9ZglKipv+iRj3AlQHVGbujUYmQVppdgqorFLUdql51
8aAIx1+LBXl7/fiPTAYmCCrKRoaXXTMFzLpIzeZYYgR1J5ucM35fGlQ6giT5yfgDP63uF/FVbaSm
lXfqoWrQWF6y5ngMi1iDcHLStBCK3+BlpKzPLZM05OscrYwzRvl3W0v5SxSZtDaUJKyPSwDBjvN6
3GnXvpg23xhAHFq4QUHaBVTEFT9egqOCdcUlBFTOBYaEliCfM0JUnWnpCCyTv4nfjYrQzxPTexYH
Hml3lDHGvGQ7V0KuoHII8IVLTLvaqft6eyG+2SxejlrMq2fDRrfSkRFFhPs5vu1On8cA728FIcOZ
b3phtKS/7JvKUbI6Fj5ABEMif9LZ7M0OeSQ+RHMTTdD3OLgiQM2zPaPDf/voFcXmR2wRsG+2+e2M
WNvQXUSEj1wJXKUUwL4HAg8z9QMGdVrzibcbQNWaXEPKlbeMkXA03rRqlYGyLqwaa+9dMBAIRnBB
aDrpgvEd7JI57QjsA1L2y3uVtfJCwQFgXwp37yMN2IY1etytzO5xBrjveqf0YEuxvfZY3yvm/vBm
+WxrHsnROe5hoadskMShc4dwnJ7AEFJVHUYzsLhYCiXOJfiux1CojqdCiWtjWxCYcS3UCb37IXkz
5yeyRYrvCNya7oVF5o4QN9bwOuDBx/T43Aqc15i7bD91L7pKh2KFQBy9yKZG2R+DGIM9JC6h3+CS
nfokQHdPb9RKWz2gWXcbmO9stnQrX8bcjNd75JhNvamuaIsGIqbU48MWvvjnM0xfZ3QOuUTEWCqI
h57sucUq8fPsxbYAL7nLj3cVS1hjQqTCIPmkgRvDY4Qlj0K/XhWbG/ZKlS8cBnrGmD6GGNFgdth/
mqA3K4DDN2SXtpwZu/pB59yyqxCtzIxrgINsTsnqMqP3BXrcc9nhYVKN+cn5RZe0fxnO5OvWXGuU
aKp7Ug+EJlgVubNjQp8mTm6fdGArZk65XkGg0pDyjj/DY+r+wq9JoMGFhXef558pADB61YnCwQei
tAN37vC5n7fcuMoYl2Kmksa7Kri4nT9H+LLVpIN7P3U4dMaJtEp58eTCpX1ZR0o9HYD1QZnANNIE
H2azgmAs/H+XxHAT2iqGfWci2u2Sb0m34ac3SdWFHI3JIkPWFwPZeY0/cbe43eJLOXrM9pkzXAwC
KNkp4nQg5gU3cjNwJXOCg49ImYJG6mBOtEmdXvS/rN6zNkUh22uN2VHZtqnd7JpLYjSxsLKRURAz
8mXn64ODbiVjtfPzpNpPyGTQW1tVdevNw3exkj5B+uz2jOmfesuALGEAltuTJ23Shd2ymGbqBcp1
94ck8zdAP5BO9IvzJMc3LJpifE1+irQiM52JQET+oQ6QF35ZcBDFYlFVTikkK/M5mMyWAmgjSzYF
+Id6CF6CYmvY5tZmyepVEvYICNaKiqEFhPNVqjyVbNat4elTygyKZbjVySCjoUytnwCZfDVnTj88
PbsOqaGXZyGKYPbc0+3sOPj2LYn+O+8Vz/A+lrnSt0dd65vinty3XH63oCtgXqvu2yQnDq9RgctV
a6tM8dUrGXk/ahnEkou9p0bGPaQvdj93y0pQPlHfC/H4lmbqz0t9Kxgpq/+O3jhbOHJ86Dr8G1JD
cEZJL69tPk35zAzTKjyO/Dhn4XZoH5xha9QGWquCWalTGXqS8cf/xxXLQd3L3K+1QA6feGnJ/7mv
HADC2ggvIOL8f4RhyJpRkBkNPKLPA67oenIUTdOwCwhQZAkFTkSdZZZNxQsHOzIRpKxBzCNIhNN0
Q83jrljwaYkrWEuVXCVwxHNY9D1MTHuS7dHKyiuyYQxXaGJXPQbpqQaW4vxV5sbZSUznKLh564Ya
0bGHuP5veRo+HOKpciyNHR/RWrr4M1sRp1UdYIdOdMOg34eJA96Vr+/50upvjd6cafTQUbmMXADi
WBWweLKH99ruZANTmm9cxtRfbrOryfZMKk3LLUE/FYspYuHbx72eVXP+8U+1NtBlq/AVWWQG/6oO
Q+sWCmzpJvpGOzGo6V3HPyosWYsZtUbPGsXIV1N1vp+FkzRI8qJeFnAcgzZeaQKEru5Esy35CnnZ
sSV+Hz95iLKTyg7R1d9PnZtJ2putDopUUn8AafuZXBtOGPTiCXs30JWHaXw3iPdHOATh6LLcIJ99
Bb93JEQAZ2GRukDka8d0llZQhoj6SmLkmH16KMo5qIgNooeHF0VE19jjI/bvwsRMRXoRkswHZDQv
8/3238psNXOm5mduApyvryCijOqvXGALSKCKEpAKLQwPCpskRqjEWpHVhdxA/m7c6UwI08SLUOP5
eXm4scamf6l04/HZncqrTzy9aGzlTpIh70ElNRIw3V83ywounbBjNrqh0hcl1sNgfVBt/EXx/zgY
Sm2i+m7EaXgikZ1brM4YViprStN64ZYg028wcnJLba+qGfrEtQWh8JOXzwv3YM+iEsrXxDJzp4U/
26J1xiTHpj7HQaAnLHeT25MeHvo/RGRNxAyrbiKPyf19cMauPufltZVkrE/KaMmQpRM03roOb2jY
ASyw1PmOWqR4Ipldcs6JXXyDqtEzsCJDx7MsfPAZGyOJOCAgqXcJmEoEU1vrO+kguPT718Wvdcny
4p7A/VlxxZgecBDQxmjPtO8IytXNGmDQ6itMcZyVTSsnkmkp3WZZHBKYKcxNhoCoO73A7BrfLW0N
99Rjv5Hk3c4g1064cBm0do8hLWPZ08Ah+xzcoH2Cx0xP26lUTruFEBBKdUZRikAN3kLgGkzW/F/V
mUnx63P+Yun8eKxNlDQHFs3ZqOpeG/A3T0xRxVUFhoCPB0fAUYP4c4PJ/8x4UrNudcdxqsCTnVVi
t3Ahzy22OsMRM8If+XAgTC72cR4b/kC+/bAw9xqPc6RWES9icJSODDxNQdd9XAAdZ6vmJfmw0NGc
JgOVmPKwgZoTCBw+Gaq4lQNczokdGhq6NEJLvXG9XQ5hvJtJ/2JgdMwpA6dUcDXyp+EKhERziRn/
WU9ZcyQJB73AsBzut8fPcAH8VQx8Z/0mUl8qOkrRnPtWOSxFrs6Githnt1cvHv8lc2IXcha8YtT0
gh35cC9buk1No0h5VksFQbom6bJZHEPndaLjQc+GjOgXNoU2BFwuioUyYgTZ9PBpqvFH4rv1cIzd
QDyFQfbilJnnAwnflQPilqjD3GzmgN9YiXluNxZQiM3E8HgJOZKxZR7K4emBhhCvW6m4GDV2/BqC
T+/Mzgs2yih97Sdr2ZuKXoyiqImf+hr0c/HpZq37sJ+aQtH2pydhnD26qcAdccoN+JSuhd7TBLnp
U1OjA8bU4BKJvA+EPZ5WQOOYuMGg7mM30One6jMDqTZRozCabKbWqyxkrscZLdRVHiop5RSGN3kD
890g+bR6iD9IEC1IlkcoPOSgk372rmzm2FSPXCUqWKfWlhyzfjuoQvryzxUpJZXzFHHcfLFjNVcd
HhB3dYX8Y0DYWSDGhxYnDvoYsNg4nPBR/VVYI8zB+uJNflqiWgLfHmcvhg2ZH7MCVgHfdWvUHM27
F402vhD/FuozfbC8vXAUyWeYHic3nAiaPHJ4QAjANFWGJifsAI2xrE8Jsdcz3Lv7zy+be9LSCU0L
Q/0/uUZGVtmuqwTV9v91VsUfcdLJGAhYF9IG/lK/ie8Fg/PZmqGoysoXs6Ml1dZl4NYOU8dk8WwQ
YVx+PveHI25wsLfmyyVxEEjDHt2kmMbaGlGOEdiqvUpGuRInXI1J43R6HR1jWFKNteB5A9KFTWQw
tHEUwaCwTipByMITpT46YZ+gEoIF50RDIZm475vAz5xhO/C8hs3MHwVLqgr4X3/1E3oKrAa3VB5b
1MBdHpc4asAgmSl/lZada2SpAyhqvge2DXTA6IZOrxTBCClK2boW174x9WZcuS5c5jZTrt16Qch3
B7FUHS4XD/2clVmfGC6UP+rfEngYB6lz5NOvOTqJao2SVaiWwKutgiKi39Mqe7mEqQ9lNHFgHvs4
1gOf0dhhbOBXuX71L73qH6ii/Ms7pr6MIQcYx6/kuW5ZxsAvPhdcf8sA/Sy4zHFbfaWPFq2pHCeK
+pWLXBlNXL/MG71Ip091pQILwkDDAp1zhlZZ2JRXOWtBFQ5lq7LLEBBWv1NHV1SSQdnedqZd+wZK
umzYZ3uxXs9mlt1Y5KQzTtvyrYdFdMqHuvWWudPn3wcPAcSrM2k5WYlKfYcxhBpZIxA1hM58pxO/
WS0pq0Npt7bsEyF2vZ1N3KSQMyV5yMlSUo/SQOiVTyCA/CO3kV2mPllQPHChrtArrYS6AnWECOM0
DxtvEVgG6eTT7IDpdbK75ThwXPbK6cBLnfRvsqARRYOkytFELmTdir6VfPSdTUs4F/yMju5L1aXb
JpG8ldjNIhejkKhSxtuii4DwNd19u0AnTbB3gng7Fd8kfs5sEPcNfGZE7+wNch2ljcGcClNvRGRP
nUgGelxF+dLePAxrxQ6BDvHvJPyb+ATknUfo5HaRyEDUgMuq11BjIXYXSIql8dyjzAwTLB8dENGV
EisBor9+pFwNOP6EX+pVMkk4ok3AdBmr9bHzRI1FBCHhgMCCYjdlgRIrtbWO9ZtIQ+gVOTVbglhN
ZaLL7jRAdaen/2KFxQxmqehIyfeyz5SfBRS/myJxatRmMmiIJtoKkxsl4WLTutzHeQHH/YJYV2Qm
RgI39gSsqHkuLGMMt49irR+z/KF+PXoZQRmVDCkeWCC7v5c0VTfnran1jA8Q/+h38kZq/xa8MOZL
NStQzTXdDoEN0Gifwxtup3RRPmWugsf36ESHIYCrxH+3PPogzEXgh4m+9T/6jOMCNE99vrTQ4gFh
x617GE40KMXbCHsahpVhiL9mQQMIQA1bbNpCTc7dslCH2zQhlBoln4D2emOQMriBTJ5DvRJJ9bAg
Ydcl+5CQ+0PF3qUyFR/BlaZC5ZRl5l3rILXmTPIJypTuDEYjKtX0Gh+Sw2mBoBE0KwT6szsA6ubk
Vc8Yx1BjCVNNQrLdiCd9kVPQXycVxuJ5zTlQ9bElUfC1EtIutEPBPMRvL1zaGxIzOjBAl/bH/hKC
R0F6LDaon0wKzUD7ERV8PjBuyotXFlNokHJbmrWdwHRTDtzddPKyD9wcI+LBKkHqJ16JSorsGN20
3LHAaQl56VyQ0xzBX1Li0LXodDkX9CjdgyMZ9SCTB4P53nYBJjR+i88J3/IlfWbBdGM4B3ZufKod
Vd6HZII+Lg5g6CeHbW9MJ4R3fQc1tRtxlyrGz50gb2hFC3xVoy6fGn2x3YO4uWKhWGQbpqYEN8CK
HHoGebPotKZGIWViEPo+ovhz2NPkp25r1cR38xMdr+TBLNwSDujCQJ1+pmtQnvJZhnQk9IQcBH9d
CWzwpfQIGfQ42lRS7Aa4Pa1p5X8aWFPPPn0Kvpgu6bcaslnrRx/9WWA2/H7xGl11/e2TN2NyzYPF
85BKfIUgw6TuAphl2NN4pfOWpUcI5eRzLN5f5XiSfPAAWF4vpqm94UixJmgtK3YndTSF+HvWwVWS
NCljmKijWKrC7Wma4GFx7uARCtYz122vcoXxP/YzKMe+puOQJiWIo3fvpq9E2RDaMgcchNMjt+VT
F2npJg7A1bIHHGGnku043vCor2WaeAe82Pyy5NbZfRacnbPcGZ7MeZ5v4AzA//6hyg/Z3K8BF1LO
cl12vFtJLOVtF6II0gVWQR8Xem0YtqAvqTod2r+3tS58hEcypQVZXqJJhnU5GTJozP4QiPGGiqrL
XNbdsKWkOPrsc8CTvPm0pLejWjpLXReKwpKhG+V5k+cTq/IWCi4pB2N7/swYGMRHrQ52OC7RTu7o
Sgh8xPT5E6u4YPlPEupz3cQKfY70TnvFjY2spMCqLzMQlS8rW9K9qh6MMxhp4IDRsDPwNsxOk+eo
6caC+wzQM/gIBfDRodQ3x4rl8odqmM6oUY5GLxgnwW72V8eYcpBjZUtBrW3aBHcdcdSad0eI70Dj
zJgKgkLhI01rLsvrIgZ3vvU63ITX8/O4HTDDSUYY0o1JZynsRuUw8w3oCH1gf4kS+aUY4V0UEhv9
FS11VohUGprbplibwh8GlKmfHycHw0IfVAETHIrMHFotrlrH7d9z6Vi8AXI5JwodBC2gWUZqtWBI
y1nxZvvCjwfo4euQjHanThdpkqVBHdSsXY9HAlOLsY27Js4JL2lHzYTHtHTl0a6Hn8r8Kw2xxDic
3A6LpsA+zY+Bn3XrxJSOXPgkBjlWOg0Y8Ph4yk4P4wMUlFYDQEmLDZKkBpc/evylQq5q3MqhYUhB
W4bYI+WG2nDuJkMuRZZ4AV2ThijGCM+VLeWVn3/xHzyFoVjsACHAFJPpVbJ/6aIjS0AiwQ0qdpF/
uGWHAHBM8/jRYBHRrDxCRlNt7nQetB/L64ey21Jf+HoE7tGNH4pTB5WyoYcaTKz8eshURLgk7CJA
9I70LamsKbJ0UHw1WU6976WjslohTpDf2b63ibrK8Sq8VjIgh6gmQE7vdrxEhEZDcpOxd4uH9lHB
gorvYFLjEsQ1UjP5lbj8+dkV9KQi04t+oA6Xj9BYPkVlUPeFV90iSOSB47mhUCZ76U6y14U8F3mk
/Q/EsZqrH/fOGbB3cf2s7dchbLynUzF9E/nh+enWfBxoJ4D+dmTtJB1HuR54IdR6dEeH0iCZofvh
SFHzIV9Nb3uT2PJj2OlcGerpSRjXSxhYG6320Aq/H6NWV1ao4E0SrsTdf5Fs2nJtLZ3Gr8QjTp3D
FKyLgJEMCcLjeAS2Hw9SzKJooITQV7MNw3PFdygTpXWK6NtCdVILEaU45B3wPeKfViWGDcNIQH5/
HH58W6ErIJ4FO4kA24dzIALibF62Nj8j1gF3OMjPR4Yb9Y3E2ZR4b4fyXmy2BK5WMeoj65pLbKjo
fp3aUniBdzwHK60BKmncc0VSIle8DIDBBHpgTGBIPOBMMdGnY3QtlqIznJcTU4xMBzwPHBiPMa4B
0FYHIGvWWe0a2RHklcDmeVY2W2pJkD4TpvEp3a8Www0Rn/6PyxuZ1KLlgh9WPYHiKgpsvipKNEfX
2JCwXNkHURXIDfEV3dVkJQXn+0vkckvKWOpXlEW+AeSfdRAQSCX85xJjEzi8trYT0+/E3fG3wfOA
S+RoQRIhW6StpudJfI5FEn3eyZO1t6qrHFnkg4bM9FnacN1zeYcy0eRV/KeBPwJn7T2Nc4+Wxpkr
zxDoj5bp50GKHbalhFBEJH89Xyi/JMELtxrjg/EXUEOUJORHmcE0fVjFs6lkRmrwnUMwHpZ4T/A9
LH+/J0PvmwTlX1NwKr3Hp4LJ7auvSdnUJg51jCdUFAGj1Eu0kUCwMgs+mhP/Rj9gKewY11mp4K+1
J6HeZSuTQ3ckM9iant2EHSb6dkOyf0/fW37xoU5n+9IV4+KJzYQ3w/9jnWd7rfFlh249u9WL4uUY
3RVVaaNk1NLMXtcA6qtrtNneliHX1W37tnAoRjbLwYFg6MykkWItsm+NHJf24b88+cFt0S6iwCsW
eBFamAnHAFWAT9qN7/1hnNsrOTVfv2q8BhwbYkeAp/0OyVP+6JHueX/UODjnAfOfk0fCo+AiO4py
0ZXeLiiAkchkISv5RXT8F+YiH2YVBeg8ZOcEUiOpfiuEiPKV+zu/lJhZ3U/CferLRGz8dBqgD5or
17mis/on+TYICNlawz4K2HQZHVvkBXLnikDwUQCPZhvHeY6l7Lnp6xwJoXYTtD3eNlYnLsThesNP
l5xae/7UaNFMG8mBu1Ac3tAx3Mq+n/nM6LDTlKWXxbFoV/ShNMSpICdQcqd/Pl+cH0xREh9ndh+P
vvEi83vQ/n2rNQ4GEInsz4n6YDPyduBM7Hm+dGIlOgDtPbCX86aGMfWLMFDcIo9FtRBFuCgf/trW
cBY4FMqzAfX5aWNGh/JeQ61epYQnmXE4dJLoCc8qN2ONc8JzlsTgd6ODlcTpjwtkj0LpeRsU2gsB
nLs349q6v/jpTy96WjsKmn83wdCLjXcEWfcqyDbiU4/weH+OChHe9stMPI4yIOMrxMJsb9+nTr5m
gL2tps32i1mjhNUtmJ6lzF9W5l0cu273CbvA/sGL+DOAq5ACiBECBxu4fAN3/f4YT6Gi00LYBwzJ
Zv7n7KDZJVn5Eq8fnVC3xvq4t5TiI44HdOm5qgN8yoZLh3+qudQTcNv5tyJjneVSMU2AF8pW34D7
HVYy9ip/pZFuN4Nyfiph/8M9DCBSkhSkMW0+yq3YTe6jEs9xBTm7aXnusUUJiqt3+6zsngAnSos8
9ErLN9J6e78E8cPsMeXmR7P2Zahs/RDgP8WzVa5T1lpzY2BsavsGyW5vjaflYI1FpxRpy9E5UGsV
MLrQWDH7plYANGirIGugsAMyyRXg+vo0l/2mD+hNYu7DppbJbnzUaGDzVv1YztD7i1INlDRKoA+h
I/c0AYOvwxHjF6/EMMfBHOb6/f+2kv77Tgmy8UHYyc+TXKQt0Y2mBz9C+tnPxCJSufsCfiPhP5DE
KoNwN/bpo1sYzWDO08p4kvMN/yFrcGeFzFEBIS9xqpkGC0B18u7n+XJAZCTdrS2tKuPTK4qgrNQU
KJ6+O2R4YwJQmc5PF7xdBxJvSE3+8hVGkaEvSe9/F3RnV0G3EayOZs3CrlYa8yhZpOdwq/21afqO
pxhCiQGIaQIjMhlb4gY5A5cjVsB1gSaIJGVD0NBN+LeubqrkN7WhErIMAPXPGLEbIk0CyFBpQplJ
11ia9eYniP65o5VNizsaX7VylduM13ctzns+EGIamnytlAEFjsM+Of62TLy7huk9hXRp3yH+k3Xz
Ek9hb2vkaaS9aVbAvAOOrTJgRL/dRVwri6Y4oS83+kSz7ar9CgbL+5EhqR4u8tu12wceseWwhMym
g7K8iKc/xt9f1/qb4TtGvw4FIl7RHE7KWkYlGJdzJtl8JWDK4BPmea19eGYYWOnAbBaHhj/SFW99
HWj8T4+eyK+Woth/8ppjXOGyn38lGmZ4ke7oWaq9+ydo7njVIvfLmY3dhGJqv3ql6sa4w6x4GLYJ
k8CfZRoNeUlOd4n6iwgB0rITrbkLPvFrSZw7fd5izvfSOazX22LeAUeKucX1ZfZQ7TZhqNJZjukz
LBTDpdG7h1vJrOZ1BhpL72POwfosgcuYY6n3gY53p5ewkaBLfrZivwhrIzPqEEOH/cuWSdJgyKJA
eT+g9nolmRO74IJf/qoVrqMyAqFPJc73zrZ9Ld/mIU1BTbwiV7x0teGZRmqwrHkqitCdfxuuDf4t
pMTymNvkyz7foXYUdM+mSQs7KbRUjhHnGuohdsJGCes72eKTWPFIvFYVhcypwrGcHUM2iqaqgqIp
tGfxOia8CDJcVu+jp/xsOA9xTji8GGXu4L6f4ZljSHg4B499DODkMyI6OUmB6L+dkNr1xhhE2TJI
A5JPAyb3JHyAWILPQMzFDqkqlrkyrvFCA206zd5ctseUur22eMQk4Bv9644Hn6hohZNukMKTLJCU
4CS7QCvu5MjJDGNgCHX4I8d0HnJgpIk9BHrEnkBraHzd7UdOepZqXeoPYYQF5J9r0dfs3pN4V+P5
GiKOTedQYfH4MWhminkvh/9thLWpc/fZJ64dfLkwInaOrLuxVfCaSajMnnDLo8o3U9wiEoprVhgh
3YJ34xlqunpJzw+l/yxbS7cEXTKv60i9hfoxLhgtHMqj28ct9pTuagoniDeq9kDuJDncsIrTisF5
ftvDbRiYPxg5eKAcYWTqm4X62X1kBdH7NU+HPF9ZEmbSFRfFxkLLeDTaGW7O1u7f1Cdknq0PzDON
sUT6MikKd9OcAXFysDPGN01b9nM2//H4TEmwyJTYv6lIe6V7Mt3jII7LJke+XDUxbjsdwZW77GjH
UiBXdGMyFegbcIsltkqtek2F86OAb+RPiJKgd33EURCSF72kTq+STtC5VmQxr3blqzqUj7Sd7wre
u7jmvhFMvhUj3/FZw0E2rXpnQUfCMfXSH9wTeBxBk30JqVId9xjhviGwEvXU8F+aH2gQunkSs/Ty
YtbErJyqRme/oL/dkUnR1GNtgJnmt9al3QbKUDWMFz5nDkgsAazUUU6J9eRGedt7d5GzK8yydMQv
NkuIPb0iHv3FBsa7oNO8XmLYejBFAntZFhB2rx4Zdwn0MqLwVbB9sZ+epB+QdIQGM3hcfwnxkNfE
39MjtkF0WA26HqLw+sBfFC+S8nHCsNb6L+PE9oLC0HX7uyGMn0Lbd8NCS4opNSm8hLvO9V3QQSlP
n/ybsRco5nfV+w0hzPYHA7ks0waCrHK/t2Y4//MNtjZhBsUgF4RHprXN53+psGcTNJCz47hgGU8A
g82U9auAOW4DS/IKt5jFCH3JCEfG8wQrWC8IAGxBu7UZX1HkDpvjNcx65Aoo4xAyBB2HZ09DO/iE
sRScBHAOeL7MMdyq87sv5yGKBNAdJn4luHBGmn1sUUeUyJ2gWWgGElAMIq0rVGafmCe+wwNDcBH9
R7GaiL1/6KL/iEnndLdV8bHBEgeJ92pt30o3ATPfTmtjg/lrZivrZGgLSQfFoipqT20fhml1JPDE
kW/D937NASgPeC77P1I+Ccd6V2ZNi2RsEibW+T4j46cymdEvh+fB2eJmrim1tu7DI4HIr9M3/xgI
PnvrTvUHtyEF8JpUyzxFpvAAEgwC3JAtoUoacWE82GsIbDS+BWm92I7lrSSGTzE13IgJx2mZ+Poa
o8I/t7y+R6h1gmpO3GJRkU0LdCL/6uvb0m6tuxERMJ8wKZc/E8fBbaagvliJrVRG4/98Sc88R1mm
aEQewcfFIbq9wd305iMr1CiW0LYiLJ+uFbbuSI73PyNmwgL5kHFyD93o/lYdkZJvdSfQVrZ6Nn3V
N2tqH37SSR6P67ZNWpWPg7S05jlC+GJwCWp8ZugWqbGK4q2IF07mD2HigTL2i+YRDPiByByWvcK7
eiJN7bysR4QxbkJuYFXG6xxjUWrtpWH6oQxyM8fX8AG//VkBIMR/H7EsI8WDKUPJMw7iVR6sVT4X
6kXkuSEJTqi1oOqKNMjdo5Y34M8+TH3itRkHXQ9wyOGFcFgCbkpri0yJqWlMFqmcXZkSTtI+XvOF
PaX09Ebhdrd34Ld0NR9aZ1ZVchrD5LB9l6b/ntQj/rnOYLdpJN8og4gIAPHnCWiQ1wE/KWgY/np3
swBlxmTAUS6hIsEwkAWNeZopwBeVFWk8OknkUY7h9WSXP0qyb+DwF8pOEyRKihMO3uLIw6qe4ty6
AEly0wumzNcRrrYjV2mnFRHxeOnPcbqzjE1jHplCXZ1A6SjvxBOntRo8+SQql3I2EPff7MTWjLoH
/reYVG2VC6l2gQI3pAQCayRrQOJo8HmuoPNPBSI//HR+yhMdrsfFcyBaYj/qrjHmObZYufpg/xsA
nvQR5HGP3jy0r7RwC+5NIl3ZCj4ujvG7r00MWMhPZewoZhNTuT9kYwUz0N4gbvAVmz4Ek4sn6HLg
WaTqMumd2q01yYp3pjYHB0aqZj1MN0ixPxPdaY25QDrAvg1SpDLLuz7+RGBmZi0rNg2Z6JJxpVWi
Z2r5lDCjKW79wKjnAvifhKwGeFTpOayhbTi+G1FcbueVPKR2NPJi1XgS7w5EQ5pm1yzRGKIXzTcX
13xFevNxPd15j2b85aAWRXQTWuymZFP+HYzfRGBecJyQJHwWt/BBmRvsf2gAou8C1ZDFEprte7HJ
UO+MkdI8qIilbem8sa1I/EMZwrf+BNqECCZHu+OyIFvhTuow9FZoE85n9gUZLHsAlkPk79DfbWoG
YyEYDasjOuEIBbpKSVNmkKuSkzn/RttB4UiQJ34+8wpwEAPujwHtitlG0xWN+su8uNsx+e40I4Cx
zUovYrBx4UktdYXR/lltex9HSY2N5T/4w5G7/l25X8iA7/hlewmvxRU3ut1Gmvcg6Nq9K5JBjriW
ei12Rln7Y3D/h1qS595ZI3cYPOhF6+UPKdJEEAnP0JZp1Rv9mQTjEkX3f99iD5zlFXjQNMon7elB
ryrZBUkv6pUvNiPu7r7NHFZgQ2RysyuA93g67bjnsNtyrlSbTZd13atIuZXiCt5+dQ4ZVzXgvJ9q
AoKu9afpnOXHWuPZrij7/PEel1IS6q89z5iGqCJecX8+7VCduwMaGjwawipc1I53/cYP9gm3KOos
O/DsfA/P26+PHBlatRqVFCE6KGupJXDGgcGWPjeJKgc9ttU0IdZ2RDuIftt9LvveAG5VbaKmoOT9
POHUXUOhu0DyXQewdS82sji2or/+0AXUDyVoWDj3pY6CcksbiFxJoD4aQLceKerJPhBt2rgcY+lw
uPSuV3syOk+22mHjcyb0upx5hhQ6I1AG4CgnCPqLOucSaAjZly6Deqhiibsa/cQS6tS0P9BJ/IxK
aQjpV8Rek24Df4PvUKW/LAGUsMHmDdNUyTrQSBm18EK+nNQl4XGh5LKJat0eDGxMIgUvXVB//bhV
FQdXSo5L140QaqsR9PD2fhU4KfZX7elfn22bjVmTtlOjtrNvBosvPV9S42FzukrrDInlv2MuHp2I
F5srrlunXtRXnKAQ93tb04Y1QPWg6ERM7W/57XEDkfhYlcaLsx1Ga4gO7nzVnkL0lUkjKPLJFoEA
DcZrC7Jqbldp8VYCsvNq4eGnrI/LtRMpRttFG8sUZiGuVHE8aiuSkeQiaFxp1a8rHzyiLjR4HzCS
yx2SCE/SckSk/8u/gXeNqAb5fhh7jpIBTc6oyss24V3yCzqFu66OZA95/QmtVlpnDiJl9SopXoOZ
zyaJAjkxu2SNaRI9r5xXZTCe1HY6SAkteRfNgWflPQFffosLFtidJkTm7P1DX6yJR1BGkG+vLdEe
yHYmV15a2FW2nZA0Nwe4tee89vpBnuAu9uOZjCWd2yuEoe+OYQEvx38kTfN+JT2VaXHuphmyByU3
4WIrOIbp7LdKrHXlRQy5FE5PUzOPHqkTWnaBxpFSzA9P5dCfctkw02ccCb1yDCmT9DksK2HgmDf+
PIrFEXXM1UcUR5ArqWMyFCHv2ijN82lS/a9ZF/96GefPPfgY700Oj2Q3h8EbexiLSeyGfcWoRy2l
RcA8WmYGo+llzl7bSnq19s1FcsXfWYWTIoxwS/DQoVCQ3ztz10vpIvVX+S8Yx2M3e/zLjaXg32Aj
zM7EYb94MKUpqqjZrK8YI71Htx4Sp4jppVnjp5PzgF1SRl804CTOM7GrOL11BtFf6s7K2wU5jv+C
P945pPeYDf0Gaghf9A9T9iFcP5ri1Y7J+lE3FLJGaxvq9phHe/8n8iAbrp7xiEkGMEskR2iR3+fm
ABBacJ3PEy3yK0U3j+ANqC8gdVkBBC2t4E0ocRlCQjg8eQG2UT88zZUiRiUdbMgHYdcF47Lfd/y9
5+15Y3vOOO78MU0Fp+ZnO2g3kI/dmqCIlqGmFZshD0detk5VrI3CxAewDaBT7FGzst+4WmcLJ/Le
xLl1dtJecAgErYYlS5Z4UNrPpzVfAsQUSRee+FLJqbvN9mljljo2nswOQKp9QkEHOSdFrrbDO5UU
8bjtDmixb3rRwEsNzhapq/KETqd5AUT9g54ZEQxRBq5AOokdzaG5eaeCfaF+yya/BvxlQJiv+7hd
I2607uG6BKsdV1CHptJIAp6T9b1J3BieAvIcF2c//b0JLFCCFMiWN3s/HB6pXdvK4J5NsIpN2Bgh
cbn50kccvzKRSaLFjb+qegSR9bgxK9OdWF8TRw1K3aHI/H4+It/dMsOezU6HhF4ahNTtLvVY44qC
7P+3lKDWqrma2nXLUgWH3gE4VRAlJ0n4t8sMgInuO/am+1amryNPDyvgTfH5VaYIK8tdzAog5eov
j6wuYWqYRjyFuLsgmHPOItLo0nuMBtgymrESss9Z7HC354dE6tqxfBOISzbad96XU0ZDQMtp3NfA
5G4i9N6GjpGp/vn2ZHR0YFx1VU1i/MyYikuSa3prsMVkIRel/staueSYkK5Whh9Oi3SqPQ5nXila
t7ZkEv1v10+X3K0hcldxTs8A0k/FL6vhpYaTW8uWkAmds/KUoNxeUl1TFyvp5E7KbodFho9bLBGI
hdJ7ZYs9lk+X1+tixLRVWWa9SKU57DoE27k6tNOi2SwpGch2HS5n9Pe+Rli/LDGE8HCbbYGQPbZH
yT6lx+KfdbjL5ued3YaLLuLEpXOzfduaPTAPLbConnOJ0cN4f6OUfeu1ojDV4SiAplYNg4HArwBK
h2i41gqESwMfTz/oBZ6gKOTvH1zAzw5RmZOxGjZOhIBdxadOmFn5ozAVFCPOicwnzFiSYAHqqR1p
AD1wZPBARjvMjpJQEuvlnhlibYy8KyUBu99P03DAezxXQzJLaVfeI7Jv68W7EwbWZvbmlg2Kq1A1
zwOoZPXraRss1R43vHiJfXjdXgKDYokCpjaRV7W1KuEExCVLB4HOaOifshko1wIXQespY6ym4ueo
gdfu+/nJ8dxiLJnF4nWzuhKNEcORQf7d0b76cD7c6zjTk9Lt71kNupqt7RyhAaLHGMYl9/81p44R
yXVvfac5vN0l64gRRowAnkBpIIMiS6pRsXejMuiZFkA4ySDmr67eMhhz/mf1OGOSctw854z7GVOm
xaiLTt0qMKxsUq/rXZius8QuEZCtShbgmIi/XOMohCogclbKhuh4mWa9kfcq0mHgAA/WQNHLPut0
wrx+daTavfQalMMkt+N+wqSgyYrBCOCoVVgXh7ctbYISgcZpcKjt3YCzcQYXMCsehJ7g0Te0Xq5v
8a9vm5RpLBuNP/myyky8g0cq/1xvXhZmZx4DrUNL+mO4bjSNdp6L8+hWojjB8SLC8+8rIJtVISaP
UOx7Mx2WXzITBeIXQWIv3+Fed/ABqNrSyG6fGXZEsXWQ1TxEZ3tnZSB340wKu+DvEGo/uSO4weCu
FXk50quQlakREWFtKx2U/gJcClfnCc9bCiLAlv7sEIFuJZ/XX9wAMO/wapZZFIcXSgntS8aYbsAA
HjnZwVk6iJ31hdfPCrw56RdN1VV2oK+mxrhbvGd7nnf44bftPmiUliSeETCSHULfj/FR59y3JzZs
/F8z2L6K/amYYSlmBz2fAn6uX2hm44T2X+NoB458/VcZWn8cmQYzUh4WWto217MAih4IKVSMm4nV
cqF5JkuTu1gHzgR0G+WOjU047U2s1yAOismyhD6eWyT0Qc3JELBVpyivycBfu5nikhFWQLoCbX+d
4l48egUoq0Kn1GrHSFlIdbuOQf56rYEXRXfzLYeoUCps+V/wpLK5p8SGyETN43p/JQw4YtreloBr
KSXd/3A7n4TLBaJXcNZSnTR9lrIMoTv8D4VDs6KPsguVuD0P8lEWanRz6eUdSX+VTI9gscl+0U4C
/dZ0Osf0r4aSDVa80jMwe9yi/QJRLyw4L4UTvAm33JT02mJr8S0Mdayb7eJMoi9g3pDnjlauoPE1
TzZzj/HEZXwmSLLkZVP1dOvYwsnZe0Z558fPxUASX4TKCuZpngd5WfsOVZIMNqlJiPy8yxFGqOo+
D7dXGR1Yh7JWOjPdlXRF9vGFg6QvD5ydm042v55NvIm1cn4pBh0GnQU3xAJXgeJIC2uLuYwA7a2g
tt+wvrYNbvL81ELAKxDzqAMOQtxDKpLHc/MWDOECtVjkm+QNVC7MozbY9K9AfqBK4LaP6spS24Br
gRgE+0qbce/KyFRRVXp/fmXoDnd3UKOE2sem38gmpmoXFBdGIr9KWeT+UxVw1RgLjMcsLGPYsQ4H
H/yM+CJ7qNV4aCjK5Dh/XJec4grdshXXmqp4o+k1tuIcnReD3uDQp1aERlFN36uFUfIjlWpPSJXy
TP8rhu4eIITNVVMiKXaS+OjK5+T7fUO9K+0y3Ey/7limrbNiprxVOQYWJ5CBDPrEQH6qpAJ1ntMr
Q7xvAnjOOZn6rXfCEyGQnSRqyWJZhm9q/oePdwNhZmgreJXO8cKGgCTbUUdriFWjxK2GYk1pMFbh
JL5pKIiN5BXd1naDAEEEcebWzR85vebarUGby/878b08XesRKTge5yEGbOymmEC6M3Zrml+u/YLs
ndLOwK3vWlaPkzmyvMb4TOT1ugiPjSAF9ceocPU8LZKxv2R4bahoTde4cdqKfsjIDOm+EgDAvgn5
y0oaUqJu1tHsgIsYr1vZY4IUe8AOvTW3seHLCMtQ/CdJezTGluUNjjYEt0T3o426KyDNWFKYsuA4
kKbp3D1e9In9+thgIhuLVzq/OrqoU066ELeFbWqK9mTuvM7HE3K73D2eiisVKvDz33dbNpz7Fr5H
gsNGrnM8ggB0FAtPmqeFqSSTARxJyhPYxZnpUo59p22TSyMJ84BKjPHvQrXD6AjHvHAMSL7X0VPy
0HZXJgq9ReqoaYdyKmmGOKhlRvoRfE9N8HDHGPyyduL2dYhqxhFK2W8TP6KLcGbIIJC+wIjKZ8wk
okM3uxMTaMNpHmY7rSNe7/vBsiQOVtPBG+Atz4ABUowiBelflzfhlaPVUKrOIeXHLQs48ZtZzSOV
HlMqf04B8UYUtREqSL5ZKNBrye9ugAZQZQ9Hx+40BB7uELE7R3X7dadEhyf7cZECuQpMjkjF6w9E
SvAJClP7CeDwIoilI2OzuFMEuhbgbltruYO4kceDE8wMvs0cqiX5N7u1Kifo9daHkmUt/VNprYvw
NJZbOr5OQZb8OxXwNpwQ7fVCAczNY1Xkvk0u5VzcVA1pq8CHL6DHOsdkqrcy9rpQ6Ep+fSIfLhpV
THWAEJoltZctyoXgbdHBqFkwVALb3aV6IMubyZLmjLY93N0HFsNpSBXRH7XOFlltAPg3IW9slE/8
Yfmu0cDUYpnFoTY0FDVGgyGVVwfdTFu7PE18+BYGs4RJFqVW38S2nCuhaBJWSSKmw4sfvMTLBCxK
1hzfeSmeY3vJHDeGjH6GRZZk8Nv8GyvB1VsnwsSerXLlkxMTKqC/m2IAzpfhuoSVCFGDXkziFudH
x4eF7B5AbDlNxpjlnQa1WlweKSmaVMbLVA4i03YnbSSvPprdng56sF189UrOmuUmUzk0A61qQim6
qPvADCJsu5WwdcWNP3Z3oC1gE1igP2bmzq/kshCsZ8BlPqPCug55ByGbKoQbVPuUyd6f70mmyut3
1lvQ59KbqQT6Awk7fRxf7Ld5xRMo9PQ+tuCPzJARc1WjPrO186IFmtKofL5svXa1OIzB39DxH3UZ
6GhiYOoouT09/OUssskq89F9/+7pziOqPdCgQbtOO+6JH62Cpb8fU+z5JIcXXVAwAbb6PwzlqFis
t7lFY+/vkQBspp6KXw55jkTvQhWV1HMY1cZ4fi3tBtZskPE6R/8Co4V6kE2xUCYiZtZBODOVkvcV
m71JeELG4/rpTrnkWwDfIZX6j86c/uTPjkNLhcC3QRg/zsnvJiuy8i7WD5KkLj9TQwd8CbU+qHgj
7CK3HWPPaIGZPkWUHc85t7iWj2ATJrToayLTGmNHcyh9cPBlWY1EdHjFGS63Cw4ukD40degbyJUo
ZAT6h4KG8jSpltapKhwgxJvFbBa/cUhA63kTAHTx9WVRhU7JfmL69fN63olBNP5Yo9jaMHQIBepa
bAWQcUi84ExmSHgohvVdnoXV4CP65bTZPeHZJVLB+yVpKwYDOM5IYX11Z+94KWkPpUpcwVQLb/5U
RBOxgTZnsYET6r1AWfKwEWHBIzhj67Y899eh53nuE5F1Q+PdafizUxBOz5snZneidhKpld1UTPL6
Vo7RAckN5Hg7UL7+6SFLb9nBwGOm8a9HEZRlIptUDASSlnBGsxOtDTazCXkteUC7ET/9Ykvqwyh/
/6X5ZXI6qsLB5HLImCQaLyv0xgVZqTvt3KQruKnbsQAth2gdUyvqNH67dV/PGcI9QIordSUKcoJq
CkH+FLIA1ukXLxIMOGrfIDMRgM13DOH/+jMM86nIkqtoEk0FIGk3UwGibWnobNX4fSJExEsJyIRJ
xKinIOa0kEfkqk2UcbY0irPJqEU/1QzSFiEbwH//tWC7k6zH+Y2L4vvkkWYF3Z5yZi0+gSQdJ7Hq
OZ8jiHp+IgwRmkPXPXhKhiLrx+jv20UBH4z0P55ZIM71m8+nkGGvyUDMEawo5SOGJTqszggSSCO8
QqYz6MhicCrDFnP0/T1xd0OD+OEPtY1mLlV1DDe9HYE4zoDwNTEkiGi6Rd47zztFVp5qy+fq7y5W
+tSkZNIjUZws2yLM4dT3ytAaoTT8NLEDpARvzjpUNiW2UUPKa8hhifrwCafrmNOAPsz9ZwKOnkLh
jw44XkBOJRNxyzrvWP9n3i99+suTRANcgJgjNujhH/y8i43w0bCbOJsB2LX2hyclGqyrH+mMu3NM
i/YjqOu9neHvr9gc16lPLxmMDjk9kiyCquuk4jx8XcQ2C0SZYepfWynm2eQM5+Qn1PLXalf1eK0Q
pwD1qY8Vz3MrwtbzoB9w6FmD1FLQJ3Qlz5+ngVxV8cXmhF5pAxSiYzkD4qRps04x99x6qlKJf+fH
+6/+R4h9kv+bjYg1Lomy5HCG4m7ut8KLctPvuCS9XSVVVzXwte7kgWm+Lv7Ctsf2fbcMQ2OtO49K
IVK6AJZ+0YFytOphaGE7Q/6OadGxWUDAWRyay10oBRj529nhQ3wGKajLGZBTjWxb+bb9AjZWNgrA
ywCizYAJx8+I0DC1OEGo6w5CsRFtn6rPREm2lITmY5Q4HjUfr1LBHzWlAFEJ0+cJiJpbF/T0DXVu
Nm2/QwNlIXzZHOloDgb67YyCjTO7UPAMcHBQBgynO1+Tjfvl3BnFaxXav7nztaYbwEN6nzNBhKOG
iydeymQeaaGjAggMa9lHtiBOuqBIJlhzFAUo4SB6EryPsdIIiQprGyYBYSs53GkCAAlxiSG+IFNV
DE90x0vzwl8PQ/h59RNr/RWEZ/t2mynMP6TPVC1iIjJObDcjHUbzE+EmKsXGD6GcAV9jxT/trpM6
7pjzf4KB7sOtCKJFbQFwYOVlOVfhnDEd0zFir/+5PlpUYXPUiw0lfcXrgnc3MHUD4pQFdlDNE4kX
OryIYEM6fGC0A2fYSpPVKwK2ld5gvNKXOjoHbBThm9qmV1/xaV5/OGs+OV/fjIgbHzNy34Y3hBJt
XE/185/gySvCDKVPAkN3AJP+OQjyBcjdbgRgo9y9e3bTfHQICxFThjPyJebckpjbeSNSYNAXb+zH
jL8vmuK/VnPYWCEX9GkJwGPKZeCE3qxcD+SIajpqPS974xUHAY4nKB7fLQ2p3/07R7LsLOgU/BA+
ACpoEgR5Vj7fnAgQSVUKkqJ0Qnrs0bxrmAOKu2zILdFEx3wnxRWt4lnbxtiiSYY9Uomw6HjpgcUb
nRcvkF9PAWOdMdCZFAEAZ3JSIbbv90Rielw2FB5COm9WweW0WWTOluC5uBI6U/jSyhD8tbm24Xjq
MCcB9vsltjTLr1nUX0qbQZ3Yc6WYthuJBkViRWzpBIhn/wDQhrCkynP6FpnHiyuJGfUHu+z2t4/9
2iSDMJ2BJMuEI/D8dYpjevaCllnT6dp8Nzp3BZKzmxLWTeFjGuw8E5lZEJocwY/4FklDuANEVw00
k/IJVECZTiXsJ7FF9ZOIWUYeCehxCOsG+mxkayLVLkzkYn/q8U3p4KXXi6hKQlI58HBt4zdMyZIX
k5MvPqDl7PFQoHbg1vVM9WL+qDXoiM5IJwpo2IL/nzPFkH1QdO6zlcz0xu+Av+7o9v0q5kKJ9nw7
WGlPhYA3iN4xM+enc9S0GCBodMbCzNLOENrFsfKVzdU38ZDHJiF88u65TD20Z6Uh1XGKZi0OlGGQ
KS/GL75xPbRLsfXF2Fydk/2ZBfuv3RWTkmWsRBrsU4nSmJilNIRxWjgOAdobBEItcYTLzUyqxXhA
tuZclumT0Im3oRwCF5Rm2CBGZL3DeFEDqQbYXfZ1PYbmxhCWpae2dJY7+C/dDjmk8gOQVvgOgUzm
/N+WKD0VHR1sKFhxet5q+Gb26Wjnl+DTFwlew4ZcUrEMAZX5pNt7DtPJ2+1bPE6Vw8BzLFbfFo+U
l8x/sw4HajidSJ71lBeT3F7zDW7IbF0+TW5dH6xP+tmDeWRTVlOJ5KdYsCn7pv2QhQsfak0V23cn
kZgNcwSWo0wMMjT3h+7VTiFakqhP/uTQZm3i/QZiMs0Kv5N3WHUe2LKIV2hUi9KTbNmj43pxW8PG
NvknuvBu+iIRjEJmko93TEbDupGeEWBRpTdx7+0baoJM9KvWUYo+zDKHWavIxxnfwNqCrOHBcR77
hYsioWrPLj6168Ys1DeGvPuJRXCDSaobaiepMGgkhZUmVpFsnfhjTU5th09t7d7qvkh2lkgvpH/S
U9vcFik+LzEcCf7lijtHoGI0ue+6kr7+jaOxi1cwy1Xhs+RC0pppFS4AwJqRQzyuxPeL/aYdmOC+
s2Z+MO97RljeyETvTEuVNLFV0uqcu2FZNT+ssVi62KJgsD7ox3jsDSWqV51W6KvBFUOz0jHbl0sY
/41bx/XX9JbTTGEKbXS7y0sx/l48Yjqw191v/91x3KZGA3sp8ZB1dbMHe3ad8wJKT5GR2cpAykrc
iqQPrikBoA6ADGndG/77KWEv1xqISaigWGrRG188dAWJAVIw3pFQk5gSC7v4T1C+t+N1Xl/vGqWb
yisWpv0rDdy3medfPTpJM4MxMGpnJdYKDOmV4Cz37R+4/zywYg49NP+vlc0zskUfVNku30xxoUw7
UcG+fHoV71FaVMknUjzl9lbF87GzzfJkgYg2OK8ZFD5wa23DiX3nK+JwPgeP45wwAzWgf/qI3QcH
587WTvl23StHfaXSFImdMrUECK/IDKJJm8gigfHJAbyTu+I/hQlRi/yzi9bK1FWfHfSh6xMPuRvz
p12kuIicsMg15vlRVsKQHT1lVdfN470JRLFWZFcHNrSfMc68d1qUqnSJNnaqhUq9Mwl97nDKtvMy
13UsJUn71CMVmwEM7EnQtNQuiG46bZOvdmPzwgH6EJH47YUVB4c0o0fwtVua1UlZNX7BpcJvyUWb
sA+gmiRKGyEGhyCqwAvo219QEHb5MDhbPgLVztPQ++SxUVsdCuDLFO0Ukkdn5nYMPq7JKKp5kcJb
YAX5Bawvuw+Y4RB+v2BeCm3AR1m+tIBLlG4819R49ao3dP+lqrpqPxk841cxqop6C2fHQR0Bho1G
j3lGjLL/Erl4pq1yYPaRUHDiRJVMukhYdXUjNGvR4fcC1ba56EWxUHWgfI/w7Qac8Jj6HAA+rWND
yX12KRwOQZ2/ucayTtGZGCA6SAIDssrxzDSiyIWe4UUtadDDhwW0liouaV0n8CtJ/FPclcPSvW3p
CsBDRTZvH6bpQc60YUCGlG6DL/QB+YDb4eMCDCCZNQKP+apyHKv3zyo99yW/Ax6X74oG9ECj+Dfz
k719flGbJE/gUsJ4dEchV5FXksSljPlSq5J32/feVzd2EtfQG4nJ1lkJqb7ESFH1S9WX2Ux1CKoA
/Dz5VHnDK/Ua/+2MGJFhnw+hPrpNjtPcZG57zIvXy4eTEeElMXAVaAlgKDMDwg7D46tn7NFL+UtE
EPjtMOo7cutfRccktLRIaqtDrE8N0bKY/hdphBRz95O0sATtwuBd6JEWQsNRGSgTZyjAWd+0RXQW
RHu+Ki9fpKOBMc130NDGi+BqLVvusFBtsKRIGYBvAB8J+fmerM3f6MTMHAoxu6oBhdi42Wb8l30c
WZjXlpZwSLM0b8VpuNQR7J7hU6bDjoPKYWp+PRInOmZ5D4B4UKU3IYO/130zwkNrxPTGBGL0eptN
rEJ9sQiEkhogR2hsa/FYJe7CgB7Txzsd5SFVxffm7anpruiaK7skyWH0ThXKFVeRggH23dgdNft6
oyCDc2GGLelOS8GHAbOz1R9QzEBF98X/eAekIBfI04ndl1FoYUaI/Q10VThLEbIm0Ils8EaNbpyl
f116ZdcUVyWcd0xYvZatvwBjORc9mJDLNrXPn9khmZ0cTnPJBmOijI7l9EMe2tcvjt6DKQYjMNP6
QqTyZgn8d19RrVYmeGbvZy1A3e6F0FYqrDR2uWOOav5UvoDWoKr2cO2mSwRXJDm/qkD8xwidCfkU
y6xqhDsFl5f7BUnuLpDM2ok/eJ+xWrDR0I+WYFClzSigHEU7y5VheU8epMjJ4bxEkTKkFus0ZC5f
LV3lipmo4suPdz3iHPc5vDrV79oRSLmRmsWfy4iDnH4v8xd7S2+3RaDbSW6/pChx0IFZsO8ooBzW
A2SZzKfdwRKh/433uwreSJudldfdDLy5VlIAsVxwA51F6qwzKaExrq+Y0Pbl5MWpv326nEB+zPXC
ag3qYbT0U2QQZmWALulPvxxbQxoYR3OLZL3gXlccoUoRInHcYW2+CdZmyzo6V4qrFOk/jjd1RIng
dkFMqDkJ28b0TzQWnKDzpvzdVRmWrsyTCXEkQLUieiBGPkzuyC1H0exyibUTqdol9rlaIfb4mAqI
0GtiwuqwyT1V8L0cHufF/rP6stlGYASdi5si1TJGqxP1yra4VC2gGx9e7MrUThbmOVDgbT+m1Dez
OP7KOAnbs6+G0Vv6SeJjdUqbnTyptOygw1QI7JDn7xwfJ9t7cwCzflRjOgJHGWzVUiebroi9DS8W
2roZwP9wmz7G4RJLMiO4eQXX9rhRvPWaMsd//8CvsBwtoGEuuUZ/ROMFEV+rlB406su9kvoV1E7n
31ROvUpzLFUNrfvng/ar+GDQgo+7ebRXcbjOpNwJAyem8aY1JBlJTP4L/IBOOeHpnnYBgFcmBEeg
Xec/Te2NJiWJo4UwAt8aEsBW9UoVl2fBvO4a2y8B3VyiSxqv6fyy/56L6+iOHRbWKu8GMpcNiuID
cp39ncmdioR4HtwoB3npyjA5G1lYam5ru2PCk44+6Iw3qKTZsinfH24oapGzoFknOVzbUyLRAEeT
kcqlNsIZBu0BQOtOg5RWtuJ9tsD2Oeo9kAtcNL//L2VWPN/h4mziaR1TkKIfY0aug0ye0IrC71fa
NNbxVYM1El4IuuALDU/dfw9q7hcBap060Mt1hoXdborcM4dhn4EC52ffpF7fL+ZhbX4SB6cBlqVr
JsQixw9sF/vzag3p5AftFaY2OEKQb0CG3/HbWA1dYgNKVti8idBhZeIF9V1273r6gvdqL/dgbkKL
iRJRliuuWMe7+TL6UrcMhl+jdsA6WY/PbXhMduQJwr6p3HhIqmnukoQDf/ayFckwSTaOUmESnCH4
p6OrlVUzZOckietyJSCPe0ZjLYOYplJzY4qQ1TVmqlm5P369C75zMsaWJhAo0xKdIkoiMDG0JVPs
yzp+/f5cVl1ZBFKRVpAGm81VZd0VJQHHe3ibDBVEei+KMgnzb2sXFgkrwUvYt3TsrqTfea6TUpfl
XYhKWoTmKLCd80tVXdH/xq8kPEUw8gTAFcQ29l/5oQEWA37rGUmKBqMWZ1hKgBCB5vqVoKfIDJaT
+Vsx/DExfPQlrp1isFnfTV6RcPsLA6YdjDrB677ncqXN5ncon/SUU88wpXr/TQNCDZZD/VP0Ss5+
Mg1ObTwyvXisF0sZaUKQC8obEtcY1zfa5eAzTFPm0ynzLJVgquzkHmHwyOMt2F42Lrp3RnPnPK6Z
3Q9898QLIP0L9eACK5xywltiXauMvTCRev4Uz3ENHrkFD2TGRpPBeiJVKJDAD8Y7FKA2mF5MK0GL
tLdc93uKe3kkN0fT2VM6P75/NLHchx4PBMSuQd6+odvuLHqq/Vp84323Qfi8ILjldGajdCXD8NQh
JrJOlHMl03H2QedBRF4zDP0csy6DZtsWt5wDLdmJ/r+POwgvK2D3f86+DoRuWqNoINQaOXDZlSz2
bHYwroG/8FzpIVV3muqXVOn3ZsDna2FE2BTyPI8ZOMnK38gWaCGo0SkLG7FesOy0PtsVRUEPtVak
Jg4Lk+EKE632efTljSrZ20jJ5dFXQnYvNUroS1UaXwwRCXy15ctswE/Z7X3vfT1U7HtmqNLM3nkX
mNY3P5158d/zFptN6VLJo+4ObjBKAzGuSPMSLEdQzMA/PI8s+oLb5yhBZpswfpPaQ3vojsjgGEtt
b+gElczGxjVJQwoOLBpR86xwbp986Hac+tIdXAIopLwmS+m/mWdJ16pCBviUIQijtGq9Z89wyV1L
D7oBfbADQPIv+NLwxgrjZHcWPvufiVRC/3+1X2hd+9zd6CFxbpU3Vth+VMPRTzh+lbANCOrrEI5Q
fOCapk4+Jn3l4cSecyVPPBNUp9/phpijX0hCadIFeqifi7cGGcVgVhAeMPGA3FNij7j1OvxeAYVw
XUfi46AQPU+OKDu9DqtR1N/Xm4Gr0SrxnsMdIOxvtttCf5IjfpuWd0SVAIbQKuGyYUy+E6C56HNc
2220+RlXqnlMf5JZb/UQJqMsrwaeaxVja/GYpauHLZO5s+5vfoK3sFKEZakmm2cvLVELFBCuQzFe
WAbBjBfzIdvnCaWs0/fnluYbNWxXIxsbAL3bk8Ql3HC6Tw2TeledN2Q4NIGbC/H4fibz4bxZ5+Wt
3gRqRGDbxhc0Md3neAVE0PDI/cWfY1r2aZPbFuO5McOs7j2j1oFAtMsSB7pxJZ7MfYOhABsPn9PX
P7MOgc1gGC+lKXWx6ydkrFdSyeC2/l+4W9QC07afLxe2tuwNqMMmghvKHGUfEdppWxuwlhR/32bX
EJx4dSrC8xjvP2kuW8ghq/+z1g77kJITaTINZeJeIitpZ6IFG9X5aTLOewyw/SJkia7PKbNM5V8M
ZwfNl0cbQkmRzX0yct2P43aq5F86YzfHz6X01vRM7JLmQp98mxw1MKA+6qmJOd9lUNMNILJMOoC5
89r2VQYDNQ4DSyIH86nTtGstNrrKROKMqpegdpaf4dOSX1O6X9gznfpZsiXyAInCh7jWl2Wq4PfS
Jn/3KkeqpuY57tWsQUIPHYtpLLqzP9IdJmN3VTbPyEV9exslPSVgkOIEYQbBEaP80Y2++w/m4frs
mTb83oAuiit1uCNXey1ussquo/x9Ud7LlFw867b/Z3gjrSRzJCEpmj/eZCQY9UKAbZ1OM7B1leqG
Mb9N2n/oeZmTWEixzvmNodzUgdhy3VnYXaSa1OGYMo5pB7uYxeGRgaDSgMtYH0faq2kaNFOPzMwZ
shgJJL3zGUEzQTRumlScW/Ty3kx3zRZj/A2V20OyGRs6oqhVgSq1sVkNgtm1BMnxs1e6R9c2VixT
cJjHUtBsvhJTdW0+IuhwhgaT4LrxOKm2LR0jz/WG1g0zzct2pBWOzwi7wQyY6yyPdzKPCQihkMO1
dLZQm6FLfn9YWAMFP+00n16IgInQrc/7DZtCZ0iM6JrGt/cQUwYcrZEU8OvdXLrOEux1StydMAr8
ihusPBanbTTc2pDxcawYiF7fec7m+2h791LUXjxFsiKk5AsIqEGNpmUa+e2VQldPDesGGOPQa88y
S3byoNcW2jeNdI+u+udtBFqiU6o9bWok41/oBDR4LCPoBIUC1XycBAq7Gw0n63s5OA2gMlSrfDVd
1PQSVcDF5+RPNh8e7ZGFXODi6ad7QQF7kjr4w46v1K8YHuiOEGet2XXewVzgUFPEEyImXw1UhOcu
S2IHAnDeOfL0/8gheUHzvDCpY3ybJ8BQVvZGRsZCIlUOcXf2sdBwO4M7oA5NJmAzVm/nbIE7munY
aby2TQ6RHF/xIZSTdNeKgls25nqDHFq9EuxTXUDcn+OjvNRpGj0ZafRqDtDsEWHs1onGo8+dJIzk
SVZT+nDZvY0B2swUqR+ro4sa1MzrXtDYsAjDbOHjyQuskONcbx3AfKHWG7keL3+aEfTLcwoNeS82
bbgsSmK42q/QPPCOSU9X82UhsD/cZCfgL828Cf7qihGjbBx1LaJ0tCj+YJSidNwsITNZrJ9hDD/5
oj1YnMW3VOTKPWmXJl9zZNjpBlyqyB5cJot590IqEYnbrXymRKs3CZ7sa1Mr4PC18gOfeIpPeZUb
+syDnmYJLw5bXDmRKXrz2Kc9CCCtt0fEPQcwlAukBiKQjWtIbmWeJpPIkAcoHvmh2/QCZST7J/3d
hvJTY/B3y/+Xb8wt0GeT1FbfMwQKHQ6Pm8MsOfkPVnixZMK3C6f3nRM4uJrXufkGmbcMqxo50hpz
nwi5Vp412EkENAxnVylNMcOzrlhhCQGjqkyJ5oLAu5KXYktKwAFZ6Di0hcXr06ZBMQ3SyO8Djmz+
IpqnHbN3Xj58HmwWA9iOL9c6kd3GnkeUAhOuS/LrFO6vuID8S1HFpmli6JspxhkECs0b4AWoJxcw
FiURwJoiyyLc3F5EsvvQaen/WZzGJGKcOXPUeO91Izmgkphyl+EsYy9+nISZ6Zf5hOHKMxFw6r9R
uU+AGB1f4VCTaWKOAw3aMU1rChysHySG49xTMcoRFuAwzzBTuueuHMFjHho2GDGr98ZpGl9t4XiR
LPdnFWFr8E91SKDhlW5gMG6flJrR+dS+LLUMszzqJfENb3bNMU7hTBFvBKQy2aJLxs1S10K5vHlU
Am7rgdyc9ozulw4jmatJjDBSBJg6hpvEZJBqUYIKM23HI7jiBRrxZ3dG4jShdWNb/IoH4rIxIN6l
Rwo+gZ7GvtzdynlbC2Av2E5Q92Zn5ObD4AyoY0aQRAnUARhbE0hEerQe0V9s4Of8VaXuLEvOvWc2
Zt+gdI8fIVtRFbdu+rq+tR3ZTllXWLUFizn/kxOwoF7XQLQb0hVfsKEcsDHSbzF0QaeCK15mnfe1
4k14/zfDrO5QngeNVWFRCjmUj+rzjVIrmrEAGWlAgvGsJgsCqMXsVOTAqKE07ddMJ4EWgZNB1pb0
73OKa8BNKcqpVMoqHQlUDHCfR20PQcERNO2bGszQqpCAbisuD3bJmkgSh6d2/AuiHyD3S+RGoQMr
FcARl17yPDB+PF0h/iE9sQpRtN1y4ZGadrsEemPrtB5SlaSQylkjbxPhv2lWoNMgXk/VwFERRvrT
p6seb3HN09oPWH9CXvylsLz8ic19kWrTQXMizlL0OiW8XtBZ/bxYXrIOvt/9Qz30mbFfIm1g00UK
jatPW6uq51V4JkOTaBFTn0FFCy1wejS4O5yohOLh7D/okVlP8skNuk+AobQ18uYMdlRMDPfCcOhb
BYFBrTPbOMLSKqagG8rCtJO/nuunXLrRTnit5KLVKPzwGO8FhHlheU4owKOj3yC+LBLgd6+9zwHT
2Yu7hysBtwbb0FdkTk/b57EBvzW8Ll205No4A8rVnx8/hYfMdp09olag8/slR6PW4H7gkKusdI00
sbYm0/fuobGkudZVyXm/t2w5bxPw/OX0cIf/wZLsUG2sY7GzSrRDo2hsebHVNJDQeUD0YmeP6jEy
zhJeN4EQ9LSEXmrKX9sxRoFP0f3uMNNcJn8zcPWNmVADM0fAwxenvi0LWGM4Jm7ghwZ9cgIusrAG
equL75qhOR/6QioPwTGzR68E9aDQvL1ln69oGiVR14CbazPSWYZpL8pfx0dJ/7IXlgAZpbK0MZiD
PtAnjklxB9lY1vChKy3QfTnHH1nltz1dPPukBVPXkxgFSRzMWz4iGhZ4PoJ4J9iN18f4QYCIEjg+
64dmp3hAX6wzhorHZKfx8csw+1Ik+Lc/f7uH00kNPmcP/6olLdI7Btta287zID1VJb0ur0Jm/Yvo
U0rdS/GJ/qZWCSh8rhe0nBQ4ZI+R0WRMRvT3e2Xzf//lg/HoxexrNV1zjPN7TyxlnBV3nj3bDmzn
Gaf6bOVgh5+Min9HKIR5BMCTwV/wb00auLTwxBiYVcNywy82dvqaz2QWMXVnGfOPfNiK3U5Vzeb+
hPXIYi9Rik8HufaP2ZFHoQLcrzI2+RKB/l9w3i5cMICnk25PFgBigKoygR7tFyfu4RdwTm8ey3ni
kY5v3iBDIHT0kGtc658LR61qoCqUot4G+MopYD8ynyy0z9bB76zYkHq6jLOifIg4ZHleGjbwBBhX
TnKnx75w+PDJZtZnBzGPecjGbHqE00DXw6mxD17lC65ib0vRxtYiep1Ycq9O67Bwk37hnxu2Z4f/
gvvvICWFeh9dHSstZ6VYKVKeOnKsDTDLZWlqcsS0AcZmQuwoXHESe5ETJuDf9rYW26CcnShm7E7A
bG5wgoSVsi9ZO5/KD3l4ZHibERXiwY4wVwoaE7ORqA0xW0lS1nB442GvA4wGwjuIYYe/R9kD9npI
Rw3uF3wwcKo89zYAE50dcgqai6Q1qvVsb2UMga144B3VyPEor9evIPNXrnbvX7eRAKmnqrniV0dF
tU+6RUVogFpa/s6Evqov5fugPIsMlFMNhA2bDddbKLfEp7nzWE3TrKRAOGS3gct8CHTrGucLhNDV
uirDNL+xED2tpX5BSr9h2V04hk6A5JL1PYSdH3JN2gqt/a5v4VlkNETlnjr54dDogivkz6gKOoi8
SHTRPRCvAbIKeHkLBCSZLZH/XgmyMKD7GH/WBU6hZbU7/zX0Sirz4FFWe2L0teoqboX95v2JrY0A
BPo1rpyr1U/QQZu3yBdFZrKMhxdIsX3VC9xMr66DCj43PjWrfnuQQPDZ2g6akR5x9t/+Sfji4OZR
2d6j58r/oQYMT3Kj6p0RWNUxhcS/dLM6JzXNv1MYAzCzdudCZkJpfQWssNlWK59S5/DZ0no0v9JC
vuZGWXYEThDg8YddhKUn3c6+GbS9akYJr5oAOZSc26dR1VjOTm408k7RpU4l68V939lFhgnL7ZJb
a5YKko39kzvwEIEzupyY5gbdFYx9AH181W0zCU7+1oiODMAPdqZxQL05lulrLSsronE4ETXeafkc
iKg3TniKLGBcNfqx2UJzhy6T5FTRqAZ3upBihAOERf/FiXUT7JYcY5REzDimMApu0mKVhsF0CePP
qCSvyC7df5lj8dMcJdzigpsOVbxcX9jI2xwYEzy7gXRGjH2RCbZSPC+f0tq/nrX84KdogN4QFKpk
C7kotzsK0gsWnd1F1/W4EMxgk5a0r+wi2gJMlgoA6+sHFuh8vOHJyO7FJlX/8XRBjwoY5+14aiUc
mau01ZhWWZAdy73uv0xr5xqNOAdMCYV5gCM5GmAjftUBkXKbXUPF48sTrjIsGL6+VR8MkmoR3A2E
MrD66iq/nPiZC6KD2/HMC3a+/Cycu2cbUMLJSKcEnPk+UrglBouAva/fzQ9naFR+d1ufI92Fr3XS
eqeCQ7/7cIAi5CHWOzqvjT3B15HliodSsbu+HtNfxU0HPC74hiBqV9tChAme0OL2X3RR4cgO6B9o
SHGJuhvwpkLdUujp0LuVYtHA1bNzGEZIp0pFYjR3eKvDKaCnTV40tmaanWWEdfD/9qi3sztI7Ihp
EuCP/4zfIosZxnOIrq4YU519KrGlFn0Gn8TVprATJ6huB+h++BCDGGXoWMOVr+oEzmtNG19Cjzk6
Ryt2vZdR+aCdvX9/+N0lMvOBm4anYwosQ7QnRWen9Q8qwvMzfxVGTNR6YngEzpUxz5UtyDGOATAh
IPyPzpk2wT2TUoYZWHTyOVryTIgp0pMDIQDnHm3E2l0bsQIP1zILBtXoJH4tCOJcWdg7qTV1csjx
bHiQxd0qrOveL3tu2QBI7+vuK/JKgfSpLz1NGkqDbAlNF3hwijiu7CsUjxcLWGC1JFIrmt/Beuea
Mx9AdVohtE0tj51FvQMJrvQdB7Z7etN807i2CCGTpXsFcoXQ8nfZZMQutk9dkDVVIfDWjCySBaJM
Qcs3a+6NXqChfkNv0nfWUZo+cZYzqI5WCoeecE4wDzvhoVQcTfUlPn/e6SEh08bol1cob1secqZM
k9eWSblQsTjZzWXq1bSuRbnBINPJ4fgVgOpON79GLQo26Xku/XXLUz4eiFJCVNCR6Eo1IgENEWD4
CbVsriqRMIbeMvuxhiKLDIunYJJCCDAabwLsE86231K/o0NkpNB7mUeB6JtvGBLzonV7NKWdyihZ
0O+dGm2MIEBGBvpiMDAv3FexXeh4oQH73/hbwiYfmhxlgesjV0Il7oKkqarGQyel0W6is2QbpACi
TPz8fIjkbfXpEBqzzpLr9qdBthYllFQvA3H8agxERJMzfAeYn4Xrq7jWkPuT6C9Q20usaoPAnttg
WKWrPuGwsSNvTbgcwPA8eSg6kp0pXR8onnEMGWIyGcSJuQpYeUhlCYUu/bSa4V+hUvkEun5QfKrd
4160cDvOjbokiF736wJpvqX0kLEuAKyDnzwDBT1JvMl5Pn7NIkrytnRbnsPAYq8ovl3aTi5C57Av
5GadJxoYB3WzKRY6nXk4xko2RLjQtOnZjiEyYC56yI/5mrwAbfNu6PI1ystTCWnEDQUYGJpbLdmW
TNbmiRsvpo/E3YvdB7rT+SR1JIHJI70qfkPN6HEHSHT+kWdmzNmgih38twMDHf+tArV6tZ79yHTC
7vzKas1c4WcUYV7i7HEFX43rsOF8VdzTN1Wf4scV5uXSLYafi3UrtjwAlNVhcVThZB81Kn4PMZ4M
JjRPAjujwBsvLtqNvyJAZwOM3vS4Ej+RL1zGAqwzmMLsoS9Hd2qxn35M7tnBUcap6/O1SDehxEBE
+lze4uB9tf4oiR5lyLZ0KeE7zhu1LYIL68Zv+FHCZS8uLahO5T8nuDHF3qPpBeA6S5r3NovNaz7L
DTMDpwGLjWMtJ/tXkF5ojtPnUqhxkq3fziRoYx9veksorjRiTZtqM/ZWaiFOvjsyICEBFpIOin0s
4llybs+OC2xrj27Psmj8cpmRI6EUR0an6PUXYmAyOPR+B4P0lh+3hxe0Hgq15KJNLRw2DLxbJEOW
TTBUl8H7/98MzZdf1LbcZDrmn78GAfGPZMKs9BU8t1gj5Dd97Lr/qIDmnQIYbQRbwB3X372INbxa
CF797wktHssgIh52Rk+vFb5H29N+CHw9qdfBWNGejS3WR2coBC57AYsGp6UXlW+I8Qnr5so9615s
58FTKlajCOMerHvW03x97SAQGJUWESEAsJ6icQdzM7SdPNQqZYNXbbbz8WbCyatps3TQHMJiXDVh
Ju/kOvd4soTSqMvTJ5p6YfPSac700ae5MOjAHaf0BOAakWjufZQcWshQqksgTY97m9n8YOTAxSXX
A9CEpc0DMuaRBFYd/reVkiO7ZT/Wv6EAYet+K/7Es9NvoYUeAKrN4Rmy0VVWNYUdnZsPzzoDvYu8
FZE97pGo9u0Mn9WMusj5DDjhOaBoTJKS2Qsku/4Ie2hxXv9cT6Il7jzW+jaek+ZukAER7E/NXfRn
6XT44y3qbwwKXy7Gxjdb842Elh9EX6EJFS4iencscBxZEq9exDxem3jNrYv529qEAaiwS2Z+WGHi
U7JiFlrlRMZqB0btOzZtIsKtR7hSyxC5dJi88xyegV4F0KRHxPzApUQEc3rQfeHx0skcIagVbdao
FK/PTZB7WVdMamJfFWFcf2LUV19pyJsS86IOr+r6/Mp50Ytg91FM8Qa4tHZgq76RNH8WukXuVnI7
yAP7YfGTeUg05ruV16XEAhho2RSGrJpyTUQ0f44peZKftawYioMpVMkFrj5bn/mBzpITk2yCywMF
LNsNiefb5RM53lNPUgP/bqSQMyvA1fbHs1B7VAQXP2y25kyLXfCmAuIc7QJ0uo+cGFf7MBBwvi9V
QpPWYbsSdeXeWoAS8ZF7ZRY2s045I8xRygV1DlU43z6AVTOuudeFJd1q1+v+LW5fq9QqeSA2UPK6
xoVkojyg7kFWakriDcpmuaHRWz1/UUlVcGtPoUzVS6OsW/31Bfc2Gxuppm3M2XVYi6jMHqgAsFgf
cgRKepwEQwFSk3+Ax0RZaSwaL7CV9eT/FgrDYYbfqWhzcJYpK8RsmzvmbUl4xWQ46HkO2JM2rQYJ
EwH9NRHLdfEc+Two+TiQJXUcZWN8we+z1uJNnhkw5QSAMz2nosLB41uoYVqnI93bmkPgA8RmaTqv
/BAMhisiRkcL31NRpe8f7N9YlTe/gUR+6H/492mHw+w/iMHUA5Tbty+LhoU8dsHG+gh+S3VCGwWa
O7ZGLkzv/dhwUhNuJVCbW+WFaL4byEYNNId7fsTzPUYbHaF7+TDoTjZm7HGv/8pL9s0JMgUZ4KeB
+X60zbFXXbzci0LfouyShqIXN/6mxQA7VvxcKcOIG4Rkx1qYe/MD5Sa9FhybWbJR3QXOk1iyM4EL
Vz9smJGwDK08rBYUCPzSqqK9yjK2XQzOmLyU4WVhe7w80pTfL0/Rt/ZEDlpNJYQTTTCRz949Yrrp
pwsxcHRb6mBPtRsP8ZbuIUaYxrh+4iwR/I02cNRwjBI4cT7WgFkZfJtISL0HtkROvl9dv+u02f8N
Cq1w1xpi6TeXvhOrkUBctUJPDupcciPu3+0lY/mwcpH1mpTKDDGOouby9h8oBNAYvgGfcsJpCrBU
GjcgIDpQC+diAhGTgyt5Etmd6QnVrmV7a+TIomBNvxEicVjMIZauRDoknJrhxDyFGBaAwCH8ZMHY
nkNKI3ZU/sPJg2xTAijN2uaPdZYuDGl+3n5rhESAXfVz+baoZphkGFCRQiaxtrYAwgNpOVHg87P6
WN8ywS6HsYKemTkwGMM8tZOzDrDF+WylQYQlmK0B51hJne8wZNAc5HF9fSP6Du58iCJoMuGW50b0
EDAF1Ihlot4aU2AoDhETdHVde9BYDBVZ6rseeizgczPxudrWEalg74Toskr6Rz/u1DhpEJH/uRCn
2PkZjr6v6PIEdkbBv2jzzrDjQfTWu3ok/YpCVWbXpdi0M6gUOhm4atEMW6QsOeHjgzgchJUQiJOf
PPPkcUJaTksXh/KzOe965eY7E3dMxzsAbWgTdtKXWGj0oHNGvd7gzjqiQkaW+uBXK+78JUeHhIlN
95fxSWm0SILojUnRUCkdGUnDlALcD1YxTD1Ygd4wg8r54xy+P4yKyPbj7I1fB5cBEq7qCFrljAcL
Z+HwBHRg9rQMzR8aqg7qYDFyTPORLLW+/toMfCA8oSmKUWdtBUgvMRW2ichmr1RdFakNu0LmX5iW
vk4JUHZH26Y/ttuQqHUsXd3H0aM8oMCVs06PzjS7AqCFBpSzaS/vD9rHq+jQbuZvIk20uGnvrRle
8w169xRUMHvBDDDxjQSfqFA5IRfnaFnxy/MxMmgDx6HcMc+uP0mn99IeesB5dMJFAeWPNuLi3MZt
yGj4QQ+CbyRLZDe6sT8AHZu/KRKwsO8SWpsQlpRP19bakt0EkWDaxv882qKQI8C9ZWUEZguI4ewj
QYVcCa4vaSjdpyrr6UDTBc6itqbwCE9g5MNgAZKzaFNw8kQ93IgTmdOgcxvvldmMsaLdsjiW3Mue
LNOtxJ6cFzLWVgu3ggZg/8p2LGHPcX/C6tnGiezpcit1xKN9Fj4g9JooFAkqlmBYSYcGU3soH12L
RbcwHKHk7c1VBpbFmXgdJwMmXW5bM2wizLvCd7w2Oh0VGWIDdBPIlg3Pu+E2jPmeZVZ1EaVv9nE5
SW5j0cPUmvS2tmm+O3oybCg1Qqyd/QZ8Xpu2pr3JjqH1lM7rbvJDqisvdO8pqEkHEMx8y8OzFJep
RvQHSTQagwl5HoudUKcgh3FgS/6YggC+O5BIVpA6qLu6m1R48hwYVc1n749AxXJNhiEblGSfaAwT
EDdQpWgJW2txS47kfrdHyUoeQfwLEmureB/CPvovAMnA0L8XgAfSDMO/Sv2uSCy0upXHrYDnOxP8
u86hdtwryaKoKNxrwBM7y7dUPu5Sxq9vLPD5XfBvwCL0/nHWaOE+7MIbAnBr+68HbODV/iJsJ32S
P82hzZVAivSgfq2gt6Hdr6rBM53WiRDkwSECW04zIIPH3iSkIKu0OYt7mmZxhSrLelqAKLsZ8Rtf
+LxFh8ROeHUR/d+T90HryqTTFqHYTpVUyf9MvTMS25fFQkEnn6qeeIylAYoNpMMkyX9JKeHIbIHV
4+cYFCoVd851cSz3PAN57jwpvfKT9WDQhOze+vkuKxX22HSkHyD/fKD+lZYJRlPVDLObHB0PLp0e
DX4BEs3AP+GOYPqYYZC8KA6e5T8M95On+T9+iRBqTRuwFuzP+yGw8cZCqUUF/M5Jb7DsEHBTfQoe
ylkaDXb88HlhxFX7aArfWb42j/3tWgXmpUyc6k2f1yaVX3jlBqAVkxi16/n8i+UidFWcwgVIxsVy
FCmTba4KBu/ADgatyqeWrK5WajBDAVUlIsMpQtGxPyBPkuQckDpcC4K/FBYQaXgdJAPBYayZqkMB
fkKniQ2nCPGugoH6OIsAEQx8qJcRYLBtG1vnZeo7KE3k6Mf5LlzdDccA8R5n6yI7bRYDvuHEBqvP
08Et3GMkE2tJCadn1YhB+sDa46HWAdlDIktm+5Kx57wNKXp7EIxbvnDOQv6+bkCDS8I2KFT8v/vA
xsZ63ZCin+jzcgGPUoPYd8DhDH9sJ1xCoJPKX4RUX+JqvTRbbsqhWsigJfD22FPTnSEGvm6Md0Q+
0fJ+/zc1Cm7RkYXHcTIzqUg9B6+LZpoB5tZG3kMYOAQHd88YzKXVlriqau7o5iV9GX0BP0qlIaEW
2eoMtQekiCTxcem5Hc3Ga598w+6u0TpCJhuJVc+3f2h5W74ax6vRDKqbxF7W405BwPJkpqknGSTj
D0rYutvs3CB0H9rS7hxS8SgE1ZyEHB1dfFh34AEGTagINH3rS8FOriCohGgV4Sui3gDwMEZc+YpJ
tDQ1m+yl+lYS0tiU130ozoUSXoLOg8EqlGgtIEAoVAvenl2rwRHCDct7j4F1Km6RbaJjLAzU1h3c
TXaDhcC5mXBB8JiLOtWLCPQ8pGHU1K/wUmLfVwS0VcTbzbJdOx8u8rjOXp38CAV3rfuz1V/necAg
lSJKquaA9zbMAoLA1Rsey/p8Cqz73o12VApt8MybCIj4uzOdJ4pcKg70upHneVdVTsPB05SPyHG8
eZJS4q7vw36Ub2lpqqQ+5KCEBzWjpHpBpA1g+tJTPAmfMqaqqLhXwKbImsbg+I4nE5Uapd+0PVel
uL9r/nyzkHDs5dL0rntBSzmyzC4D8XLwA3jZoNiCb8iILdcWjek25e5zRqQjwnw+Aum5ZnnPRNO7
CZIiVYfs6vJOZPwGAmhLI7nQgnd4ZnBF9iaB4d8sVe0/2fjzMJ7aMGD2qohPFTrnjD9Ia1Xomqrj
OCXea7jKPx0RmFdbmRGMoOZ0B0bL4EbYycFoyHXScjjYrikcxGDlLMXJGxBjwURxPGaVFHkbbHKV
j+tJVsZqBNiv2J0TBUr8tt6OSN0yRR5UmCm3bZjh7+NMVcaeD4PkTF+ZiYX4n1B5ZsAMXkrqP5aO
SFSkj3uM8mtf49uk7wybfKz7J2JMIeEj268AkNglxv9mPXJZDizzGtzZbn9qtIngzdFB+dukNMfd
zRxfEiVrFrbtUX8cwjfl5HB3as8a7kfUft7z1HpVauNtjtXfJaqTV1CmXIfixeL+i/TtPE2z96nd
VjF9PjjzOk3cJPStpQvYMMXGIgW8u/RxpYGBToA0XWqVwnT9+ZdLeuAGZbLCB2otAyvECFDzZrVy
E+Md2h9IGq6YABf1e+Q4rqIuTzt3qsspfZVx7WbjYjdq3WIhG0+FPR6iE5dKZfCg0CtKv49UVGnL
JMlk8vxY3TNUF5JulPbj2U4F9ilAi3X94AzYIGgeUYGPVLrx1AJ1v+EHhkmVJx/vWrnaKjb0fAyY
+xc28aanxGIFZ3Ztxk97fvTJ51wdDOP+AsKpSBorZaS7zv/aPrZJL3klpT6eZISWTYpe7Q3wh1Yg
dZqfFhQv9geRhdWAL0Y+mkOileTrpF+C4YIa8ER21bVS5DonnD9m7nm/wdP0V4ROBNK8zx3mFS22
7W6usTofSbaGKIw/guFtaFLnXf+UBbeLx4MAFKetwiw74CYakdgcpFj9NPgom2aZLDsqgx3x8AW9
cYEBGj9U0WtpvATSNqK0vSu/KgLcL+zk4qTtwVHau9NWX9AQYbnr9gVDP739oH67p9B3fcOiPAvJ
awcxsqZ2n30vAxkVF29kWjm4weiiHEpoJtGkpPKg9iRDyaAsitm+tsPzAhvZoe+YFsStZCPJ/f68
6FZ2CkJKVWErQ3F4cCZP+temF+jHVCV0CFeZCNKd8LkZMzzSbaS6OU05vAQUk2cLRBR/73gL5if3
EyKblHxA9+IhLqiXil26+pe+nLd2RvsiV3k1wP9VaFMjXesBP6pp9ul5OzbOz/rRfhaxxSsWcnTR
PwgqAKCGI+Xy/7QBfMp8gNg9fZDPDYAq2m5izVPgudmqcSEkMiSF+8V4mvqCn2CSBxnOtSk+yGPB
XhNprlmtxiECQ7iVqF1Ypr09KZJteyiJOzCa1EOVeIuMBP+CXfCM0G/WFesbD8cFlF26hWQxnTEg
acAgw5cE1VazhP0HAAxGVD/8DbmPLLsBrVh/nvOLf7avmteJ6boiSmDd/weU0YhBYEVeI8glyCJZ
XCAPDwWt1K0M7Eqiaz+ldnKOQulh09deQs4aJkAc2Z8CFh7QBR1GDbikOHavXVRwLJ60fe0Tw6YG
KSge4Ck8PbsQPddZMLTGxtPl2I5UpX3dzPYjkuE3JLOc+ln2mjtv4Mid0iU670YEq0A3ZZfEcQCh
UtzdVj04CFffI+kqSgOena0PxOWU7Kf1ooVuq5R6gxb0zDiqtrCFq3aohG4RnB5ynZCvzOMl1GD4
/LutU8IW15yMqNqStqKw/39bkhVhHC8vx63YODdAKUiowS60rWsSeZkAIwJQf79kYTvuj48B/4Ix
SIKUJWJuNk7gbUp6fQU7eDVItTGt2vlgw47XOzFoEsxXPHkn+KIQzA7OIt+qElv7Yau+dphiZNKF
EQCujHYfB+pVGDIyJr8F/bCKq+jbyFcqeIqdpgi2y/T/pPkYMj7Bn5Yxo18Y065KKwx4vyj9YPNO
J9VXfpMIEiYURpT8T0RjDO3WsbN739GCae9Hrn7qTBVWpNd8LFM+3KbjmDdXhArViUCVxfH2wccI
irzDAgZJ+h++33p3Ew6TLNWQeaztXe2k69eyjTk4aZp6eL3eLFtoMjrqi6pxStN4PzQ/q2Tp5Wa6
Vt9WWl8syxTEhpRkKVnzn48rKWQb9FqJuYssouF/lq5XbVs79/yCyGvvkJld65w9fh5FwoZKO4fF
679xiBVoXwTHIODdbZriM2kb88V/tFmTcNP81iBc3ze+NUEm1NG3blJbO5l8vB8GhL9+TOvF2QeE
ID684NvQikJSKEvsX07zNm5yp55SZrcREm8c7iFx+RvfjwS6wcp1GalfkS1tRhNw4JJdvJUD4Kum
7EG4yHzzKKSTv1znMMN2ctEpWzDdVbLQKseCx2tllHPireI0e3v/upOuBHhS+FO9hoKVoW66SceH
HMt0TrCiukmRMsK1uecmLpLH9pXSFenBW4bp+LA7/Dhn7rx66h9HNF96DsCwwn8VCoKqwA11mvgE
fhnqOD+Aav2loiGJRUoxMVAwa4UJvBPF49dM9Sk5OQzmSlYUGNwgjTW+sNpVm55w3A0W+qE9Hwhe
4+WBV/MuKp170SOMwJO11Pn5mCyzPaYt+TOq2RVlgX2HHipTr8jQNK9/IsFCpw8zZSyWLA0FsvtX
B8xnABiqoyzP8cSkhKjKK/K1tyUTc4Txjo4z+cGLQkMlt9AJZdxyOaPwBsMpmuAwIAHVWoeapJoM
uRwzdIVRQ2YRp9iX0H+3DTr8iwUMyk2s/CQlBBBk0RnEBstsyUwpm5DrFr1qMfmkfIwiEiqO8kzH
XEcS8qO3psPFVjX2JBhuI0DrjNKAvYRk9INIx8WDJoHeeFxlO9XIMKVzpJuFeL+h6V3c/yiG8tLJ
pdnMbDk0DO3VzoJ6EqGri1KsqK0sBWqD4fIBRhiKMbWY51gRp/W6uIP3987LjRAKUuzwNrrk79r6
+6M9mG37EMi8zNuymDOrBaF7d23h6wkZ25RGRe5y+MGhl5hb/CtimVAogyYLMvUEzrO0uwzI4SsE
M/VGFlF43z2kmogPAqQ2gY2U0Zvwddfz3/AMIB5xD2/NPJI9+cxv76kJ5hG6m3BAdoBBEpC6RqSR
xS9wnvKHXA551a7+Btk3TWKqeFSItJPA24UWUnV09/2/bZAGnlz2NDtfNkHoNPHcKnrhDFMVnns6
smBxu3v4aXY3EekASDx6O1FHyDfsfvjcBmb/DwbHY1xZUw4TOo7Zl/HnjhierIDNSt+MxXuMPWeE
TcaqR24sH4pIR+5gmbnbVCOo+pAm56ZXxYUC1cK9u4iSnA8Wih5Yy7gqAMDOh8ykK79rqjr1YM/m
ejoMSW0OGn8/rRsCrcwjg3MrjNtcIkYg4wsLYYVgRE81rdbhnHIne4ECHIJzkCbZcMH61yIqITSI
qjA5MfykBbmJj9CtSF43Cda4S+DBe4N+qfJMaVGS9ykeVwdAd0uRt2BIaF/SoVqGvzi993f3UjeO
Ubi3RNaDbL3nDIxCvn5wisdbDeQUWDolpYpl6rg8jBPMjpeOZaEvHjDbGDufxAXjCf8jV143UpSb
loKTt6vhYBjUDgamITo4F28WRgbUad2OGHzD7+/ZW4Kno4LCVmEBNKE34gxhXyGU3etTK5l6KnVD
dZHjoqhEWwVQyg2QdMsBUoz31hSkhrrlt9a2KJMROLawRkMIQbMtpo/J5JujX8mBhUuncbaOsZoH
UtvHcW72jBnitKPNMJvWHhMGPj0fr9JJ8iMihkMzdnLmIIMBoWDNix0ZofL0B5KznXyzqi1l2457
ZTYKyt4AMUPwDHzNoDbrU1l6XaRa19VWBqUYSTGj5F5bPfvf5TYoaV57TBPUzbioK7+em2++xdLZ
Uf3GQ8rGyRABhEca5go7aDKu9yyeCXgkQ65sBxB+SNZj9XGZAV9/SE6k5xE3ldFdbo9jr5NobTBo
Z1VGpjkHG0Xe6G/bva9ABf8O2IYH/w1naSaeACqElLKAKbrZHXzisjXcs9HgXRBd3fK9aB2FJrmp
mYYia4jeo97tmA7jSeA96hn3x5cvkyF9BwGXy/YpmF0wHDTr4CgDO41e+0Uh5CBS3AcreD1BOl2x
/aqdpLfyI94aC1CpyACKxxa5TKbIxY90GULUMi5y8xcFOB68lU8hwpmvXea2CZZp46UMCBrmvtSh
huG/fsR1uLblsN7qQ667n86lZw37g3yPV3OnoykOQ8hPc90dW888IIWIdI4N128yWqPhMbB+GH+H
NWt9ifJD+xYoLiL3LQfQF618OyLBLJ0sFgKOji704lOioYwc6JH7jayoSdNoA8HNVS2OH2hZCWF5
pF+z3Vtks8PupEyw0mkTde02cN6+kPKpPMHQ8d+9CM345wYLxJCJEG3giXchFhVI8SsoeC6nyjQY
A21SuTQTFowk/beBUK0SgQhhaEMEYTRq4sDLoq5HmSlmZqvG7GUMcbSRy6gIsyvJVEBpadKlc68/
6Vt9DlsU0VozoVnzIYsrm617DKG7wCMqgLuYi49o6SDN5AXx21+Yocz04Dm2NitshxaePBcD552X
1aj08eXN7sm/lLXN9LGDqsT0DDEwPfC7FXfy1iyTBFgX6DjIIAlE7e1yzIMPAeynNLfaxpEoWTi8
sFnbjof0r7cD8ljNytqlhTiiQFl1OV4eZTcmAyn4o1Nq1tO2POTo+aMlZTnS4mnS8kFOPIJLnkoa
aqx58Tn3Q3KDS3lu0c2VBD93i5bBVHqwPogP/OEHrHsmAzzl16Ne/CR1Y9bTeSPZRv5BfxSuN3Rq
NKivWVJOz570tOd6j38MhXase0XZSMicJFNdKsc6QVyunA3aMGKzc2jsdcQjX4dxuJSmkfvWws/A
ZUN47dY11zLwQCoCTANecc7baUnNjIkWtwYQXGgd1gJcOJeNwCya/Hkxc3OASXRhjg0Pu3xMBsna
Q+7/66Lm3xbZ0xXfEQYWEXtNcVAfUBLQEA4xVSS8KKCzirR4//csIo7mxs5LaHyuB4ml0M+BkqyE
ds0QI4zHWn4utz5/XOHS8TnUmNkFLUZRkmIPyrCcYG+jmQOt3C1YA0JCcGO/aLDmnVh8zAFMM4zo
Iqx81ghgoNDY8+LqOC6AT8oeyhjR7ZOekZ2VxzZZNg+Xuw2E25FUYtuQCvqEch/2Mmyn9bQk+yuo
p6zouU/B25EKBZ3JJcuT0w9pAeh/Ri0z0fFmIUI7JRs8//U3iAPQGDdaiAk39dOkCzxR6xYdjR0O
/+JnqWP9qvh5aixBWdfW/jmXBEPpnPvNFeoYRPv9In6MdKLZq6BGFhjBmxI9HCeR39jZh0GC+Eeu
hicCPoPOqYCTTOSqrbTSX6ahIDrzYXQurBQSzlWflnUzsEFS5eNA20CvKJEtrF4Z+e6LSeAkeZRQ
uYMETVaoswqRlzIZcgPamy8Putyz7EnO5croRDpwNM9Lo6L2UygfBD+xOrquo5hegXu9mm44P8jB
LuPn1lRWN8xkrh7nP19VrWuXchvOo398y2IUQrtzei915DV7IUttmxlHtqSqcGMchhBeXV1GTdM+
fQM4nRV6i5tfkimwi6ZyIVhqI7DrrNNGmIrYCdWtMLX/Tl8+FvmZAjSXuN0BIvMviqSrI0P3/HOH
GP8Fc/TO0imx+WrEmxGv2nZPN2ZPUNKj96jquVnp3HM5Mxa7CTOQkFNrZDAlYpalRHLyJUurDXk4
+vrerfkrm4yD/OZF66Ri+aSlOtdWjr9vthezPci1u/kRwo76yrLxszaoRIo3S5Jn5vo64sAk6ICR
RUT9W0DJ2befyByYXVZJNZ0AmVQy0ZMj8mDLFYgFw2n+pL7MMjTG7BI7lmP8ENr40ogSNCrBbVw0
aDXcR1dGbFni8jJExXIqjdcPPHIt5pDSBojGlkHLTHiQ8JXyFW1XkYXXHvRehyFCuewyhzSVMttV
OIhZcD0fLeN0pEDXXgsdt3M7pNIozkGLCpxgq83tkNang8ZL1VZ8ZMtjVKWtIC5yg4GOxq7p9QPd
yTxwcBu436Enu+abSSeFvb84iBq+Iw3L9CYRYoK7tjm/IUU7PacaQ+G/H3BqgNH9tt5tmu8jTv1c
YNYg2JQdyyVawIOzlEhrbF/n0fqm1s2ZSKiuP7IkabCyt5l0wmn7xE8Si0rg4RUOdNVAaI+MX9rh
xNPBXHzbwdZ2z4231dYQSG0AtmPJkfhILo9wmhCuGLgyf+9GmDGhh9ib8ge0viYlA/5BjypDvkyj
4FA8TUKPBXveEq4q/nHrhs6KTOKS+SSJAi3wXWMteUweL/kJuveqiiTco/B8D/5TUtH7Qtp3ljG4
P/V3nSEloeG+fxjXjuM6DOXAdnRQ0roXOeUpXXFVsk/vqmVbQPSq+9kxHN5nmLXyFJPS5xUm+AY7
167lw+W9jkwEfovEGll2kV1o6b56PZILI4swphOJqyQTI6sVAfMoWnOsNrjor6T5IG+LOgrAPUH3
tXOGSlAwjLLF9BNKbCQc8tlu1JX1IXZTY1oL5h/R9cFhwKWZfvONNQIrSX9xntVbPqCxsb9DZqfX
CVsTTqwi40GrXAgO4+1TLC7k/UhwU33sd0yOpdaP7JqxyAkCwg6ijFFNT17oAEVFCNo0udNPxlSb
vfbI+oU0YZBVHxlPhk1yviwKpZ4NLIYDxwW1KhhYrFOzdfnphw8ERQW0yKCXzMsuqaOJXxzBFmhn
C/dIntT6d8eVc81qbF4Xgr3xjRhzJd+S2CdI/cqb6ZLgKjgT5Ki9iD8PjTzYjvZnkATnuB65cLn6
1LCjIvn8JHhW90BEh1K2r2GBEvHVnn3HyIhsR59dLorhKwjO4hrsDR6F+kRAFdGJmUiMkEKwwrwa
cOVqEfclF+oISPeSw5c+hFW4f+rMZbpCGdD/lZ8PXAQgoQcv3m7CjVAU+ERJshwRfAh64U4s4/D0
r2cSYmS0z+B1ggpCOdN0Vq9xs59PHiS8Nng9rjX4XfPvaLAutN/FhgJi4Rw4R9rsmPmU7ti9gJ9D
J8+Ok3RfWTSQgnKSyKbHKidgg5lkPascV+ZEv1XakN6v5lP+F1RKoozfEENPqSoJKncEH4nmNI7V
wfg56pPbv//bV4FHODxyvn4WF1b7OxE9h195awCot85JLiegGmbTyE8Rr0xHghyVJBAEcUpg26Le
R6q/JqBMiEAKpUBXG8vEiH41Dz8dHqXfdNhPFsZUHMQ9QMiGrj+T2mGIWcYtfejkmHiWI1auigKc
4z9cE9soT6Is5XM8JsqdwruhRkG+sJ8Cr/maiRtm/+mxP4utYS3rQgcsAnID5Fl2d5uefJRDl+Tt
XTSpWWiSGJ+2TJCpO2FS31+vPkhNIOQRlz6Cf5v+pUvc5I+Vtqw1CKi9ZF+wSsaGc9Rkij9Qe7O1
EkxTs1ivaZ72oDWeoTELDFAJ8VuXMhGILDc1PpV3kuy0wL8Js7V8NowfchOavd8TOcB0hitaE5eO
nYabb7vdpSgsdiFUQQHjfWH+H+URtv1sfOmfFILzhNRb4aVoaXSXqKsnGa2px/0WzxsXjJmSsYwX
cYFrVHLtODf9Gj1CzVcEbMTlhN60pyouALT5wf27Of0eRV7NjSv288k0VY9K8CbQU3/99jZ7hb2P
+9ZsZhm573HOoiNk2UfXSAZ4aq23FX+LdW4dvHvJPiMMMUrxVEZSJD5XqVvOvVVgN9GrvM5xQm30
LDeJimdo3ecTohLsarfotvawv4pCFTGkiIisqR5PJukIT9pXWkzh8ewU4Re0qke4dnSXMFcRRxMp
qiAhxmTtHR0ZaHquKgzjjtkU/ueGgMMBufBPoM/c5zZ1ZcWxWvGpVZ1N+9IRiHxvmOcSDQxQ96rw
4rJQQwfK4EDuXWPtNtVCXFCdajL/ycu8PYZGWWcIXRWp0qYp5Log0zOAB0LGIjfPlRBBLDjAGEv0
N/3kUWkCP3HYYSTmgrie96P8gt6d+SMFFwTrr6z9cP82lbQgOgYJyYW9whH5Ow/bvFgufSLZATKS
mBnbsW1Hs2zeCxx58AJH5uGZMMlP0x4MBIiQg8WvnY1MjUrv+Fha3FHxFENuGLdcGEJvt1iSLEN/
EQ7qNzdFwyoZ5TDhcWFv+59utupRsdcE2Ovylo3xLO0iyTzcEcmiENWJG88QGQ0MRJnpdl8Lb3RS
ZBjJhbv6lDQncC6q6hvUA4Wq+NJ26tx8MAKCIltF239NF7qzG+3Q+zN4SMHNVUbUXpAyDuhwPwo6
dwF+LWwGvPEnSN/jMv0Vx8DWnUig3zFOirAzOMop+BfAYf7prGdUK/JebLu8IaMK3pFM6W9GCFVm
ua0hkN6bc70TbZjAfNo9poMdZqDhuogh93rhRkYaTJN7m5DnklPt7IfChF82bWhpRN//lO5VTQq3
jAeaW0LFFK17S5Gg7kJzrH07mOaVsb9/zQ3UppFOS4TEQ6Nvw0dyeMcIQhwM9GG4/X0EfCwLVObz
nYikqmRHbVjxo+7B9ueXQO6AzKzSGT6+dKu/xQ3IeY83zN46ixSNmcJlRaqJw3Z87/DyDPoOCqI9
aq/CqH7Ms8CzpSG5IcoXG/SOc+jvSHMZk4ycv09jZ2+NuetMP3z9hm9x1eLMDOCCfZF4bPu433Qq
+2iOxgzdjJrK4jNRpHRb8+QIT+fVJ5eFbenBd/dTBsKXa4poeTwa87OdGk7BVZLclOU1WlY9VeWX
QEuAsEAeal6q0YVkLtLEm1DXqkq8DV7D5vZYdnDfywj0Z67fFL7K3fBiud49ZjtbbCM2MMCIkXQ5
NsPoY0KmJc8t006q4ArgRQXqllrZH2e/F/9vQW3ELECQeGUZ+7NE3V1ivrG9UEoCtIBzJYP8ApDO
zXk8dlOzXmoXrYB4IjTUgHVTPZwxASiibUlEiIryVpBS0+D/VfCWJljmt4cKZDO7Y58GWPAQ0xsP
/UJ24os5cwCvNu4mB27ZI+/X5i+EVQppC2wYWpI58JZNH1QoYDn2reIg9W7eRpRnx3W8va4X8MHD
kAljjn55Gv1mFArMXtvSMfx4YaCqicCPScP+7BSAQ257FrdyAAE8I7AfYZptZKbuNpgNODyBmyKs
YtY8KetOglGt4ncvHvtFpnuCP1komSZtT6hxnRUE4NL54iQPvrpjlLkTUDEsbwCHvrVFy8g/c9gv
4q8uAcZAO5Na7a3r38m7OCZITicfcrLy/Ad4FAW6NyYEX31yKuyjTlGwLx8ZV1feE127bo/QE5/E
qRYUGaLoBBFC/cc47DhEL6Tce39LVAg3l0EZZ8DaSInEu25Bg4D0ibbOcH8qZEDTT1US5NW0g1nY
o9bf0dlE/6A3juYgK0p1iDFY6VMQgBOtNhnwRKfXxGXDYu49aVXHTBAoFdVANsPCOw64joQ69JC5
slnFr0bhTIhN1U0siyPLmun8SIhYT15EIR84GmaxmQpHEWfhil3/52epnNK8m/eGbYxjoBCbniqF
NOVekmjAsjtW/YukPuNKwR8fPk/BJ+DN3x27AFwmesA07kEN+pExvgD5JLhOh7HmjXeMaW5aonGO
EDMGgU6ogBxm9xcVAf8xk2DIKbsbIoJnfy4sR7ZTc3+0UGDGTv17wVMqR/ggVwggVKlQsFS/P2Re
e20tW6bORXPirI52FJ8nyki60XSr0J4QFY+leE4NhUuJDvYZ1l8LlMJ92PuKFnnBhr3uxxYgcjBG
PjT7C7PHp+Tl8l913eolgegAUXTGonB24xFHN61P/wYrEEW8n/pzPsptZZFOhSLGoZgR9o7QROUs
59bBDqvCzYEWBwanHKlEwF6pe0d1G1ZaM2hGozoALdfDNTprKHcj7UV833d27aIqSTljGWrrT4cq
sRNIOd7JfLUeXqluCtKCP1PmaczBuVeotNlo6uf/WzQNQdjJzo0WdQYAXZWjQYT+RZAxJ0nUJWoV
EJOVsocTp26ZYZT/Q8prpwBxSwk0eqJZhSd1WuErRBz5NiDAcKW4CjMcYvyROYUiPC0Wd+qwX3X3
fNVOLOPHK7SheYsVMA97DVcP2pcDambLsFFsVpixOEztdQZ+THY6edH8a1dJWM4B8gmAYQiQA6ub
Gjvbaoh+2KKc4+guL8A6/JD2+asVFmxJ4rB3ctQujQ8ZSMHq58ZR3mklkNwji0mjQNB8gJ0o4Eyu
nlEJVjTXJB1IyRdxHeJrXeF+dquPvlCulPKJfNqRwLXef7T3ayuVmaccVcRI44xPkMfmdAowQGm6
qMoI4reu1Id2pEAwlq93vRYYGfbDH4+lkuBJToU1y5+bH5DbJRHQtBjGhCwzE0+J0cb84wqP52ki
NMsSaq9epsKAPsGlbubfLCLH8XSIg4VoCkfk7CFrRs5aHp2yn2FJDJoJysq68x+wGnNY9yli3uf8
am26JT2uBXMSN7xmtDOc35ciN0pyM22Mbp/I3UegShsMlITHSioYPte3pDm0u/DB1YUMM2K5Fumn
2N+OFhslNJyC4Aat8LC69TKl9A6t2C25MG56tlTY2jce8p3vhL/4RAjLPaYMY7879xczlHV+FXxi
X6Bw70xnH1SYRPswYNeZ5/gFPJNWn1w24jXk0v6Ra0KYhKkCkLJHD+9eeKrF5mgCU0KuaIeLD4x5
/89ODKSVaSTfwl+mFQ0q44t2yY8ZsuyLRvC1FN6RRAEMo4QOaQM/sITD8ETBkxVZW5a6/1Jhh4Kk
G7r0oRFygpU+UBQ6qyGgIF1vEzMj38AZD/NQn6CfwV1l+tptBKH7xfBTApv3DzauGWDBkI7Rp+iO
Mrzkks6meAY65a6IA8QNqTF/4pozJrQNZ9HekxoqDaeN8MOGNDsI2g8Z/+NteM810cUD7LqyXQlK
/DA5YuLeoSUc+eR1wkcxge6Enwni5jkfKomLXvUFBu4iQoMkFLbhnsCJ/uZjIfanNJbZAJH/nS0B
+kGAToKglyt+tE0YXA7CVK4KCyWfcf8NbBNdKArtb2IJJfdAaSfZyD77Mrvjwt8Crg0aOPOir2tj
vVf07/sQFzrU1y92jdqZNmV2BOOdlUVmUdi2Jym4+WtD1TMstwbSGvla1UbNoEMV2f77TOJupoHw
yd7ytZy1tdwl+tDqTP0fogS4TZZpOm1IkH4RT3y3/B6qrA187nIRSV6LRWr9yoD1/jjIoXaCKJwu
LYYoAp4XCfPPfi9YSnEO9Pza0rAxVO8dUrAmmYWPjM2aSn1BaDwVY2M/Z8CZsIInIyTaKaiE/dX2
3PXv7t4GGNymmZnNyT2m5ES76sSb5kPIjtoPqrxkipmGv/td+xCpo0TMZSQAZQO3329v1bKoTFXC
VysUeglPoNQz8AgLO8WtCmXSQScwlHTKyhooHa4/g7KC0cFavazEhOaKFTsLTFCmjkAGTlk1x1BJ
0TKEs5HsgELl8VuTw8pVOT/3hFRK2FRins9i3P7fzb2f0KLOh5//13cEDvHXSMt36Cz77TsCRApA
YzG6FHDYnx1ymSESdCwPU6JyrMp+J5WxEWkNRWOJhN6AWQ3JtaKzUgOGvL4+06DtLBn5xKMQQNoJ
74nir4ud9YwlgBtBKMfs1CU9vrGEIlj6xq8gp+54AQdKdjUhdsPo8ml22F6KqocoFYNswJQvzzkq
BO8QYU5WpJVF6/7+RtYA6+I756gV2PQhuEMKiHHH5HZkySDASJM6In7NZJ9JjprTln6dKTAxOkrC
Wm+N20RIlFBIe7g1RZPaesMVm28a0DYEwDKXwmhKKJUa251l6aPRdw8z991CNEkHnMZuknG73bHb
41VR966ltIwrNv8WKC2b9snbt6md7kr8yXVSu9QwR7laUwpmmCPaJGoMLfRobpSB6i+2VfFsc8vA
jDbyuDHLh7DMMYS3A5csRA4uWuIdPwjfU/jfhnV6U2sWjfUmFcB0kIwD18AOJD75flLcTqLpaF9O
T4ralFUxjcKE7pgCGTDx3U8gPTJdNvHFZVwxgx+8WL9B7Qolv7ushMZKp1clBrU0XFcZQdrEPhfi
JD/5SMs67/X6jqi5/OWkaRAdQvGXEAH6445aQ0YjhusQYt3zZNmEbYnyYa871opInaABQRfG+3Ab
8xixu7lHVjgk6O9sL0R1TiTiLbMwZOzXeJZ2vwUQeE851dBVebZ73o+jarL2osbXccyAOlSTgXfR
e0vN9hGOAe0jBWSNbbTANJ13JTWuB49HKe03jN9p5gSl0ztyZmeLIyVjxmPH1UO/kt9isMXLmxfo
USmE7Os2Orc/mp1d+icTfFF4GX5p7kfHRcjFNiTcRfpV2x85SHC3LxuUwltTRC97sip35DBK4BHS
gkzF6bh2zpJRzICaagXjXSC9qQphmCsI1NknxabwiZ1FDHJYj66t/6kMFZTX37IAZEE0cfHWosCc
KKIgy+laQpjnmdLFcUrdZwiNCkGQf6bVzWEx9fb+8zKuywncMy7QfFRQDLRTb909ErXxz8rwJckJ
LglNjDmP9pW4uhJbr1ddMTlR/r5xF2TQAKgIR8qV5ROts9scW8xDthxdND6ESuELnf37PiAN5a8N
BRwFUa7M+8jAv1lgXMffyaz8SoA+45kcCRXqhA8LdaoMzLOg0qfJDVHbXqJsNYX5nm3SMsoGjMQF
6X5IjTV1Mlpj+mQ8+wYH1Lak0qUTMXxfK+GeDU1Bexs04cWmMPUvIFCok8Wt4aJehZMTF6VjqAuC
71NKKd5cmQcvnVBdnvXL9Xi3lqpCloQISKw2aIu5BR/XDaEfRrHU4VAXBR7k/uTlXt7HDeKojmQ4
3FBuKh6pyDKNgYi8w21yEgYZzXUS6d2+iZ5KubiDji/r3GraQTKKJsVu2TCQI/FcDaAE6222brf9
C2FLllHJ49ui+UE5xoTP/uQBe/9pgGJkfNQkPqoT+lVjD25Pr8spOK5klmCVZhYpZCW3GYGgaf1W
Von+bDiGg1lDFV2joJNnGDd0NX7dWTvh21YHcH5IAytn0YKPH5qXr2x31/T19uSWTowpSHhKXiMR
hWNj8m80ZDa/U9GvHX4fZyY37gnxv4+WkV5JbaiC9/H1EzCkv80JxBWmk24lY6kyZeG5nULJkE9v
Hy+eqZdeDRQrN2ERGaZ28gTQA3qn7rskQ/ttJ5cvtZzibKIVtLZg775prsYSzyTSS0tRi8ivnm6x
fNzN4leMt+QBBT3G3LIxak2w03vaqznE7YndnE1B5ih22mZYAWM7YWu9WWGLYNu4AawlqYKxcsGI
XWCMNDxTgtCqaSnbLk7aY4yAxVXdXcPt0rP6YDSYRa35nAvjSlLca4LtUbRD4DAmo1AJ+RIoYA8/
KYPv0jx/Q77e9vevl81gsPZTqQrL4qpw1tY8XDC/RWcc9zeRXKxUwRnsLnbQ9dMmlLM08MBMOiAm
zGzmrR09Bvu2hl/MWOcIWtfUltvKPrBZMbuOL61RSfqy+faAoOq1LK/faYHBn5s0Fd33+fh6Y8x3
um+bRb1xVClVWMlOqCwQcQCvSX9XZcjyBB+LBJYOIeyUhVzl8Or/0mWoxx4FJdjZd2Pepll1xk3n
NsaF34pUznylrAEfPwzD2ulIRKIuO/CUhqWWtrjhEUpWKSnLs7Wc9zvdQZsZVwEVOH2/HoxXAx2s
myd14YCqILv3n9Od8f9mH9u/DPFR0Yj0dVKjrLDKTQHyv2oj9OkwVRB5VG2YGOHWUENqbz+Hl1/q
FeOGb6bt4h4lJMzi83q/eOLxeRDd/oNRTC96h3CexyuBp1WMojSQtNbxHrRIkVuLWQVygNh3WNAH
NY/ISiJXOy9hZ7+fwl2U2X6dTlEv16gvKtXTDIaqSZYDoVVtGuo6m0A1qmFcNfVTuUokr8XoN1YO
aHwSn8dJ/N/dsvH9ysyJicMZwPgUkRRZxQGbToJc5lfRq00yWlo1BPcdgkHnOCdiymDiXyTxf/y6
n79xYINYYY3o6cN5p0hIs0Gk4GNeKGz4KEGbTXtGZSHTnBst1q9HmC9tc7yJ9mUM59OW9HFCg2KB
0J9T8zwG8+dO043EASJ52BQs5GB1tYU74X3zyAHYKiogAPxPJOITDAZMx2Tntu6h1YB2hveEp92u
nHu0IxEkwzK4ybTmBa5fp0dXKJx7N/FkFHnmZ5Ei1/Vhw4ei9p7JGHFZlmFrZNRcid0+yH6FrVAk
PiK3oHBD+jebnZl0iAI5NsFFIKRgDtKDxf2VkLni57FpGnmPZAgNdgWwjyHZoT8llQJ7dGQRDrsd
Y5BVrWTFMg6KKDCs2HUKp2uyh9J+6KziY08nzOiMQqnOod/earHx6DaaoAAqk8BnHX+2AbT5r2v0
hO1mXWC9Uef3lNlpusdX8pEI0do4+8u5C2a/KkuxxoCz+/rBjIQETpEZpwCR1mgLBjD+xiRIZgd4
83GOWzB+3yPQ0qa6vi1oMTTXNmFXgxItdozAvzP5WKXXKgUcsunDSbbxw4gtcX+TZWEk1C0Y1pRS
CEYwn1PKjy8cvEt9wZsKoxFkDQ9hyqYqPIvsSiwxduMDmELDp+0we0pxPer7mvgrFIkkvhFmge+5
BMf/LqGLzYfHm+YJaoxWzag/D3j8hB/q9J3un02fDzhTVlIyAte1XAWcj/l4MWL51+z63q7b1Cxe
Qph6o/oGBHyLh4i/F9rqT4krNR4YAqmWhdkiTGIkKJ0pWWWrj1zG5lBFVKELmrG45ah4kR+0IUaU
4Gy8cdFpml4t/Zypa2qM+PksS6rch5/sUtfLPpsFmqTgTpNC/K7GRJZtT/MWM/XCz++XGwZ3fTdp
pZFvuoWrj7p7iL/YsVmOsaLARja41Xj4PBquO9lj9ygyqIhsXAhPqwLbE1ywMQrTgLpj7bXIzbZs
nEWXKZ/K1POy//CfLYsCgoVpm5vWl3l2Urft298ceWlAaW+ojSB2Q7p4YXEF3l4OYw0U/GOtXbDU
El0JsidIdfBNTFIdsvAcIKgLuVdP12lQVeVmCEPCMS/I28LCi5dgqgy5ejYQY4Lg372wUfTiBmZw
o1O6ZHS0gOC8jY702+yQ/P1ud9Pb+xIIhMwr+5tXw5beCFZNRtZleN0GHoAef6864apPGMwAANY7
O6f+e8NPAWk0SXctgSjY1A0R8uQn0IIVFX+LRRtdichWi06Jmvrm0Rdgs+e075Z2xXwHe0J8E1Q3
+u6e2epGnjpUklRLnHoBDDyy4CA/W/rij8N+V6nxgnglSRUUZDMBFURBAKu29wjuCcVj/rQcgdc7
gfDeYzoNSwX0/CRQ2g4EfSPy2nq5DztIzOKVUfemDkVcEC2TzoL81X5P9LHG4WRYGHlJ0CjEhHUv
RACxXFelElNrAkug0WDDsoM40abanRLUyuy8p2JfO1ZKjcavEIZkFTIGX4VSGhRJtyQR6K6Lix1Z
IOhpY+9hsbSw7IXC5oyQLUhlaVJv6ACn05QJp3UrS4RSIxv7mJR7xTI9igJjTRdnvZKWc98vXDga
+ELco3afu4cRJD2aRw7x9UpzpjU19qYTQfA0+H3EPkVlx8hAPM961cYiRk2wqEgOuZuxfQeF+Wlo
Wh3hytGOL1R8o4ZQ/sk/3VgOwt6rTPVE9AC+4q7bPApCBrnkPffob4WCxf9Gsr+7StesgVhr2vfI
qHq07/1AoU+NZeylXBYADH4zPKNwVOj+AkesdDwYBvvB2EfltGAuB4F0YIM3I9Nsqslxp2tggnyo
VI7Ke2Hye8C/axT5nqHQAdODIvncIoYUad+5Qp0hZRCUKxaPXDIzbagA39NBxMhSUWdv0dB0IFqo
lydQ9P8DxDUCUn9cj6Q5z/y9WXlMGwVBD4mshWEZyXooWuu6xwj7PNe4TpFUG4/MpH+TZJ5LzV6E
r9iEavxgEt36KJwKmKvuJgnl8thGnqcGduMP9XIDCYBRiw/HOn+P/49nbVRJIprKpxiiS6lZBvXX
p35M9RCEZtLdmivIJos158FdTNDTbBz9QlZnhNEA+7czT8us9gVsKJeucwuCfMP8mig5YG67NbBw
f1qYUYE0jNEfxH1jV6XB8su/wzdbaONe5K/QVKWgeytOGxnNk86o++KStn4B3M9HM/o1J/15eRBV
9dIn0kpKsXveNslsVAkaPTTxVBhAGQH9Avd7pNNyE1pcj67jGmX0OHIiocwUrPOfi/VY/3je8YuH
heT4cIvS5he8QNmEnsQT8s84VqVB+em7MdtX13SdWybVyyH4ULvOg9ZiZoCkVdegOzGeXORTGT0I
3D2rXxfgl+x3dBWweOV40pfbRSo3lFSkxqPpPhX5ASWwccd4CRPP2ObIp6/WFWhXoMJaFXVSNTzl
b91YFu0JXWk2t9C5RWkDXShfA3XWr4U+QqCGh84/eQQuM5+SohInKt4T1YiWrdzrcAWXp+FoHFMu
CTTUz/O4PsXQKs5zF7mjzCppCZKgvAE6DNLAUjwBr+QlR/jsG28kmIqAcScyZCswvYpu0NtViTFV
uw0NNlOny/WxKVBqyyDVVD87tMXtBhmRjWXNVhbh84Gr5MsBPlYtE0n6m9+Kb16G2EGkICYLx5Td
GZTAkS07RR47Ce6bg03GLdqKxXEwmKhpYGEXShfpemvkSt0m8ipfW+Ax6dydEoKLn8NcfFwF/DvL
/NhN6fgOfDv/ApEBbloosjW+GTm/eq2HgzBiJavXosreSplBh4dj1sipY9YGdNumkysKvmGGSPMT
5/udg0dElJmg6Zx80fZidN7fhcNc+xNeTPT3yUtAwwgYEYZ7Lf5zlV9ap0INFCOpWHHZEakpRmk/
jAMo7ojXHH21+S6UuAexjJ7fnlXnxTmEh7EUcm7e6qVEhLbabXf+TJUzIRyO+p5FAbr+r6hBd3G7
5aMQhMAjWeHp5Ls80YzqPi7V0YVWeRa2el853Q3MlRNXo2PhsZA3f2CIYFlme8f1uevRRZRGKAS5
PW40gjzEaheU7kmUFVTZLLrqFPiTLY41FVkkcpvAqybemHBp0xIQqJpsnhEIDjpiSaomtBwphG+1
YwomfnHRlqbzsn+nxB0HIjLyj4pBgGe3GkaMCHFbhU6Atr0AU2mjryct3Nd7f+dPn6b4cO9HYqXE
t1alXQBRfLlMfCTlsMHz1p40UHm3fEGYMyLbBsX4LmGTKBdKzl+Bb/L0G/2eZK0URI2wX+jhEMcy
gQIwV+sG32hUbh4H+JhsjMBLcxIjbPLQrCCnGs7tvsi7wNinIVHoKsWakYOI6KdUKhUiNHdEmBLC
invb5dfcWWTKc6Z9rlfEfcajj2mem43jAiixLV/0NcQEypuXXlSn8z69wtezqSPsnkKmSUtXIz6e
kUF2WV1nNP8SkMMNzRppu8Grrce51tfzOeyS46YwP1V3dT7FEWL4TP/f5/Db1D2LQT0FMimnYAy8
sbfzH4HCFx/ZeXuDnRTyEr1UbAbrgiCK73dHF3U+bRQ/qvBAMBh6TO7soz87HFH6gGtCRrzYY/FR
G0j38CnpzU4Nqg8igNxsFUlkZ99DuP5/0y4jltbaVkDuyUh5MrnGnPFz0EOherynNkAM/g/qaX6c
Tc+gMbt+0rPl+/HeF3RsV6OmclwukW2C6XfDY9il+5EWB/YhoujoXFRwa3cT1R7oR4n0NPVdc9lG
5r2oKPQICi5W9eVK7METUkrB2v+arLz1NWKo8oBXR1Lc+BHvIT5ukGnoB5JcR59Gh916HliHAxD8
TM2+QzfPXRd3Vk03tUl307pqe8LlLtD7JocQGcimxN6hbdFUkXnBBDo6sl3IrnQ1HgAoXbclLcKt
YP6xUyZTz0YFZUMK0v4C5QhPvZ3mj2d6+5eFsx1N7h0Opps8hz5oAP12MN30/yl1LAa+QTSzUBDq
9UrlwAoN411u317nSUdI8mkI2G1cqMLr7LGUSyUWb+hDQkN6EzfxN7jk1Sy0nCboG8Di50GgxVGo
wqt5tDG41VfIlFktrwmyjyhhwQKnkOJlwDtfUV2uqsdujxVrS4bv35bt96raTZVTOhMDEXikCbHp
8sB8lGWNJPRdvk05jZWJa8V3+1UeJZFGZyLaCiwg0C1lb5i0S3ICCghd77enfjdRBCZF8yXhp7CW
xTstPlgrRKy7XKyXSgj+fKbx0JjVetBLf4Zz+X5Vt5z6Lnu3CTyQkHhTJDysingpJAk6FVV9MVsp
/++e2kZNeeIRiBGmcX9scbFLVKMcE/3WLGOymHVJHTJ3p2XmCSh9w2u3LW8awgQ0D/5pfFyr/t5R
YI/2TAGlo/4zrjqwCkBuH4i8jbPx1uA5Otn4n+Jg2ju6S7ysl9K8Ai5pscHiV6gYigjo3bJURIKh
6TJyA7Kwfd+UWbeSFNK8UVD0UOSTRpLpUSvtWGpri4q31dIXYM08uaKlYE+SHY366cscDgyMIYZJ
OzWOawdLnYg0bXQnmYI9yurC9Na26qIjcG1nGBctOd0vs2QgtwXoApvG/YfufHQ5HgjtvqFuxCYF
Lf+BIXulHn7D/Cz76OY5EGi/xiWTt37SCCzIvHq+mqllYCu/u2OcaOXT3+5bHLESkkox9BilHZBv
yTKBoe2sOnZTVTUK8TQUKqNsZXmixaeeCjtKOkyR4Plt2o7iXHhzJTor4yT0H/kR6uSgDysh/5fq
6/X/y3bUdP8RahtHwNY2YhQmB8xFaDBrRQqq1Ru+f98wI8F5S25fTI18tH0IAbYxcB+t5Ao9rqMH
W775g1rUImatXOgy3qe/2emLnOQmEqyjA4gUhWsRzrQBwuPlnhto2OFi25JicFvkwfHWupx9JLKD
r+/wuDukqc9iTskiVUA25em4symjVdBSrYswhulLFsWTPulcLRVrjjGhmtWnBdlyvtb0TuxXtMfx
GrwBJRoIYQklSFIaBFPTxZA0R7OPWEOgPYTguNCcAO83ytkq/BmvnO8f28DrDy8r2yXyEUafOqzp
dTr4L2jSPYD6CmV5Zh9DSp4V8PtCIxyrXcSKi8m3KHgeXL5YScczII4sqw81eEU40lYHKyO210Y6
+yLetZrHqxDk7I8Vr3FuAGXyxFmjIQcnCYBu49x+hqF0DQVS9qA8fIs+UtKFAKK+WmtDSVs8NS8E
Exl2cT0rJ+TA0/cbIPvK+jGxZYKWGvjt8U7aCaQMNG2BJN0182oltuUdoJSW+9o61Ky9mxA0F7e3
9xC9JYaXhSodVk5Vjy4ZezmkvR8RKQ0GgmjF6wOkZHW5ulrmxtUwi3b2o6PqlwXRyZXnYIr/BcPN
v4u7TaahJUlOZp0ioU7/OC774sZLIIk3eC0940Fs+hoDzNzTi/y2/ssSNYQW0bdB8ZtAo/AjQmlB
Rt543Ie5NzzwcGI/AQx8JHV1/aF4sjTjtCYU7CN89oK3sR6EjjMCh3jjCph53/LfI/zVNCqHT7Ko
hWoPqUIxL1fmVCV2scuJfJXUtfYKncWWfPcBgf+2AaKe+jwEToLgzYL7B8WaFqBpXAh91zPna7Qm
PFXgUdQFFkx1GVEGlpBsv/Y4G5bvzms6btwVqyqcTcLS6mzxBmAiwNF/30DaMbkmPjNGtMteDECk
IY/8GcREdpHsh6mKi3/+lGMqvIfXaiJxRnBkmMM7UizeXTB73edn6j4Rw1Wyz200FuRObA53PtsU
V8/vWPZv77kzN4VmGtGhE2KGYP5gY2Uwsgj8Q/09VbhXR0C/F4p3BOdBLoB3FYQpTHyXSeNZj2Ar
lBl+D1ztF5THkQve5pK+OA+pYA9S9QlzSJPX0ho2igEomhC0PYlX0dkkEUqVv/rmM7VxyrboquAH
okmgZiabBfx38rzQiB+ewlKXcfyx2TQct+6bvTIGau11pRwXWcAOLaBhOUt6iMDmESWupMORWaht
y1f+WbjWfoR+HRI4H4ps69yUWVRv5O0tP8BZaLlMk833UFl0EE4EYEj+cs17Uxn+xIS7Y2Jsd+Pv
rzgN3W6bqbtlXza5lyLv0BPBWHFqHySLlin8PlcpRRht0A3g5Ch/VQZAH45YX0gNooSQjKlotl+I
Fa38Ix3ZYrpHaA7N20cv4hYJJO+0nhlpDaeMxy2DWTAXzQHM7Yhvl2SNZnr3UkEj4awkzFE7oHok
EqRXOVu3iwcTRuxdwjz+BwVR7smvf0+rf7V0n3MXjD7Ad7WLsIKvqHwGmFVfjv5mVykvtJjjv0bT
pg9fGdlPSY5F1rG3ZI3lxet0AUbLOUywpqlG0idk1CSqUytEvNJkSkegrFu53lgh0qdaOnbvc3R+
b3jmR8xzcB+wVxsE1427a5MJNvcSnDz5/+Lrxd0hVvOGTn3BkJH8vhkP9525xWhnkaBrK5ftj1jg
S4kIfs5rLdGg/h7h/eVdPTMd4lY8QLXjNZeYuFCbQhHwAdgDz8nRQiUokeMcC/zt1DCImzTjE1Yd
Reaq3mGBp4iXPvTtqNXHyEoUjyLNCWRlnUyuOK4d84Jl69QtF8qXUVP3y+S126thi3ql4p0InZNa
jsBc7rUCMsXzqjzPkPfrnT69CAPlKVjegtvsZ2eVSrCX4CueguDds73wI60anukw5JphV5adIkdt
8iy1qu9w1+Xm9zRG/Faplmz9NX81mj2sl54G53aa/4BonyCX9Fv8fWngLzMYnaI5lqJx95EfzC3p
cSXQRQE/DNKM0X2suJH+NkXNM8f7svZd0bu+JSqmZNSx50+LPBKRMU2d34xUiMXqFM8JYGMwbHIL
QbsxwxqbIi7O4jlLydyj5QolxxNVHN6n0TEWidOg/6zqIhASQM/VQNZjhGqwdKqEKwcqh0LyKxwr
W2uKiwvKca/HlXTkDpQdmMA477V9ISUZm6bTp1ipS8iSzUbbErufew+krEuqYf4EkxwopYcVNvVG
BMQHXvE/p34hGNq4iM0yknRTgZlenNcVBClBTgciyA6AJDll89JieW5Tp6M9YgFgEc3aeCRfDwgZ
+HGsDtzGkTliD3hI4mn5RWrthZnGuKC3psUtD7IdaE9tS1a3+6QCnBgGyKFqJ41/4GMrdZBQ9LyZ
nrpislBd+bTMH3CqEUtPeEGLMjJ7VIeSiB08HQedkAS1OPXGloUxvbcPYyIlzGXl9j4nYfzD9Kfg
9EXOHBuyG7lO2XpD/VM1Jz8aFDqesf1MvLD33sPHKPbykZGFb6QbVuB155rx8G434OVqmWcXSQz6
8XKtFzJystbDSsQvYYDQZUfmkRoVxcYm3t0YtHK7Rb13MpmUhOdrZ6zO6k/5yTD6/ObGgvd50Ww2
6tIEGyibtD6wUyTMjWCew6voj0QS3N3YMG5n9f4FqgJaXi1H11G4DiEjv6Z7xnm0vXqLPuvj4s1T
wEA3F8YRFXwoJnHiqQx6AvqTBQeJEwk2+cdTAvP0Xp4+pXX0xv2l79MH3VxaN2Bo/YFxyIRWHZCt
v3UPr2cT/nKu2ZfwNo/7+XkrNpr1sZ0bQc8p9pz444Vgi3gflFbsUg0ILHn/oSHnVcUfUnqtVwwK
CeW6x/U4UdY8ss0Nbh7Szo9YVLEGmRLZidnfqzg/IWsjTU6js2vOXoMb5oL0fzcgIGnpddD3vSUq
gySRlmLX3QKWgXrgXS4BFTwaINXyPnKaO3eyvyBPzIXCPKrp9RG94Mo/rztq5HbLsXntjwj4Gp7L
ThJPRbj+Q/KB0IqGUOWSQrPGN5L3llPfYx1XpNF4mdVfFFjGfoxeZukMbS8T3k1He8lau+Q1jFxb
upz2ggburaJOrstfFDJw9kD4QsEpJ+urDlhzKyiB0i1mlylSTBoFvKacK0HSZ7/LFTObGQGPxacv
Ls7+msc3NEwQoSObYap1JbwcFHkKk6NQBV+bC5URfsizT0hGdaNf9oxFXNDfX7Fqk1Pbdwxv1tgY
aPrHk0rMuIH7XBx8uPM1CJjAcmEkQdO5NK5kgpl9hCTrKmMpdwPESIaWjpoLp/WUMcrbEfd/xpR7
5utnrXPi3svUUhKvvI/N0+Kl8SJN6ieZ5YAYVSWbUkrXVAa1gHr/U6wNbT/SuCD44ULseDnLNPyD
Gzl6rMpXKpr806o0DumDhmG0dH43eJgwt6CLYOeRQSYv25+53IuFdw3IFItlNbgguiraerlZzRmr
rjs5q2VWI+E8IyYvBRj63miVz3lPSdTCBjee9i5GJibJbve9O5RP6noP7gqHMbCr+OAlBcuiuCcv
DXVAuOohpZ+r5IyX1zoYyaoy+dfq1Y7MrAyUoJYzRRUAMx3ia4Oip2UrhnTfhg2zaBUbmnPjv21Q
+ytjNb72xqIyaQJPskTM6ItZCaQeveAGm9SVtfkLlf5+bncPb9A9gP/Qo6CAGCFH4WCHVnE8sBnD
IWaTXJBs0E20hCbex9JUwrfZV8qsyXm+pt0B8WcrLjyFA3hhKOLPCxTys/QQ2YICyAMJq663DHSr
tSIMLFJAuXv9vXxuWfSNdYrrIBATDfumw7VeAoTKRQTS24hwLc7tHFCHYP5fBbzQPNy4YE4aY+xO
ulRnXQrdyYcM3Bj6aaZob2f69AU5uXjh2jLDzhR2wrHq59metobyFCkvEGQ88qv3fVCaHkbjemko
Noo/Agsw0C3vmbKmDAnldlmREu14rUEpCWaVHBD+zW5+bE7Z4dM6Z3yjTyUP9+DRAJknf8oQ+rVE
+q4NkDkxks3e5UtLXHNrda9qh8WBwxLpTTmcOxWR4CzSH0UgyW+TybmPQzsiPrvkkFkQKHMtjH09
tv2kHZ2xY2N/ytpARgI8Gx51lrWX3+6ge1RRfdF4dP6Fr6lrf1iclYt5fbv1j6FDn5eCum85rCYj
vw+jtbF+rouW/a9LRm3MjI6zxer6loH/sdySvGFOMr+xmEgk5SDg/tcggX1ZwQXcR/hu+cguP8y/
DFU9MPQsvpNbyrMeI37e9Lk/fFXGjPJf2/3l8FlyUJWgLpCoGkRGw4o4YCoiY6j1byWHC7Wfru7s
Rjt94oyCtVbiHBT5PAY8uBzsBsvFZIKedHl/SMS8I+QhYZdHXq1n5P7F/NSXI2A3dtLr6PeaVL8G
F2HvzM9flqigAFEAFefmeQRoNinxZkXHLbMrqOP0drjrYtwLcVP7p4cTdzNYjTlnoQWaaA+NYS/1
j0LpYrOzkgY879wJ89t/eKQ3b8WXdA11N10fx+ZahguSu5/ya7wkKRpumlZhnCnKwa4eioXysnrk
22/VWKPUeIkXQwOMMX+LnuXLs75csscZ3gBTlOUgojJfHkthGke+2Jtfb9mTI5NSp2SYm5PbT5DA
NHEf0Yd8V7mJ+ltlnFs5z2BYN82L44Z2UiVpRZpRpDPo+UnIIRcfntPvyzybIeBcI/ma4jJQkd/S
tBu7eqxW16NXsEAVHw3L1xWdxyk7dXx4w5B7jvOuFYF3d6EzZCURj0JamtwT2qXlap9Xt6lgbLH9
F8i4Xi93DFRFiqYslRZqqs38/NG3PKtNcp/sqx4FnY220+5OREOVyCTIvSo/aM+9F/3JRxk6Y0Lv
FI7cwyI9exhAwHezsTKeFQX9I+NGfx+m50rdk0k6PX0tqRE4cBHa9DbHa8N63vs2jj70RL5FKewW
/lynQ/TI7cp60/pIAY7uVLX6NiQzzcnJGwn2RUo1gmdE/H/+J+VcBIoZ2FaeNs5wxR635dPE5B3K
8x5uKCjpTBPY3dy9RTRhqiawPXAlyCs0IfIRiJzFrYe8ss69o7yNIE9h3FNLpP5qDZ5+Ak7OjYnz
wjnrTCAaNzXjfC91b6/wvDATUHNyoBkHOoMEkrVwrcRWj48s0cKDMtId2HeWKTACTfhzf2w5nqM5
L8yfPyCssZNAopDidkOlU8fdibKIJrGY9omf3vOzLAV0DFgLqtieHGgYbAH2Tb6DlHW5eDYasdfW
R6rKJVczdvV2TtpTHPTN6g0AQ6OZRTFE7+Czi1FDK4jK2aWi4jTt4k3wGP4R+GavULXdtYVu5cH1
Ts2sogvzXzIKg10mfZYdk/lnUvE2B8X6JXSGP0+9SsACvio9eyMZq7p0SOiWFP918646xEnzLBu1
Xg773o2E5trnoNB4Ds/qPFXG0nwJGg3zj88yYB8YaWlGWk7I/2AYCi/TB930GLE6V9UeyiEtdYk3
om5BmKIF6VLvqPgvVuGQW3L5SnqjxaKnlEqeCrUncrOx7rxf94+OkZwIN8rVfN5b/SZk2wm3rMqp
0f/FTkyeHOdrDhG3CPHWgTpK9+YzizEBtjlChDq/aAjp7b9/ztspnE+XF355I6H8Rk0fn8piY07I
1V2zcTXwflH7gY5zd5Mp9P5is17er5gXAYvX033pBCDox8Sko3h40T0eHfWbVVenHEt6SBMG2h3K
vmaut+LbtnRAtNJf5+uI3qgf8qACwMe//uUQbEfNfklCGIojJGP2DGGJpoX5E11TN1HsfNgkVrev
13iitAVo4I++xTPHaNhO39e5x1hO2aukqXw7CFny2Zbef60mBwxwy/Irpo8d9nwpweOyGNwd+F/2
eXR4DCws2rLB5mx9/cHA0Jbkr6Y4zGH+DiaeWkOLE+yNL1EHQzp9BmDXSeAt8z73A5EZRf+KT0XU
JbPk2M+NWRJV4fhPO63Byqef83+vj18cpVOxf76QHUPcmzEU6h1zprYAcdGxhYVi+sJRjCknoswn
UJBKwOKrdlDo8el6R2vtlxbG2Yd9yjaLnE2qkKuizrTuoksC7cod0bGFnFVqsd4hpqCBWZ9L5vBl
Iw9kKjdcbNQrqAIj7GnolQa8vPAymKqmR4n5CG128BRT2YdD80EecgDBjt3Ato1W3yHaqIu4l9uT
g7Z7Ffi6jpew1bBdME9WHPuJeYZ4qogQ95ZnKB0VDTxgqFfqIKbiiUlZpvUAAUnGCI9k29gqHBTY
yt8rWQruN4hekCjRQoFjkwEacsJZd8ZmKVGhuGYROGKRdDkqBF85z+RCg/+NbcHvTYisDc3Jn7xm
eTQ8z8t6zdxgqzvPtjvhOKVaapFl9t8Z+JCQ2+eBsp+VkIyDXiZjpj19KERRtHe/hoUNhKGQ8FlJ
Y2UzJDE3nzWzdM3Ls8+mTO7BUCE1ej43ZlN1ILy0HOe+58BXsPF8PpQShXHcGpjXVlx6okw6oilZ
0yhK6O7UHIzE897KCm9mj3HZ5N4cymBa7IHkMkzUXRqXvUqiGrbKQnqqC4SAg/Es+GOaCHQFwhqD
yC5yTZzXvruHq8zSyjoJ5ZWRcyBVFExOxM44lnltANqpABQkFV57LLYAQiCb7ByKgzCowDyDejtB
/E9p6WVW69OMroKLPuuzb6uxVxIwJk2BvHKajxHNXiaZ6zKcVgKa2Bv1yBIUNo9kJqW0lNIrpcIu
RESfHWbjBvdFbGuakJwiUtnc8mws6L5mJalKgrD4cDn3JYVWpSVWlP/rzjggmT3aY55Yk705fsqb
/Ysf7mjM+XeOHpfZ4jqyko18kgMoQINsBXmY3XzVxLFJTkaWFYtusWG1yrByIEVfUAJoWqiDBjKJ
PldCeCaiSx69XDrDwa0ynfwpq0Eu7t76SP9XtKa3K8o3ynhA2Ga7lVVCQ76hTmZJiMNyhq/dq8X/
noFZ/FNBwzNKG4OUFsuDO2LctgLZ7TndciKRWEv3AwXUrkCjSnnic6k0tOAqbV2G7zLiDyaVxDNi
8FUs8x7sc93YaAXZq3bwWSRB+8Nuw6QQ/n/CJyqha9f+8y1uIN9VNkryj45SrBSTIRpJU2TupUKz
ucfB3lW2NVaXr1kyNWkC/gYl7u0o/YN36LYtIDTgIvpjSV/1JVVChTfqafAHze2VOUqq2GcwoCWK
eRZdHSejQ4r+aOB7ry+gseA4z56DWD7zomT3NIq9ycTMmBjvT844kt19/qzhrBwDWy5+8Mad4oWA
7aMWyvn7ZfGMMbtLlwCqVSq1sJ7meiBDimA7mF52VZz5OQXcDMLUrgg3US8oxBmU1cUHJDO3RroR
rH1rbID69uaDgQWShep7sJm6n9eOKM+Po1kuVOI+Qve9zvP0fvWPJd4ezGx96GtXRdYsGXYRQxru
Bpe5nHk7+wUSLguKVZ2DuwrGAGt5jEekTFhHPCQJzOYSm9v4q7wxp8mypMZ9n6LXGD3dxUr9DSvO
P0R7U0shMsxLVv6iAB1u26o/456AsjvlehB0ynE3H2cPxHvLB4VLxTESdEXaN/dMD+PKYAJwpp2W
WcuH2C0ijAVN11W/mOJqh9o9axIL63/1prx7SjK4n71AXGo27W3TNrQPeriSkg9097eOHepGR7vg
Zg5hBYJs8f0IP/nFR433zQTzuHx66yGf4fIRw/648yE2DvS53VBCAZ9qtBa3x4qgFCZqedEGwHUD
3uUbcNxi7hgS5zQsO5y4halET3FdMr3bdDGdmGDkjjCCQikZrsskehlaIxwKD6zJ8WQvdpr0nV9U
+j+qO7K/3fOZODERsQPFQh0mU7GDmSlGxZJCn3NpSdCKAUxQ15XhbVILU1a7MvKeTkt1PLYwzGJE
7K9okynx9DQ7+HF6XnCVGPABVrlGiSnZihrlMpg4aEyAjrBTkxktb6Wge3JZj91f+KnE5+AhtOmT
fpUF0FHZejmTD819TgO49EFYaafwmmNmiW8aK6vK+kQryg5U2Oq36H2xx+m0pdcMplE9FijD3F+d
BwBWcRqzzqf7ZUsJxf8emiG50409T7QjY0wyayfKTo/G8xUjlbyjrGMMRQ8j4HsBNV2ILnTJuS8H
ljvLpdhF0zeBDWxD8GQLG6HBSevYWMq6LnYn5PYbhFfONnqD4jozwh8A4S/uwhDSOSMddFJPkPMr
ckhvN0hiJ0bqgI+3xB5EbLTLJDp19K0sEsovJ0LlTC4FKND9ENS5r9ISwfeCAgcDcGdzDQHW57Rs
iAccHSF+Y9u5/G/QIwgpz5VAfMfK3eYlc5zpdRBGQ5jASxXul5ozbvHkNdPvYc68EvBqLfEcDWr/
HD2gCtPYQfc8GRJlnzj/KgK3c7zIHt+6QTpDkTbskmFhXixcDiUnm6/iLzmvp3eLZAR04MXomITS
RBnPnIv66dnLC9LZOjMgcb3Cztfueg3U5ueppp4+AliS2QfaS6gRhKVdkXroVdLbrhLRKwXvb88K
c4jTzGGHPH5ZqChztM2pWsDro/uu3JJF5zu/kb8Ehb++qYUdMNUM9zNfjelcAxcG9GQ4O5rN8TuY
tWYgarq/p95eUNMN8MyPdcH9uAOEmozDUp0Usojmk9aI6tyrmhdW8ywbRuPGLMgS3kicB8MqwVv/
BOkQyR8ZzLv9agatJEUIzqxF+tNKpXgMFt5QAgfpb6WMS+Pj5T5CtdMylovhJNVDP5Xbnv5GvM71
PFCbQf0BMXC5uskE9xBzjhz+713j74qzKxcFCvYMdSz8CO3zeYXYBWqx1+9WMXb0e96eKcOZjLLa
TtoRmgfGiglqkDrDIvW2XOCyOiJWDhyGGkcekBJ6X7EnYQgWyL9kEc407G7NfkHgwA5A2/tOBrRX
eWWtA3yJbgYydL7Gqvr3HQyqd7Hwfceu+bcy10Yfh5bXM+hD0M5QNgm2KX4sPnWU3xy3JOlklMdf
de0CV+aqU/bi+GzxTyp5QV3MBUlm4oAJf7G00lwyhl/C3+FVuTypLzIJvSfEJ3ghsboyf6O3KB49
DGGI6ibVOmJPsFjEO1P1Tphjk0jbSnv3rl/hIlwPGFFALPLqBSDoUzbpUWj3Xv0XMHSBL7WZeBPb
KuIGoMr5SPg28MsKVPPzB8mnzBXhILwhNEWqG6QwtKRY87wOwj4vbHDL9RCODCWb+Z5Csv9X5XR5
Ygi3Oj66AxOD+/kThXVjiFgybOB+vood2qs7Lm8d/AOIyM5983zENRd6kOyydRQIjeqYkuH2isao
j4EM3mJ9n604ogXx2po+PSLF+kxCZyXQkTt31zs3hUoi1nB5BkAxoN0V356WB1xB0Zr0M+kzpt2D
u4A99AGbF0eZeUkAqMCLsGGeFhtcrKuL30qKLOCPftwBDFUwUQV8XPg3Mualiy5OrG0KJDuCl+Rr
lO/SRAXIM5Mb3AaBMc8JrTcVQzWwGARcpaZMWhj/C3hTaxu3QXdSisyFLfx8KypAgQJ9PnDNNZY9
pUlmzstm+0XJ6CTjrtJcyHxTu55U68/L1OVeG4C3PuXTpwIEf2AGbOIKF1FwHMpcS9kVihrJk/UG
aFCZya/iNcOrti8+LbWDWcS6HOkxh+tjAS26G2D8tANCNTLpnpYnVOTScAZSD/EZzTmWVNtbRlUR
SAp+LmbkzaeMVbXVZ+SzX3BZ0IZBoxmiRotPDWsmyLTwwAwkWlEczKLXzy0NP66YLzZ0EP0k9dCS
BHmmwS6CqSrt085X6lOe4EaWVEY49A6wmDnPL32PHFJN5HFxB9RKa9gcAkbgoRNgfYWOortzuSwu
ntM0CFUGUx7qZZIBAHhDT5S7J2Bq/+/alcznbhlZzL5/IQIWxVEJ7Jl94QliVgk4lbMvE4llbEdF
CB8i2YI7wXNwwZnVx2pTe+FEeVOu3zYv//teW0wjeAfEVCSZb/5MUdUj1/sFHAdSTaHMrhEcaRas
wTKLrT6x2POz49wDKHwC6nUEb8/qqwSDt51+Ks2O4W7708Gf9hcU4BnIQ25Y/2VnyaDlcDj9JKmJ
2T0wRXmw5cpLfCrDbTVB9loYElM2Cnh/WLeaYLKLZsTNe9wYeEI2cNFMi2zqcNaKQjl58bMy5BIj
mSBbatKv5CPsrC/HLo2gvuYJ/4s5r5bzcnRxGLEk0ljYkG4KSLyj/XM18suPQVvap+pYp/paMGLt
qcdckaxE+rFkccTcJyV+C1jjq7ibV6rwJ1JyBCH2ZS86YQgW1b3rH3zvZzaZLDR+8xL3xVFHy5qE
NQpZe9TijcK239AxazsZMhhCFFqFzEa+EW21GuvPBuVO0mxAvUHdUektgCyjeaRxzJIrAQ+mR4PH
rp3TaWJxjlNjMX7u4iB/X2nQ22A5oVo/lVUnUnR3LAQD3J8tvzMq4CP9YoAA5Bytpe6yzNcAa1KP
ujUxJPt+S0UFpkPhF6w6OPKiRRSaGXIinWW2SgpLY9JUZje6z+okfKjWJ16OYF27xYmgkb5avYpI
gUCHTYTv1uJlIEDzVS2DZqzVQywtHf5t5SRGJvYv+xDrPVnHCAG5xiOG3CkDzTIzYdWQ1ml0pK3o
cL5ZVSp4M+EE3vZDsXufshQq8ajA9obp8TViQa7eGlKfCJGj/51hRNvHGhlVpznCtbe7e7t+/uAY
6nhMmPkGmZ43PSO2BRQNdePB58ABdoQBGOIlwtZqp/ZPeXvnNaLKvX/fjQqESUesqeMOv/2GYeUn
CJDr+gxrSKuZEm1rfUdM86hS2jShggXPNQE/3QIrUuVd6Z2nxIyZHI0ND0IMo9Pyoz3AWEq2z2gv
S7Ci12Ck5VlCmavFLnPt0JGwcVG39RU2A9VfKk/3YW3ysdcpA8lRsYGCv78S4ypxRbQDW+C5O14n
6cK2iSaLuvpTnaCcmIbw0+vxRzQsSg5ZJqYtLqJBQU1zHoVMf05ly/wrOVpTBpPOSmHxyNzhNn62
YWBwWwJpGCoLxNfD0dJVsU+FYaMf9cBH0CdAht2zf527grnPJDY6P1fMRTcrh/uf8eGnhVdAH/jI
NvO//f/ZQDpScmXfiCkLPJaYJKMYCglayT0t9OOFvVDaLu0Sqa/1gBMRbJwT9DkmWjKjfzzFDpQa
MjgpRcpppNbByallBcHL2rWqJNOcNCF76VKFXqSUg9yhWxMHLvwqT1elE9a2VugL+Sk1ChYTI2dv
BzlNOA1PgBCLM8+0UPCTGmDmSjNrzmj62ZzCsoK+j4BY9v58pKbn1rz3klaI6RIul9DYwlcQqGwo
ps0KiYu8y+rr/D/yAjoGfC68Cj5qCD1Q7MSKgMN0q0cmI2lUCOQxuZjCstTXy4UwdQj+Tm86J6at
vRnoXneqoVC8H5HqJ66u1lQOtCYYTC5IRId3E9N0MEsi2lcTud6YEnn0YVA+ShTrZipoDkICM090
nhXRNeVJd2ZVxS4eIEPtrL6IIYHiweVED3QrYkURnl1iw/HyHCADs+BvBlTt1gunL9W90qPPjiNy
335OQm28Ms80pJzpTDJ+YxEl7jip85Umj62giCYw1MBuOYiLHmljDTkX2gACJFB3yK/mrC31dGdl
chvLDuXcgdl9Ji1sXkXXC7A+HCff3WdbQiGF5jID0W66CCzliVBMg4TTN+YdkalaAxlWeCILa6Mv
XLwfCGPYlhIUzeARDYkd4Cf9X8fpojkhE7kkxxyKEqZ76AUI7t10KXsniNwH7qrmoAYejCAYGKiT
2hcJ8ybXoObaNYT1p7wsnktbtnY1QGNKtWqHcblE6h4ekx1tbp4PizNnmZhGmCLLvVBbT5LN/dk/
vv5Fdrah5n0EieHmkKO2YSyRflDsAyI+BqpXTRNyUHUMF1p+EDbzz3JcQFjjkj2438rd0UPtdWZ4
yF69eebnyFrVR2GO3pN4doQNZu2TgG7LcsRTQM9x2JvdtLfAu/DhcoJXRfpyGEtEUAXSa9Ajc5rz
SMUlT7MmubLnHuNtj0fq+pMYDbm0T7L3kPb0rrIghAx8aSZu//4MomjgMTHUI7huSi6M+3emH2Rj
luPokwOJCQJ49MFAjG8/fZtLzSuiEkYDVYl6VCUC4DjxzZolzEv/CpLlgSjR7HCCIsH0WLuIhL9F
YxYR+MVTYM1/hc8icbUlX2AfaLDKfW4nf67u1eOUCL4ASKfOXXrtabRAvTxt/E39/QlNfV4OmPbU
hN7jQNYbM0pc3/23M5Oo48bEGdhTzj1Mh36DTJeBIgOfVepq3xyX0WztAFxqWkAVsIvR8nZbZGh7
WvT4YKYJ6j9wakIMFfIBgX7VTf4CNgga6kLYtWra0bXLf9vdB3//QPpwc/t6UBZuzyJ7sIoXGCSZ
X1NYAjbXZESRbpew/rN8y1/ocHeKUmteJgsR90EFYQKKuMuWsPgyIyV98nxfXKB6+ry9AhMntrR0
eQoIwQjwMFcLCylrI9ihFi5Co84sDzrbGy7huu13F3908X3bKZEnDTcPAdU5mpAyXfIksThqTSZM
uQcR3Yadg59nb7xl88b66lxjELXnchvnaiqclMd7GWA/tbmx2dahlQJwkKGIM/i31fPnLQbqDf+J
SvSIgQ0pEo6OrvwA5p6N6RKPCNSxbsTY96YI+AMbfVn6vhg+R7Nw577+Jij7eLX+4JL0ukO8aScd
MNshlOIxzWTVVwBdWTvLnqTMNwU+D9yH5IwUhCJj7O7Ng81WRseXYj6SBa3e8+jc4z7HlA9DdUvy
gh05S98Z6gBi9Mn+lLSvleQ9iqQZQF5gslWE947BUUgqIhuwHbei2oaVjgzvCpm4ZhBzftALt9Lj
zyHqXthn83aLNolc3W1MNnhSzf1ObwOW67e2WZzb2thDmmi2YtjZzRvbG1ITLTX5kAZF1oa5HRMP
ZaKnjnrku0p+WJSKsnwmDwNmX0SEHBMmaEOoVJWOQ7QcndhDb/9x/nNQKyGqahFLIoif0uMAzTlA
VA6JV3DMBCUQDfkrlleEi3KOFG4UTLUAo0ok0AABGWO71LSDA2tmFgc6NGZ83ywtHfoKvRnakmpJ
dN6fMjE+hKrBzEsGFkRtSfJy0AyN7V0H2Gf3bgkLpR/vvDPhW4LcwVZtKW6SWJTx/Dn4bazCa8gT
2H6L6/WddulmWWW3UMKfa5VzMWhLsfSdkeWd5dqkXtKtkxZFu2hz1y4GA/qLtrtyxlllKXzW9BM9
mZP9T7No1030xXg57LGch9NHDiUWEluJttt4yp9pcMXVKOwaGp4VQNQsAfSy3JU+ujUeeTG3d4T3
NQ/Z5Xnk6REJDKK/5O11HrhjaWo/G02cD3QQLntgJlrArtRUjILWOlpOMICuoPXkhL9g/ZI3momN
0lWdKk3LT+zcoZxxGfkGZ8GIEWb02kdPJUHZO6866awLL6ldWlekPwna7neyH8humaod4R5tsMC/
ML8RFpM5mv7pqVocE7+i4fC2mJBVC29l/QGI2LH3aaAA2oxv58L84lpmsmX/EDMrZlUrn4o0BpO/
T0qq5bR/k4tHC7wvKfGCoA/4hHx1ccfIc2nDLhXpBJV2cX0yC8ssCCc5GiOoX//YJq156U1sHXH/
c7UeBT1uOBhCfW22X8arrgtgSenZ5sBG5LAkEqWXDnckBGHEBhsaID7bPqRysnd+Svpxm3RcZP8z
wQZw5IEAxTRqub7FJ97IYbB7o+WxjjEMpTkCTgcmitLZHmQgiEEh/U3W4Y/4EE7emORgOX4BdM+n
8T/rR88Hnf/KVm235o0ZfyJrHtIWwuKIrPgX5NR7rFG1jeYhbwdakApukPwyID/G/hBDAEYOHk2F
d2eYkSFaxCLCn9v6sQxrZNgR7iIExXkoFBApE3eqrL18jmqXAF3GzwCP4iY+8MzbULUR8Jy8Zmxm
ChGG3ElBIGVHpTfBn8HfDDo66Ki5zTze6wnHa8TDaAlpe3sAjxk2XlKcjNgc/7G2DxVF5EtO7RRW
XbmVTFacM2XToyABLlyBnjwXBp5OgvxhnvZV9LNTaMCJks0Be2KBdEqKGVfmdXog3+wHcDPFKGn4
cuYqAMeictnR19aWFRu3QOrsyMs2qJOR/xg2oSrOLk42nj2bAYInuegOd5YK+anPcFQw1cXBaU07
mlQfBvIN+HDHyz7csioPHjGX+ivntnBsRKAmZGke3qXiznUsZv8h/YNlMErglZpYG772FvCBCmNt
fzI2mHJSr/+oiRISwCjnLCd7K1QH1rAoVvVLGkLC81i2cl4svxQCmVqNcJnKjNq1Xxj1132QCwSq
w4DXdkd4iXruASLvPM/r12A15s9JVC7ypGnoO6vcQ0XVlp3LaXOykS3DArbG66NwZbv+04Po/768
RvTr6Ld6UwFSyhxSwEGzJ4rMVxN7Wm5I2kvIoLhBdZABKHm0iAJL4dNlp7mbFe9V7LpZM8X8lvlh
6NM+I6Oh5UgcRcWzxu+PFZ1LSp0btNiv6yOOA0zUIVm7TcEB9x+E99qlaVqBjeuodVedYneKHKX5
vQfdPn/CjXq+C0rdIVtsyn4/rA4oFmuIPgLYpJl9VVIJZz0f7YmeYpoQ7qkWqQd6AGtR3Xy2z8+U
g2LEuBkMJ3ciRbCsHVbC3P9+EVSprvQnVXRHVnMg/1Ag7AvjSOgcp6pD3Ju+Urm5TFkVL+lx0sNt
RZH6twQ0epPJzasPxeTPTwNTR71yFdYP/Ndafl2HzIDmqF4sdqr7F4CwBTx7eBFb06MNyXVgV/wG
b3uQ63rxrFw7SgM5aAcAhxyxppunncAQOKL1d0fGzOXhzCT9XP3PzqrIP5Hzdzru8LgigfJTgjeN
jR6Ehv2vhN8pJ9rHr8Ybf45bqTNa7MfSRHER7PGT3wyEx4pY5JbHz2piqjeHEqfbC5/s8ZpI3O5k
XG4vuVNoIc+ycROyjNIIkdH4qfOoCreyPmsoZRU1TdXpvIdQU/jt5HYbtz+DI1qyeZEh+v3plVoV
O6ZJVzOXKzhwEzGMpjugCtS1ryakxma+okZu8OQlR9fgiSQ+ztOLij+RLcjSLOOLu+/FfjuLBeIR
4LfblFxylf8rSxBA3MiNaXqtfyKa52JagPy/2/uSQgQ2cPlMA6kQ9TfTt2Bv/0pbuK1SKluE4ABs
txxJLsF/E3bmP/5Q22oxm3VNAdyuiMHu9+8a+6FZnjyXKILGfNpru9fjmPZxyvkk7oNw1Wd6zHp1
E51fCC29hr8lgf7rRI97AeS1wG0ewBhRGDr6O8AflUyHxVyeocD/4j+pltrvwIeXGuIphdTQ6P2x
5MyLtW15jhuQIYn9ND/BolwlwEboTi2XIvpYCprRKhptGz/3n+Kkt4KH0VEOvgMsFYZ6XZxRQPDS
MhgjzPhGvkuArR43MEjhGWcEcviegj/ZV5j4W3b/qSXOunLZscrgyucGxcG8VBR7lXTn3KN1xvqX
fBvjtJIN0i8gSNZ4W2kalUolJdqJ/fps3EhOEh3dfk5fYs2qGYilcEorQmcEyMBA5ihL95+r4izr
VknXG31q+DXMm/UbpDelZ5wwLkLAAaq+vfShT2SmsiueB/h1mOPUy37dCmrfIY0uu5MhP6LSdsg1
SVFGeTpbureRDHg1bXO0LMK+p3QeByWaB30dohzzRx88BMrJRPnhITpGFfowPFeTIZcl4OGMRYxm
37igfGiyHQ65UP24n+e9Q3REmmZy2qOIJI9sNw6q1iEK5HewXgKD+rPs81AZcDEN4/cLuGkP1NB4
/X7QnTDb1magpmFfS4tY1y1V35kpul0SgHGC0EAmc4ZwSng1VvyYaHg/KyiTNmo/b6BxjMmq5TOh
Dz3nlBuMQYYsUpvTbUepdppSRWxYWhFtMIq214CAHnl+5/ikZtjsrVGUmU+lbufXZ6U38DcDuLS+
O16AAFgzFJ+2tRZ34OsK35C1aKQidf0bM4z/fgaN5ge963JhxwNUhMDN6thFWVAFISvv3aOLkcsN
l80IFf73FrpuhytkyAQq/2rHzkLSCXQb2P5vgjGhDiqS0u5dHPVBDpvxqERTX+Bv5QZXQXdvlIma
LIxSt67b5bTEehWP7hGRhjtmQdFP54nuPx0qYmB5p8Jlvkw59n/SFEm+c4v3EhywKuikr+Tr648l
mVhGr2m29M4jdQP1vyO1ZdJEM+dNH5EFT+PukUh/Aaz+f1icpYybQ2lHste/BnBe0hv+d7ET+VgD
hGz+QUkfIKSO8lu397Lc585AObzntp0hGOf8KmpjytcvALPHZDJ6rF+GTj6qDtQXGz1CF93o6Mjl
gQks1h/rmYuCJNxnpWy0SC0WTI1kKJh+RCVSmwDIg7MskSHU6hSZScQimxYdlac6WDvZW4oRvQSh
hlWXuHhNPucsrHSp8D1M/NTVvtw5m3OYXWWopsMgSsx3tkLHvJaYAC2k0o2UFEbjiqhiZodPPXqT
idklyiOXHrnCgHp7zXQbpBi+oCK41hKOaJ9R+dYYF30VeHVvchDSQNmoLFPiuo/kavGPj7W4OGbl
ZjvCWPKaN6mUrDezKSLMPNiu1aRI/uLcxHQFNuDaOn0yZa6nnIJzjmJtSTUIxEf8+QRndK2CQrtf
hO3HjM2bQZ5bJ0y5hhZERIwkHOHs4MuSwgtUuKK89uYVlfu6tQikxZIFv7UEZNWbXhz3OFeZloPu
ZBvqcMyAGB9rX7FcPt4NZOfG+oSZAHaebe5RSlCewoABPrG1/kDa3HPFB+DqoeV4/lRe0i1uRZ5H
BU1wLMHWCgHnOeVsC1B4V3MLwSJamK8PwsXA2XMUWqcqEtkSfXqbUh9tLbbyZ0IlyAYBRv0njCVn
n6LLvzoghPN+LDxD57Rg77AJzdUyzrGeOhkB+50oOvXkeVvANDGl8EsJV0odcNl5qUgWd6Hc5l3g
rjX6emBxDPer5KDicbz2ZtkL0lWYwWcHe7h5dYvDySQkB7kdPRePsvVr8NX9BeJLHnbFrTg5LpoC
bjX3MDj3lpQadovk7Alhbt2RnyhoYjbticjZAzsFHB+22ElnT4YlfKgltRN+QCZgwRnSGx7l9MXh
SsYwsugfhPUUabgpogX08daU6xcQASuoDPMO6Ob2fIyurWiywiBZNUdtNj12/2ilRvsZnITsw0Wc
QnGBgJZHWz3kq9fK1KNNRFu4PqHCa5/jtJ7tnk4KyZ7SITywr9lQMDmI8uddYrmHlI/nGyNUNIC2
T/rBM/1E0urSssyu7QRghdRUUNyafxCkNvnyN941GYAHOeAu8HQ1m9tE50wDsVA+1VPMTxEHVNzx
d+LdoYU+JqcfH6hfSeSfYR7UhEvII5XHXcxgTInmAEB/ghvhB2uym7DM6GXK7x/WzxlMxTSUHUtl
vwjd64ojK439TicKmeS51ja7AT2xauSP7+B5juoN0n9B3xG9GZyC2h5V0uvj9eeCQxLE0SHZOu0L
IG7psekuKWJnBBNUOvpKVZwKgumySv+jTM9Czs7og1iwNzi5g/b75C2JnK155ZLBe7meVrsfx4vV
pQQKN/tq+/aSMlEVMAnkzlVW75uv0czCV1y+mAAcKwpjCzrPx5zyWn0S3dgEFCOUdxacsw7Vm5J2
IrSlRnqb5hjreHdGG658eGb1Bnyg08Xw5uklbFbI/cDNKjj8x/OkM7Sq6M/1iKUZ8mi+vxHwcONU
dH7BwL8VKETQFC11mVh/+VJhvLZQsBJ2xR2jCEBaXfvziTbsSedQ1+1wVSF5yL7WpPjA8MrViCaG
AmQRgqOKT+ysS2S/pJHYtGLQs2x+mMXD0JD4B/GEeuAnnnLrpH/eWE18JigSwUwxZ7M+8V51UF3w
w4Afk8xwoIOG9T7B/AH+g9iI7q27+vWRxSMTWWxuEkKIBkk4SQ9VU7R70Nvu7a8UiTboeUXvXvZj
i/1bLfkJZFdcok371HXZ75o1t6a/KcyVGqog1kDqeXdgqNPgLPOr27dZZg1O5mhzmsMWfJFupMAu
7HCGupfyDQFlNODeeqQrRLQ4JfvaVkGGz/5kLnhCYrfONqImRHDdvxcuAAm5i7m3/mjbQxjakwC0
0amle972Eg/pFs9d4291RIvrPBo5kCAP0TVAIOuZyN/y9ZuNpdFRtKfVCmyGHZ2xVpmuFpnsp7+r
/X+a88+ATIRyFPNjH2rEFgUhOUSmndS4Q099BdB3j8L9DBfnAPtQ2z0fG3w1jyOmbSk4gRgF9UKD
Z6AaEo702VJ9bhvbjOY13sK8n7YSZzfQJJrMa43uGhPwH305+zOCRjfv+oeMszXnegERyTYkEDcK
gyf3tCEQD+cWK5mlmrPwtmXLchnFHjQzECOgDEmzUxwRbffjxXJC25FzPvGm679cAPVnsnx/4x3Y
m6f0bqUWW2+WK5F+yC7ygip/rkWaKACILXLtmhNRNJdlxWHsR1MBivLwZoAAtEwWi6gYWmeNJL7D
sBbCbPAEAfEs1gxQXvtZD/sJSjSPuYA3P+Vouk+D1wEz/L9LYisNwtmCYj0gqXRWDtqMLp78+VGm
IUPx5xypuJ8rbVzQHF9z/fxNy6SCABJsQpTzbdRiVKvIIHEQEXt3Q3FsSJvS5mqEkd8x1e2yFu50
2CsFX+g22srgQiz/xFilteqWxyiHl5g1A3f8n6Yubydq/aWDLeNzRKgAUWWPLf9Gou9ul+6TNCjK
6tb99sCJKjZH76++sy9Cyk1obKW8o1r11rKfD2srtQzvDziBQMC5+uF16dTq7RP2u33mGt2+6uui
VQkiZh7ZKxU7tkxeo5XDr+Bxeb+EJ/x/I6ICP/q8sVZUdYUQTTWJwCx3EK2T3AHMS1hdcDVKX1Fo
RU3eQysnOnwZuahQ12LFGw432BtAjlzPmDLqrX5fxpmkGXXVGvQ+2VM9ERwBDByBnEuen71MCia7
xHhAOSRdmK/F2vRZqVmSO3iyFRmG6HZYSPlmBMcIZGGM15Oq/gRMPl11x6wF0t5bx0WnQDMu5Eco
c4D+evwZy3wx+p5m0nUspnNj3AwCrNuZvNYlKSBWbp8/e1x7tx1PX1Q1v9kVwqY1Ck8ZpN+pVUDx
d5cBnTlV1I5/w4pD5SXkkzx/4vTLARTyGwC0bYF1BYEmBEZt2m6fliUjxJA6lJ1uSsfXfAxbstM1
wb+nf37iL1n8nPquc5/ajA3LVEWGBA/hfKPWT9iq+cjHuAJlYC0b5EVTMGO974XaI6MeqfxrtXfb
vWgMmN6qgh36HZhTO9mQq7vrerlOjUb8WqJv3zTOdSPvBRrYhYhOHakb1EbMfWZBB13WN/rOFsc8
aFgmLojzQHjEIZELc4NUi01r7yxn0FLS6e/SOicgvyj5gKHpBLPy5/hSciAvC5DjgMIqAoxu2ydP
6VNV3Z9cqrPPYrGFjc3OEFItZJItKWYMBG3jb4p7X098dzBalLksOvWYZhnC9BqdJzM8y3GXFMLG
4o+pEz4O6bAod0+gtMuWY0PXqdphEU45eTgEC1fBLaaaYSSvjM+5sOG9ADeexE3mTALRVWqEBoTr
MS/3hUFwK+80iFxFC9NjWFhG/+SWdBQpGEadv7jcnx4RmZVMVaFILyOfl1F0LWBGejkSibytB4ga
2mponOuzZZQWhRfYbViz745xUFGiKrNX63XKqcdMzvPM7xaFQflBm2abuIFkZArAkMjkQat13nPT
09dxGK4LKD3g5chXbZNNAKPC68y5koLfpoMYOwjKqTW+IThKcFmEMIxkEmMJS4yE/XIONZZPyA/4
kEFfpRjE3HihAAJUOQg2yCJdZEIWeJuiJ4jJIhpt7Pr/8Ey+vtiqHMLdCxFb1K+gH3Qj0Zen/2mI
dHsnQSjv6ScU9qIon11yMu3ajyudnaKq/8vEg8eulrvoP7W/3DdYORrg5Jlu0O941A0SuulUXi1q
TMCsbhScroRdxjWsehE12ED2W0VoaBSk8anbHIYMp8uF1HK97t8XL6Fmh7X+2uA6cf9dXIgyxeaN
IwlUD2ywbI2Wl8rTntPVaHLkEVW4usu1r4cs0Dc40YGtKHvL+sI3cE14SQXxeb/MCRN3c038EVck
j5xvMpDmysrnnuO3wiWEc3/AasFmCRBmv2V1FOqjANvuBD042Psk0WzOTYvcbBWCm8JtrA+0uCPi
CijXIp53aD1RBeTfUKeWFNDvK0AyrnCBZcNblwjLsQ7umsDep1QoRmVyAnJrtWByeAN4ftdWMNn4
qYtm9CFKLbxvb70cgMZGdbs9YsorlKw6MEn42y/3B0ynFVs2yPcdLKpACgkO72iw61ATAiiRyd9b
0Gi7h/Bdv3RAMpNAIVjDQUAh6vdUpqPrmVKEfEfpGDW+BTZXUEpzny/5IBdl1JbKWtQFUjaOAg/s
YFY+3cgK2TyV4AVjWnE+CIf7EBsGs070WS31wWfQAITTimHqQhlNT9+8Ohoar9LJTnyBCSMScXJh
TWd6RPN6bB69vgOrcV23p6TznFjbxSaG8vpe2+nTkXG0xTmo5FM25CqVBL+uo0kj2pbH1csxs/EA
37RJusTOZIqb5sUCCgz+kSVXfLZT427wEvAFyFHoEfcEX9oszIzh6aoCHESOO/5tBjTeSSxVHDMU
NFfPo3TVtru4qUy+HNiSWc4feUbrEm7wPsCB520tacZATi/FMOntDCQ1ilvN8Vmf3XrM+pd4fLVZ
Ij8KR4zKm1RXGzl1em+2qWR8qpyUL+bK4b5JX/h6W2Tt9oI9YM05ZQbLnwqFfoCjgreoIDtgr4Wt
5+zQoX2s/cAc8YI3gBoXW4BUEtsttS6towKOiFwaIrdXA57JAZ2maRz+SmBiw3qIEmpeegRkCgIH
l2po7f06KyZP0kuecAGDC6eh27y/dgw0MNHRfVxQthEV+QIANgO9GASGmnN9Xe35MR7WuWN+5/g4
p3Dpf024+02O5f3w2+pJPGhi3pR2XYmii5JNKAP/VHAb1/huGov+G+jEOTCAXfdpHRe9u/k+btSa
t5XYRxIcLmf/x4NbzljDaOTkXF3gx6gGiXbDaJeGaZmERlEJpn8kWl3oVn3ErJ2sikj21tlZZDfv
PhVLNWNq9aSwzeBv9p0iV08+1BN9qcEpqRFkK2c8VQR/qHThS80QbrKdhkC5aqQBhWCCoUlHvaPM
EHTxp3Pt42znqBNzoO/Q/bODzD32BIYpQhvFz5FmHkYmyiEPHJjPuZvY/2MSxO2y5JS59mvXRs6f
J2DX2DimNLOqjqMgU2BbvPqOFsq/gz5ozE5dCNo/bEOxQyCv6KAjOSIX4rf82CDdz+f/R0JkBvbV
bl2kwHPSGxZQttzB5lhn/xxdFTLSxxdPO26ZF9Wx3MyNoHBqjbc/ZZ/JP2H+o+g+2ylgVgYOm5c1
YlrpVdqrQJbHTd9pcIWOglj+Wp9WL3UbKQIOdaz26O1ORLbrRsGgdOTQEFMSmPU/g1kWkrwtt9yD
OrlS3cLXdV8JVqoYeygq4rW6h0f3MXvAgto2y8UxfbJObyKDuNYJaf8GpJ78Xo0Vd//CMjXjUDIk
5E8b6wmGPJMWSG2NInVJGjo9YDvGKH9hdODxuz1kBLLdEPjMK8ucljUrMbWiPT1tL64dh445vCRj
WNwnOjFSjlb/27Oed5oqqTtds1NuOThYSCrTvVwvspWz904SuH9yGtNBUZ4ZKHDeKeQdWU7Muwk1
dF5GBiU/2FI0KkXK3LkFkNNdDTTwhqX3I06HfhSk6yLCqePTTDvlEgXfuUaQiS0YVnAldGemszGA
dznRdKAHMAQE6HdOljhHZDjB+tb7cLjT+Lpx+ADomozDvw1mVTVP9qW1nj1ALbl8v3mkdmGBgXX/
YqtIIY+ZYswRy7JOZleNImTLs3NjA+D265KvqTNiqX2OsKsHIDith7/kytp77pfNZC/GMTjmoYxi
+7+nn8B+p0UcvmWNoGbyJrtFDTvcy5LMyPpBgGluZ/SyYPRFEIzIAHlCvlh8I9clvRfo4pnjV1i+
j6Pb5QbLahxLW6dEg1nsSx1zJ+AXA8BNvZPoZBwU63I55tDZd0IACE3v1UqBx9j8v47EwwFuUTgM
3jl9jRU64m2Q1N3MVO9LkgwPUXNB7nI+Hf5KuL5EbdERK/4Eg0pTm466x+Qj8MlxT1xLZHRk0f3C
KuXw1MPvSx+1swlbY3pN7y3T3DLPTslMkqrFjp+DldnmXe0gtymf53U6duDBrQsVOR4wHbr36EJh
hrTyDU/NKCtuOEKqeSl4Z6Tco+A5PQqIxo9chLURniXfxy3quXOmMAc01QvvHbQFmK17Jb74Ar+P
TLsemJyVw23vScWO8WGrb5YjI8y7sXiJpPnJE5IxHIK1ey5xw/0S/uwFw6gLPuoPaO1CRX4zmD4J
o0SWMC5TYbxqxPb4CBb16aS9b6SsZYH7ztwoaKzPWDVSdPxVcNa0OFa6hmUAn+elDyhvkjEb+7KL
Dq7g6k64z6g5BZmd7X+Ml2vqEO61dVpddSokVu/yaok9v6wAIrZyME4HAqu4VlIov+P25VUnY1k4
8vYDd9LoNf0/NTGapxXrhf9lwCVjMaUSYz/3wEYQ5Jz/31k+J8BbQhEP3dVUFJ3ryVqQNeTIGvMT
WuycfkCkiG9tpgSYiGl+u60cJOYGf/qVTnYaqfn66dhqyOfmT/DdXPrLno4saH1sJJNrH45r8EHM
obn7MDNzYjOvmmqYOmj1YZYKby1QwtdzUNhhqtbftX5ERyM84X5HeJ5WzLAKx4ydV760Be0zhzNh
e/VDv6+7MFdtG0LCxfsYfj0HYLEIjvyMLXZHRYFCzUgvoXj4jbifnUtkXtVS3POinpwFSEPzGrTa
L2RNFUIgy9/f5av2abtDu5kDNeV7V9tIQ9KA5fZ3q/RD2WrC2s6baFiWxXrfRUew7slZvWjFOoiD
VCREOx6OoujRXP0UGVDB4Lw85jAMLQAHiWpKj5Tvq3cUI6F2uE4LUsDaYt78AcWyFh41AMmNhjCY
pXtAuOCJJ6k3h4eR3uB2/URxjExTWGejleshnomIJrmWFx1qrNOhGeOD7uNT1JlBJhdcazs/3ZFy
qexx8BBHMie/H893vwMYx1p3csGVPqRGwkvwX7OzgsUamccLa/xHQ8VheKuvtK4fnABOkurhtAMA
cFPv5friYdo+NSmEQyf1p8JZ8I2fQMSLa110Aya3/YUM+oojoaF24fcct+7pRkH1RLlUslS6puJ/
teiaYjrGVjxb9iWtRkvBo9v9GU5ZaW+Kg1jrTuQKvs4BIjvgFaBfgjA7vKlOyLBSus0OlI5PtVQq
RUEBnEPoTJHC4Otu8zh3djjG46w1HbXCfqUuX39qyV5xxVXsSKJGQNVHBZPmPZCtmCZJi0evH6s9
esAYBESNxCUz3zfLUczJETLWzgvvZtBVUMU1J/rmF52PZ5SzmQtQ+3gUX47oFbSvk4S2SS+n0oL6
42u4VDjRfFWgxV5kf3V8uzp/gjz7mjexUOkHUYWhSrl/gUk5TxtBYvhv+UixSeND8+L26p4+WgOD
ACLKWHf9GrEQoX4GwFr8VtqKGVyqPzrBGrcTVc1EN+G1Wp8xlutPG0k1kg/86JQtHBrfC6Z+h+br
WSoInGcBOWA0yi5T3+5MkPUtpV4U+Tq0yHpnJDtCloatoxVxaeL14JMj4Hzk8VjgjB7iYx2SNe5P
t3S21XBte1eepfKX216idwCpWn00PU3BCPwuuFhWYTIyhkhrDZyRksSZT49ccxTcc1RT9zyz5VfK
lJfhgcxi3ZT7sv5oKFapLP1Tt631TfSBcXnvnRG8XbVhiOsZrYeVWg2DJJEAzTPc7uXpBFGnAGho
6/okE8s3A+MIhlPa95mkoQNVSqdU7I7LZ85ya6IirO9rqaZdu/Wp5FdMYySWnSo7sepYP5JU/GpH
pm4YeQUGgRRzgUftxjrjx5eAa1L2DiuUYqBYFKsrHeVFUxZf/I6vNFolRs9JafKj5M5gMU3dXPB2
7wi38+REarkEsmwio4Gx/2Wk4osNMH1OVBGlO06DE+tFcawX/8mfDvFVK7WaJu4kdLp7tF7Y0GV2
bYXocgyEjBRkCPxLZH7VQShSXurgYa74U2zvz80Klfg1wA7Ch8FFRqGnFAvn3Gx0ycdodnEdcbXZ
vs1glEfFVBTURSYRysrPSMM9vSG75jr+x9zaVPkWXRM5D0sd8oJO1L20C0ZBOtxtrO6bN0+nLkyn
FuaNdVCgab/YY73ecD5X1F4anUg0HZqvUsMlaopBWboPgDj8l/aEzqyWwIuZe+jEAl9NzfPUCG7I
JbT8jXsVGBwLoQ1kh8hDDUgOKbmPusg9ZwM0PGQ2szFR7jQ3b3AMzJKc0m9aFaykZDWeIoj0REVt
iQe/A8MSi50uW6v0dUVNUr/2NLET5+NiUsxFvw7z9cXGWmacDqQc6HsXUUHR8DaeOyIxRoyS100U
J5RokfnIQehAXyJS9kN/sqQcIeOn8p5A8kAV00NJST4yJCdsquinYgdpSZ4ZvRMFv3x2SAkBk4T8
uzBD0SHVJ2VR93cRP4R5i3DscbYTldMZO1Sn+YjxlFN8gpqwoi6rseKG24Kj014QYGkvJxIDxiYT
25DC3PQbPBVoKxy95xEB0kDEAQP1j3sO+iONPqnepdWl3Qw8F4hDIzNgH5y0pSAgzhN+S6caOQS0
34hMYmRDQ8dy0gntqL3GIvZ5wxnxOrwGcPblIBWv6gT3nrr2IYxePmLHR1yE3ve9keCE9J/inC0m
3JSyKFV3jLCuoTyCZockTchwY/UA4NwpIo+AQGQpd6zRt6NexSviUlmclBggFjfbWgGAaUKU21nM
9OPgRqFXS4i/3pns8SIzUPV/ISdfEKJu8EQ3uG4nrQjVUUIF0g/EJYHjsqSrXirFWEC+rUtWQgIJ
5ljPoXK8wtxmCIktoG8OFOVYXr1jBXDTLB/Pr6RjLe51KAmTm/SRiRTKcS2JHIzDwOqtO9v8vn86
37mjmWKC4SMsQCuVCbLE1t/hmJhBpv4wiSZS9OpBSzS7XRnVbk6W3AUzd5h7w9/FDDgDHvE4tHtc
utNzye6f+IAMos+4WRT8piAOproVOHvrYIUnePciFmDd3F1U+4UQeTiznYQQE+Qvwyj1gN+cTAx8
bbUkwKGqCLeEbBUZisWYdUM8hUDdVjKizNuUJs76rEXeWXupsJyD6sdmddMImXS3pE4npb3jZfuC
A70A7jQrzUSe3pESwpLVNm61jPM/zQQd49vhKngQ3j76uHeXSrZbgeMCK6w8/qVyM692XOcYO1bL
WCO57G5FJSOkuYHaqwjDB6Yiuw+NRhO6mis09itLMbB4Cg0G0pXtkPh/YRQ0snJRTjmul4UhA1kb
KhaMBPwMc4CFAwzXqf3vbTvz1LEZdwnbRjwAJYhAD0mucxKw0PTRGOme4viKVMEQb1ucGZnG1jqE
a7axxRMZPYwFpTiTwclYh4W0wb+iHKorsrd0U+6MDdSyWENN47XEQmBOfkRfeyzvYD1lEHnOCjBp
JLc6mlkdLvrnBJ7WSjs/XT8RyXMCkbl6HRmqRTsRNIqrZeOJq/ZSfR6Nu9pWXaDKQk5Q4x69ZcpT
Zp2YoKCWZ/lCeDyIuNAYLdbAFZ1Rge9Q3IRQa5BL9pWlpRTEwkCUCg/4IKgcnikYhYYyhc6TGQ/r
xAcrAc5TIPtKZWSOGx6l0ICg7nPGYTmxTIiR75lmQBTjRT9nx6Mir4m9WpGcVF0EI3ffNmmTjLef
2viy631hFN+UNIMyR/ZWoFH2Azbe/sRmzJ0bDKER+77YjocwYRjo478Ys+yWI9S4tcN4VqCN8IrE
KdP4A7sFeA2LLX8FAWoR2A32M2BDgGPBODjwbNiCVJcA9/mjgn2xBXz4e5OtB2oDP1Z0mGBhB3kt
H/reYvNnp6FP2vLIcnesvFwAv0ACfIaDjBE3Ts2lnV/CzZXRwNjr3mMCLXoN8P3Bm8D+tUG8KXyU
OfnktxC2+JNJ7vYWTxvDEqbvWme3FaTlJWKPNf5Efi5MTy6YeNRMvTN9IGr84kH/lOEcpH/wRCzv
CcwN6bDb2Vm28WMvFyE17EYlQwTbh1bVTEd9S2bWW81pFUEEKX0CB/6DRj8Vu7pzTZcpLjTUOcu/
8bCxXhJT63KDpxFEVPWf60ilMC3KALjku5qV+N1PlGrKfiyZmd89gF8bAU5vKXGr65bpvnOY2FPn
4lQx5DwS/zBoYvG0rc5bvAoFScGPtoUjbF1FK6IG0Dh0zuhK6x7sc0FcRHveM5GlnkzIkaq5MKhS
tQEVoIBBcbCgScguJElxMEj+Hk8X0pFtto6aT3vTC9gLo8FbgSaMxAtsOxilf5J8eNYLfEubAY+/
FZh3UKEI/ljaJkUQ/e1kKZniOp8B8mpUcNNp0E9hYqftLuRjsiCc00eVoDbhmAQy8HypfSYbHiBg
6S0st6/UxL7CNrotUVbcisnBjt+vBwePAnzwwkQN57jG5WYWFps7/TaguMJlVUEj713hZwcpakX6
/b/BpHEG50rPogRUxYfacHB6r/rUTLG4ZktpUo0F39HIZ6ITS/Q5WTgxTTi+z+yHiuojRJpcifNV
VPvdYlLn7SC9OMzzAtD03CwlSuyZeTvp5ZY6Y2l0baIxeDxTO81gXLmTY2k71MG4a7xha78pC+rU
s/Yb0nw/yY6rzpnCgRfU63MLWV0oEtLAB0oFbRtImcgomSQQagNz61PHTlJumDEGeWydsQEAs4yK
CB3haGXkmhE9TBXdEg5walnSugfaKk/nz8Pg3qCaF1LSASYJFW1FKsMVPOC+BE2Ec0zs2+B9McAu
DnG19y3PB4wWSAbB2vTZESMvDEw8W6r4TNSOx98cWpjbvbuF5vGTphNQHziRAA1potvxa024/NAd
WYD26Lckqmk0/HWBeWEtswfjZADcVDduJ5a3o9lc9zlpUBLjHIc5TgvX8eP0R3oYCpsjnRualgv8
es0vBNkfULF3edRnc3yj8/bmcMv8tzMcG066ET9B527XXVGEIf7ezD78Wcl+Ym6BjC3/FxT4CvIw
I2AzDdUyW8enD3zSxYlgNl9l5xWlZh5Mbfs+vTNyKsnXtVduseSJ9xUj3Y5+TQ3I4FRSFo7QzM5b
0i/qa7W8/ycr/xb2ezXupTAY+ZxT2OS/KzJbuzmXL/mR5UJooJClw8qhlD6ggHqMM4xnCkJl/SSi
vW375jfc+mgVveMU62NBkgLMoPGlRQh/NCKYxtWemvfYJclZU9GIncLOZybtIPzq9AffWwLdpyRo
/5VZFmum6SafmyoCVRZLH3qUyqBegJUYOmG5OL6miDNcI0WXdSirLhC7SRMhXtcAyOlayOIrTBwM
KI1WMizI2c/xqJ1cR35EyxXAcH0Ee5t2AR1RrF+RcQATMJtAJ6xXMThcXwzbqqbMh4gGQU6QQrqn
fXT41yLMckpOiHr0exrJ6oe+o4ip7SXVXyhMc1ewD5hV+a0pcmTXRk35oQw0ZF0a56wkNfbx8Ar7
wqXgUqde5/CoSUp7IvVU4TFD3jpwrxW1Z8du0c2UWtN0J1e/KC/Gps0YctIib13BYOE6f0aJHA/F
0ckptRK277srdvj4cpMZozEN9dt0s+IbcVOPy7V9RG+HwJKEsmdJFEoeaiECisxNs4VVLiq5LSLl
ZlG2b63O8GdYbNcgeaSdnrNr13o96Vb8x6ERMXfC5du31AQGiaSdnWuoePVgtmIDP3hSPtx9qiH2
PdPTEk7qaCy7FkEi+or2icm4pWknZwZpBy6EtY83QdxjB8rPqksTrPyzqiITqwI7ZxVGcz2cQVZi
vna6yhcwZysg6+5MRbsu5H4ELVUvGzGXkndrhNJkPMKdGMtUe2W2xaNJpExiN4+pcnPOUqwgXS0h
CDWNKVw95XcIAcEAQByPFRuo7F+iL1Yv9UFmqVe2kZ2KnuNVeDE/6b/3eEOInBSFuMr7tynjZ6m/
dVCNJSqrGsfxqo0pG8rCuovEDWJB4+j40viHXGzp8UcB0DqMGjtCn3V/BnvQ4m/z3r+DDpnP40Zz
oNKSGMSjrofH1PuGrAXvwusZ/hu/NDOiFY2nCckQU8LX5hHpMSyszXcw/NiLlcWNhZyiUePKrLwA
CVaCBtVlJ9nMi1Gw4N1LvJxE0go79kq2T4/y0vzdZB/6SUK1LIanB4v5Mc2bMlPXGoPGQBzEl8mH
j6bghGz11nm1xNBPiE7XfF0QaStS8xxLZniTM5T/fAMWy0XBiNfQg95RwxIWkEJ+wa9U3OT6MEak
qg45TT+2Ubl/7ZB58vC9Kw2A98Sq+oQ1niQdDP7RbtE6wqNqSPjpn820L+ZqN8s+UCVmNZJPkIl8
AcJ+AuIJT3z2kTpk34Bda9rEVP1CXHTH3sLOqZ06abmRciNnlioT6kBo2iuSpQLFDDNokRfUaGnJ
edaH9rh28HuWlsFwca6bdDBbYaLJkmBsY38ivvuzOrsycEdWaWe5oeFwnhI+7blCpFgwMNK6o6vg
gI6guCG203l+U/LrswfyYBhtfpBPLl5I4+z5GxUT8LmPta8eM6FuX/GybbuFlxJlY8UJmDYl0I9n
m3gdiYhBYCsvbMWw1X0MjEt3zpZJAFp92NlGjw3P6u76k2gld0Dkvtve8CfZjXRpjFTGYiv8u0Ti
bjRPrutmm06gAlyFAy5+miAe57GtlOWVquTjepwMdps0X0S4BpN/G4uUwPw6AWzu495aMopdE43a
bhJBgzvh29J9KW1zE0+ZCdm2KvF262fKtYHYo5cEUcfvlqV61pD2gd9cqWnxaf0z5HaY167vrba1
dce1wiY8eT5A033dDD/mkLCSv+BKh4F546YvGlWorM+zPW2czruCDHXec+WOAWpMwhzLsaTm9e5B
8fuDQx0qxfc8lIjEeBubDmIX6eUthkC1NBQ9G0T9SDVg6WHdSf4WE91A5LwhOl0x/r4wgxtgEkod
Ki7NVQUTh/Cv/pBc8eDkDTAd8g/yRAUBCm36DlG8HCKdcYhT7+mGSpFMMH1lb2bbLEdxKkHCQvSK
O4QPCxdBcuXY+85Udc2MjLcxknpOGlFbMDZHqbXS84wZkPraSpMoll3kQD/2G3b8gW9GQCETduOf
svEN1KU3hH/BLXcBZfE4BAfALhvHLr18pHGPxV+26G11So4Yw9a6ifFV2VV7Eh/Jh0g0jp3RteFS
Uav8VlJn5XVNfgds6aM9YTbiR/dhScXospSkMhp5wAzUIDsjcLUPLBLK5WsRIUGsi0bndi5qx8o9
pLHTg7g06ikN7tHqWam3PErXmx87qvnYlDs/c7D9xriR55YMgG+3gBX7yFcfCpFtS9q81Oi6osio
57mlaej8S9rZPtgxEe6cKAOdCkdGPTQsfXDyAU3RuGghn7vzxAcRMFNmP/xvaDACqdq95I5XtgAE
oFndWQqgMbJq387BFpRWubyi3tH6Y+t8AN/C9ypQcz8H83KEuNZcWsFlVJfkkal0RzGPYV4crIMx
WYT1b2bn4Tlzv7S0z5uxKaXTzUbXhMnHc235l9iObYkr9ndxveR/cOpsiqAQGuEFU3MAF0h2lJtH
w0LpXgDorkYxyG5amqM1nVz5fD3+GSniUfD9pK4N3p5BexuDnTqoqazTO1Rexcs0yYGHsguBwCRd
uQDJZb1eqTgGv8HbuqA0gzG6GRVR/HX4Xq8lJbP0jPtJqK5oSL0sQ9QqZ9tkA2+kiDO6C7rMi+8z
ckDvW9N5neZokZuOpj6cfOlCkX0lSIlBRMdeVKHiCNOORyfI+zD6dhUEJYusZScb/i4ho+4G09AZ
53ueLmzlum4RYF7bx6zwIix6N3hizzREsR8II8ExrLtQhVBkNLP4/IDGGg5Uuo/Wj4/91Ojkp751
bpdpqtkYq+TC3GXwxYo0GCPF0zIcy2ZlmVbaNw0aK7VBfQNuBKX2bBWUehDEfWCNFna4K2Rw4yfv
hDeJp7etvdhgL53/upgMthyqj4ZegczbenXrZOhPkn+aYVtEGKmIMY2wgrfRpmVPziqA/4Olvp4b
XdpIuS1EmR+i2tfknzfUQTilw0Hs3Gozt+m6Iigl777HG5v4o0iwVNHWju/DL4lK86+zTEMmHSTT
S9rxwa+1gy/1G0zle+UBF1h8Igl3gnoo5UWL688XuM9RVAY3VifxMdVkblDsgQXxQiVKj/gbjPdc
IZadDGZrQsxRdjUyFzFzkdn07mjgBGR6IfNB7uXFvoPTYpqO2zz3HbMONa1j3lJkXQ26pyYf1dmx
Sxxrj+poLaQopg4J9Td6RCzCSh9GE8YRDQ8mWZ0iOWsVKV+pGCVb4aQbQBPrMJ6qBybSsMsxmtZ6
QLDF5+vfy7Z51r8uVjVZrDBnD4ax6y8ibPIRbvMyqp+ZzfUf5i93eHhNG8OA8fyLlXedX9Ddhfna
LlL5a/aIy/zZD6RaR6wg32v6ia9yQTekYOyLDQC6ma+RSuCO0kcwZOrJnh5A0DLCZeWspmWI4Pyq
00m1s9q3XNTv2LLmB45x94JwXNXa3/B11UfrPoapxC3S/2CRmHDPDmGjI92UhhJZ1gSzIqECr4V8
VmYCgse3RE9naiW5dshMSInxd+92gWLZLeNO84bAzQy3isODcfxLh1/Or2twcmYeSizKu95w2zlc
H+KgSYMSVtM2PU/5vbJhSQqQHupAGfHgiDX4xtF8CLgNJBp1CZfoFJivlnJrc+IQzeXa+3kFdG59
66ta/Xq6DrWe+F4vLqgaFnxkXUfRWe96yVFY48wl4t1A9GehzE7KPFzzQ2lDxAAaqwD7S0bUGRk8
RZGxUZIS621UxWBmMNxsuVu9dTi8LWGoyKDCN44rONimxorAJB62KDadsD3gTzh6GIfPz9EMINj1
kEq8L04wACRUGQkC7P4AbMsgAOtkcdY5ARO3Qjw8QFsO2/VeLcNLA0mBGX9hU4B3R1pzvVJ/Wgol
3UpfvE4eyDGFJax1SfT/nha/6e45eahlo+/SSjqmzOGULwhvO9Vba3HU5MouDzwQEgzKyAtAx6gH
2cW5ij4Sr98fMbaDTf66cEEimiGs1iGgyR11w8FWQNfPJtKAo5LicoNLLvFBiLr+FUTajxjhvzTA
o3tpMrcrkjcTc1RoMSTh+YA61KWpKUE0vTgtn8K0CZw65jM7r+6y4T1LeWS66/tIsM5IfiIITgqk
uo32C+IxFnCM8wXBpki3Js2N7VmJeEZmi2dbc9tLZXMtedPxo3rY0pN4kevL48qnlyuVtTCsycMQ
gfD6c0Emj+5RwvHR5gkewjwE7vPunWpRibNMg9rV0bqpJMzqTBlGUw9gnNAFUdAequlhDpcrZ7xL
jgwScRZ98PU9DfFcFXHT1IlPBZ59vBDPAAWwu5j5rOKPEL+2izJQgeLYTes86gofEW0sEX8HY6hL
tM8hsbNKYsBos0rIJowDDMmf/Do2TzFSdHsUVV2E+H2cm5drdaTkxw3NnVtuAwuvb5kqukfxgHCa
Z4nIIR9h3IhHcz/L19cUVgeeZPw9eJakJTxvvO6iGJmAKG7/5Jm1oeORQ1ZYu4rfXZZgV8j0ibZF
cXIZ2V4LV9e4/CJly0VDsglPpdrPPQh4Mtvj0VbaotuSVAZKFCUzdvDaTJ8Amgc0CaWsNFJxIu8+
35uikrDjUOFkoubpDlPGNyBC3iUYZLXy/2g3uz0yeAwjTokt2YnOt6Qm+A6isBSSyQ6gcI0/U3Z6
mhgCWt+RDFZy1S9fAo1E2xYLkP1qaqelcBfGbSOvGGmwst+V4GsLpoWK6axJ9fxNjtahTj7p0VpK
OftNE07CfSSlc9bEsIDBEsPAJpxpj7S25pjP8arydAZGSy0uRKfemkIInQl8FXrO5j8g/eSfuDvd
Lv3z8rdFs3U1RKpjfWFC+fPALNzCs0MWG1AawA5TFdPHluUOtR5IzuBypGCuEyPqAoZVMrHxULja
9OWbx9nR3mcFoSTQnQx33strLYHwenhlYy5zYGzNjpQps3mFFUdKSivLi+exWiUfTkCt97EPY9ie
IoUUi4E7Bki2HM0IvibIRwUGvrokf5Cqv9ylXUbokbfwTeWf0hag92bWWR1hd37dWthTJhLRJbva
qQhZeUVAl2CzoPi2vUwoyO0Lm44dXS4G4ilP36G6spwZlH5FeNfMneIHi4yqLzp8gp1M433+h9mL
sYZyWwOjv5CuG8yRVi99oz6YxF3VpGtKZCj/MYfjtkBvJWhT8honnXA+SzsgRF4r+Y1Bj90H/Hqh
hwE7q/MstIYRZO5KAu4H5Kyk2H4kTTHFRrK9nRa7S1116w/qCHfxA/wX7s+Zq59QG/4PaOnU5o3A
4bRvgfqwysq16MgXTLbe5CUeYbwoY1hW6I0rmaPaKlec1xVPrahFCHRyAQpma45w6S0/YYi3JQY9
n90i3wIBgHf73icyjj/6G4jtOdAWKQNFcFMhWLmbEZ5KaUUFKdgkzQHFY9Bpymoo9JDvwoPPaZaz
yjFi7kIvSKcB0A+uDlzDWCcVbNLGrD+Lo4cyvQRo9rkGb3px72lJh83X5PDGpN+j07Cl4kN3pXrt
EK+hpnQp3gxUYw0rmT0rE2BZ5VZRRU3T5sxmFXvRamrm0mcL/DszqpVDgtdKKaYgI8IIcFQwC4n3
1Qj40sG09pFAWP1BLqGO8J/0zmUe+0Y+ElfiM69M9gukUHeJDrNZfBzF0Mnlbk5xVWd5VgV4RzdU
ra7yQnpalPaunRQWw+cO+eALQpRig7z2OjK2LqN4kroZ0hy1Dm2+XTOv3+46pZP1NjMUJ3ZGWaLi
lbQT3xQTeFcjOrT5hHD6EuOfH/g47wprgHvkGRrU2wahNDuXqZxw+tMb+w0QjRbZ8N3X5CEMx4sc
DPrnU0KN2cV42RcuvnXKISv8Fl4j2FtpRBDijuen9m4Iq9K1CnmnxIzWVwQ28cW6W/T6FTfa/38g
VVSMK+L21JwqBPiGsgPSNUuXHEjIOfj+0CwkO1cGciwvBrueEojTFsy8eTgOYmkj1PHv8WWvTdXk
uF8OO3CnquLYDP4mAjX0rGjQZuT/dM6ZCvv/RO/j5lPjbyvTVy+I/M1itHM727W8pDixGcOnyGg8
LW0KJGL6pspUlrC3b/dL7+frAfgyjg0MApftB870MMYSb0HXHuUaJ8wuarbLRJWR1MBPp5K/EJdo
Ldgp3+tiNQHWug52e6Zht51FjP3rhIe6jy2RXXlgoohK5i57fQ/EkoNiHsb+IJoHeMFl5PMFKZMW
0om3NCoemlVYbRf3GjUlVXgMELu6ES4l/7myQ7dNAO4Y5UoPl8nZFva4Ya9nbX1F6QkOR9xWK9st
OUkUMl3itb4jAc1Oct0AVIn43R1r0evTebLgLKvUDWVhsOAgRR5itMhew6fqv6QkDN/IXnUxp15h
2A+9aBSUvc2HmOFqAxEI4KlI10R4LqI4pyfYCodqPwTe7jbfQCgjgBgQd4IZXqw7mh3vattSIrfr
jKgygN+H+RhYDb16c3P3fMOJHR4nKDtMwEc7JuVdVF19+CiLAtUAsGW0UrRhuWfXhapXbRG4i6fB
u3LXiG/wWKgTrdLS1ELLGdxt2Uwi6/4hxClTwDezK7MiJqCJPuNSAk/hmZ08+AArceHidwRyBsxb
60ZStPks4HTJv8XZM/kaiGArsrSJXaJwLXGZsb2xQ2zlCTUdg1ZWj3gMWK5UlJAkEMVGBZ4ATWO/
s5wxuGGRxilX5ZgQUsHWuN9/LpsEuTLg9O6+Gpl4R9qC/5q6pXanQjNC+MLrvkgmtdCQE9M75XtJ
oM+eLZB2mrzB7l7sEmG6PH71uB4mIwZySkZQkRzyouF3BwlvJx9nif9eLr0TaLgRGp5cLt+SWbk3
PwCQ4oj03lLepIl91vdJl5uAVfV4e1opRMsN+mBc4l4+aJMzGN+Vv6DpbFxaDjAUULUu7CoOVwld
LZuClhsNKd0TKyVEZv+Sa01tyUOwbjcPuUHeoElP1IFRkB1lLZxRP8HeDlN9bvssjP+UIJJyHn3y
qDj+Hqpa/DB4axXc0aaVkQK+ETRzZ/1KzwFBvuwS4vbOPr3meLVhatULQjy4C27OlEu1ewtHcwaW
FnS9yUEEA41QJpSKsV5+89Co55zX1KSZKhjh8XHjPVovGaN8QM600tXK15BiXsj/g7DqP0BVJd9/
L2hN4GvQt11Qkj0cFlmT/qdPUE2XTH4LZ5r2EhBXfZz8RtOLdTugoXll9FRDlstmL9LA0maHuOB7
Vnl3Wl53jSKLZUUHNYdAb1gLjSuGfIYbPGaAUj4jI525YbJHHyCMxSt9rpc96uPOKxPYtSO/WqJL
WM7bowALVi5IRB/QuRzrJNt4YYfqQAFOE5dnhJEuqySndroS2r9dOZWNKOJ6i6Ab2VT6iFsgNZ+C
FQhTSo+j1Y6RZuu7XHEV+BP/K0/rMTM5rRtxcqs/sZ8niUrvu9SEws5hYDQ53UQclIRWqam/bjBw
xTAiALQDnVbunjWbBY1Ooqvo51i4JNz7S79dm17z7KZoxxmcZBdg1haq+paUbHxz221BIfpYPXUU
vIkQ8FbE2GOanRIGI7rEZR/X6Pw+YbaI4JQU5fz6+er77NKbClGmDwWIDVV5eQCDixyT8vKokakE
omgWujlS8eOMa/J+6Gm+QrActSMp1AxTPqY3budkvjekcI+rCa5HqI8WdiJwg9lCCcVgNeomjFUA
qtglgJvwuyiLHtuU7FisGEI7Lp0stQ5I4hvaRpaaxX90Mi0o/rixjkFcicYrboYGVQIIAUGeHg8q
h1R4EMdp5RqyNtjH9ajpbX3UBz+3+gSWx+GVZ45Efp9jXc/mfV9nxVid4cYWQrtcrykU46s16Fki
KuK86FsP6exGMVWumQ4TAGPF/0bqDCjVyxVagejkz3AtC1xbTbsiV+5PFW4fpNIpGNMMNhA9iugk
53rf1VV/8KFheo7ffR2jc+XED+K5Wn6g2x9pI5Vma2yTQaqBRY6K72hDrJq1ZVERRoPLGACCgV9x
eemb0PtQlXRgkvGvFC+2ayRFZ9EXwXmJhYVUIA2e/VW2cnEEF03VP1UClPoROZgFou8KsWNs0BDQ
IUIHdr1HZW1tFMcZ6DUgcE4jV+hxCanWCVkOJ4SBTyFgsDw9icJWFNzublldYMqw+4YZw8Tl1gVb
LJ8084Mxq0QIMpFD0o0k+TV9zv/jWyt0HWaLosGX3s1Isgtx8ztcXrezCGJr8DBee+e+CNZOXD7I
0zmyn7B6iKE5FEecdCrxsh77W5jyqST9MZ81MmuOebDaxdVU7JsgjoDE1SIIKoqdBxd4dJLXKS2L
LFXsbXJSZFZvYdqTZnG/KXFVqKf3DCtQA9Wt6z4VEez8Nqu/aUfibKQKOf+OuiVXn9DxagrdzRb8
ZdoNSs7nKzD3+OsIqvue7wZ9eUrwZbHQZoxRIKYg3UaPNbPzKfvsRbFIkN6NdgxIJfSeFa6vrEk+
iD+8is+BOIsMOBVZE6sqSajBR/oKztIclnGnmFpxGJiSU9Ih8nCqc/GaVf8E3sf0TcUaLSzsB5V6
PYiK5KgYZb8ZIclYs0AZiBpADTOWLu9P9lLk4oJzi+LI2ABGLBBPj22elOLanG2QJ03j+hz75px4
dsfM6sWwviPkWtLkgV7CJXtJBZO1EaswksJhiFsGmmH4dFBMlsmCwIDEvaC5BWGmKf1x5XMOdI67
9ykkTwu1pUXllsOyiDICwCWpYsBuaaEWo+liQ1LrQoc7IeOL27XoFftw2JSkGVkilrrFYu2k7kGt
6wMVWoAf5IIMTHYSsFMNoBKaCzvgXuD68BfHMByCynO3kHo+IC0QQqA8FNv3I5lVJGZOZhTNJtNm
1QeCkpS6AsRHqnc9ehQZ1yGE1+tf8d4ywCeTP1h5YbJzSx7Iw05PueihfBIGHWdBp82bbU9hfIkK
JVCkYbLbjCBNsr+Q+7F+I2Uvcus/CV93PfwxxB4SAjuuPfgbhX3UtCIIAxFPtkUmSUg2XC3bA90b
iQS6AavrdgOUEnaKfiSxbKJkr3+Ic98M777/hSlqLv1bkes3RI0kp1thxehnpEhz2B38+Vi0ChhO
rsg/6XHNCkM8BmpsY8iSSzqUUE6RWP+x7snxNYMlNfB4UGeWbEdfgytDvsS+x9AgSuNSX6vq6kKi
HPUQpzRuBkmxAIGXZaiw3rfdDfZXjYr2cAQ0bHL9BfdWDd6y8YH81cssoEIKwF0mBgBvz7ZJ+dHQ
s/v4QBHmHMvj/m9+Se96QejAKDciRjcnJYOkJza7ZveECWkff+UFt8VtMsKJO3qJaYYAPSZWK/0X
pgEXMUDphhv+5J6prjHbka2QHw6ekvdZdprc1nE0OrLlzYuynTc9YGzxbrrML2MW5itFcoEHMclu
W7B+thezohusUTGCtWdkbdPa9yB3NguwTTIFPFXu+c6fsQijWRAbTyVf16eKYWk6EhweAMyiNN22
3RXo4qxpuBh4DW38clKQPgwCyWbgpYspY3Opn2CmVmk/FDXf5c054nKqdLTH/np3fvbqiwoNbgdl
o6Stlg0LjP9GU63GoEkyD3y96bWro6cC/iDGvumFXOxmXLu8VK4MUrRmZlfbs+SR8nuzP2HxJv5+
9pNZ3Xq5tLxztQkQeA3wftCq7X+GNpCSfnS8XJfI1lUUSJf5B6I0ZnWSLBBTjkYid4+xccSnx4S/
vPyoqfBsnDgfR/Ctd0IqenksQylXgvkCyIkO/QgT+7Dxpfd3+5NO6cSv++f1N3ORVDCtFToa9DyQ
I/9Yl2nO2pjNMSJfiD3I2DPZXBJro6be3DIsXQ0Tf/6JfJcKyGAdo+nMH726gyv4sF/sn1hlFUVv
URby3qpg25wrh8tW7myQJ4RTFbklgoVIaNa5b5y+gxli/JW5zPLA1NBFQv+fOw7zBcR/kU855DnI
daJ9ywYB8HMTroy3+y6tNdCr4irHYnqxUUPxsSp14T89PVMAi/ME32H6IXQF6Xb0t85Iu7ZbtFY/
K7FHuk1LU12+AwU29+g+CIOU2lM5iJYea8kNktsqC2uqGN7Xuy5veRcWKMoJ3GFexODe5AQyaHuK
sQotQ6Ai6YXEDR3D+6k8eGu1U0NxSprT6UaR+9HzlKwCpTBW0M1/hMheiwzmn0Mde4HyAliQE+du
hXcOtt4kLRG2/RuoAQP7aJKNCYkaqhgJBG/060ACN1OOFzBpXdgQskDBGJzBCUJYc4x2oX7Bq9P4
5mqfKh0pG6DflqTB0dnRENlnXxyA/14Cg2zyoG1mysuZCYRRnk+NvYoFoQ3zicLRa+6NBTAu/a61
7ujf/6clKWW0TckTp3CvZtLMhRCQAqrWiO5y1rBkCgHt2undLbbJpyo5yENYQ3Rb37Le59gR55S7
Q/hUecG5OF0wYGDsI8AKkn/npXLO23WCyyW//CZkp0gh+95kuaL7jLaucQw2tE7J3mCcvke1Sne0
xPaHwnCD2aiWk4A2Xv+QUjNxYHuucqOQ/GOJirDDv1DIEWRJTraEqNActbqOU23BSuBsjuxXcP97
pC8jQhZM4iMAFbWVTyPA/BXroJ9EiHV9ySIiKhscnqo7IBTHiW+0S9CZUN/xM4AW9zjPafDU4vTt
L4Qo1knXwI7SwGFkbpmxOY21IKVShl3Dy22Ou/MbjXrj3mlrGc2WI2r3O7If8hXWcYw0zTa0jOIO
GP8QbtZyUWCoj3wiP0MAemZyhbqOZFmaQRUpPtPFoU9qssGl6DQpV3vZ4XOPKksuaXKMh/XxwtW2
qZt8HgdQUcgaAIKx3sXU7GzmXkQDkY1sGMG9QtlHijPDVUxh2fFp7DNkzUew3BPF2RdnooSbkX4X
o5NLM2BVMAhPU1Xm8uJnC1PrCNpTApVKChNOZXjjZ2zv927eC4x2uJwzicpqZwh2d6YDIY5YFUgx
/bKaTI5fgZji5eVotFwaPO6eB6Aa/rb4dZXFI22R4/F/0fQgxEF4cvyQSzXq0/Q052ldLTTQPObt
hHamIDT6chjZ6mqk982EMCosgaw6tUFwUezmz5kgGgVXccHyA1SVqbcEIhW9hupPpLJS+lE0fT2e
Nzsx9gRFMCSPG0/vyZz8frt3ukRKxE/ZxjVqDWntktgbHNz5E7wcg2e7sHE9+7/BlyPpLzCw4xAQ
jq95mObBTi4Bcc00dixNpgq7bM4jpqe2jDjzGhjcIThQm2DHuVAl1zOL1kVrST2vSOU7OYcdSMOU
khel9kOuvh2teap2u+bUpfK2zpPUPBfE6ea0YtnlLKUlf/6bQnzo60WuZVwehFHmgL1SwsW4Xcj1
pu2InEWw21HvmjzqROayHbqgzLWYgoK6d4GrfO5SyTJZKBJmTHqfedqjxJDcMcsYdN++eW6XbJXz
K+DiLo+nd1h1gv53uVggKo0DRmW7+49F7PHbJrv+YvgbsZ6XZaPdqAqAteb+CTmJUk8AUdTeEFW6
a+NuVRYUYkt7ahPUVh3XC/pxWCBuE9+dt0uQGnC60z4vxGtkHLK2t84sP9xkjDBLECKYUKrX6H7x
UhkT+Q6MGzMhpdVs5uBrT4iR0jg+G9RMuWzftmSvQul+uAL2cTiEd5F5vjhxxeuIZhPJlPmT2VlM
xWW0RbIrfhe/VUucOQ+NWLqDiVGEEtsmRcj9TWvEY3tUnDQxUvtUntrtbP0Z79/65JYl0zZ8mr5x
dH8Qa4/QMb6C0riyu4nTpv7zGM3GhUuynYSX/cu9sW/PiIKUb3QP/c++aAr04UQvgpyzBJhgdV+U
/XktfciAqmaq2hSbSRPyNpj9s34hYi/HrnZHBfDGgDXKbN6ckpOCQFcuGcBwzOL4m18Hhm5zB4l+
Mp3HFhOyJx3jJjN25WuSKbqGIS7CiORkeUhZdoN2h2t55KDfZ0fcTjQvieTQGyMnpVyD7+QzHMoI
uoq4tAqIVK3SkJn/QajMYQzck0RDAwZhhW/+juBPIyrLdepO2g3L3Uh81Hk8GUqt8opL1CKKq8eX
WrWQoNdEK5tZ8pQO9V87FKGVvs+2t/q1jLRvhTIwGQzxgEk1RqWh05KaGH870iwFZgZJ42PQoeE5
hzdcji/FfdO7uBeWs8WZOUvV6sYNDpS6XPKt2Dw1wX8AkfQUycAfPn2q/r/bP04Z8z9WgDzO/Ksy
HsmSfjC0JNUzUSCWyw2Cl20nfCEoa3/NAD/MRpUZ8aXDIPIT5ubpsxn2yzYIyYP2vmtUxgiDDnHE
NXndltlMF4hJlJ39oZ0PpIRnEBnwkLga0fJC4SoK7SYsSSR+3XQ/tJADqlbQJCkp0mdMfeomxqYK
nyflil4YN1k5HNjdY9UOssCc2kAlYM6V2Mhgb2Rw1VtjzjPdJymbao6vmV+h9ARSDQ27Tz4zNOz2
3cYoH5PhXbEpoDWlWaxCDHK9vVPaDo1ocx9Drjgq9IbESWdY4/ZEb+AkFYQ9L6FbeKjDcpptpuNB
Msb1eR21Gwjfkp7f5OEVhMz2AW1XMKChzPvWzHoIAzpLIFwrt7YAbTfEWvGGSbLGMu8+2FVNXGeL
aQSXzcgocU2JYOlCa4druo8TkUo9SASri/ZUnsD2y8sDBavxZJ7aXnLhMvCKUjyv3xE9LLnFwNHs
TI2Vvor2vsMobH4p3Ci9pXnL8M6DTIYYIxqoMbjJ8YWfU33LJNwAi6pDCVvDHC9kOFpMgMec+Ls/
FrU2ikRyZirOdVG1zgfW7fPSwKo/sfVt8kLkV8z5iQmh/6wz2QPm9dHPp9hMioS4O6YKAWQlnwdf
eS8sUxEjs4CZbnyOIGGohkrXMtXdlgjdmYCcFiiAezRtkvZmh0ZcM1fQGGPm4wAgDmeK+s2lFSxw
9zrUcgnpj5fXmFfiIZrdD9O9S+gLR8bWLKdywgkwFUdasEIHyNGMhL41WRnD3b+GKhVcQh8HstFG
xEhhlUMXkf5Bi64QbjQ7ko8pwWOgdH8enOR6iupp4cGPiXXyFP+XkpUcSs0O2WCW0j9Kz4ZG563R
iMtahkQZPg1MrKVPKMSn+DqsbfkFQ74BnxR8SMSVv4qmR8W7bQiGCdSR5YCrDCoJ4bUgQKX3aJMD
yPVX8cDBiFPKiO4LHexFCW1vmTngo/lrcqycAzjgYcetA+wVMROgcP+MtZ6esVAd1/nybRFM27vZ
l60mottrFl4frtVUcM+JF8iohikoFo/8vnssKzmyh/EkBZ4sihwc5DUIbxi3g1ok9QY5r+4EtYsT
5eWToW/5miXOT7syU1BuVQqIvAL8KjOvx4sP/ElZta6q3UlH6r/WRcAlFC5agAOdvYKBgX3vCHqc
BUG3WAHF448lMiZ1BdfFlc4RoRqMnWRHjeCPK1O5gJx2dLtNQwA6TyaaCcISPvQOuHZdkfhBwT0k
71t4IqxDCOYlMBBThWtsyA+OpQWbgIvQ9q13Pdqjji5C4lcHRujoVsN+SZe2JqZ7c8TuvLMG3oI6
4AIi/vtrcsUYQw6YG2QxKec54efxTbL+6mIq7hTmSpWUu82gUOFLBckWoO8T1QiaYDF8HnPcP4uN
NpaKnIVUnZwXAea3Po4zfW+xi1adbwLJXi043cqAwmQQLCCU6bEE/9GwbSTDHRtwmMUW1WJHu/M7
V13fZQ0gYizxhlZhbUwK17l7J8VHqD1hQtldhvWUWltsgue7TJhKdux88YHmMDPoPV+J/nRFqSBP
u4tTKFNnu1GEtZymzOi/CYlC9pnrmv7pkf8KYsF3NvRh3XvgeVj4yGKjxlBJpS0B59SpwiYjxbuM
q84DnSzK/mc/XHlLLfSxIjjmdAaoJ0KezRLqxjK109K8FI9LIGojUumRxemsq6fKRUmnA/Vp2FIx
0NeNyZnDXTYSoj9oFFEieIJgehdoARzi+rHzeAorC6DNKet6XReBB7cHHaAjop0brIA96SfrXMOt
w5r/mqKhyux0dfFwEGTvRtEBZyRkulLk2e40bLBDovxmSniDi/WSiOCvBlpB/P5uC2v8MsXGacaO
eHMgszyboitWvQDPis2ZJXfnfGKc+OFFpFjWdH04jiSlmDcwwYxhcnmPRLwKWS4eV3e0pOpvn0pv
I/cGi4u8jH1Zt7PzWxdr8W4FeXZ7Bv9NdiRM58NWQOEr8rUTXbtN+0OcTwG/TvACZ5ug1A/pMAe9
GRc5S7kiLBHHZ2VGPdIlSQBIEFqmjxwKbgnqPy/p4Xi17f3vsbbVAElPBFbHpybW9rEPuwQ9yKvT
depcvanHzwzn49ys+zzJNhkDZieCXQWy8JWzqJI+onzadaaGU5539aWOiDZEP8E76njEoIkL94lr
ESPOa6LaB5aWFbRVnz/AyAUERJ6ZmTRmrs2ob2S/ZnuvWbo5us7SZweKjtcGJQ71ghwQrjqBK9rB
QTWmFuHmXaoJVlc1Nbw0UL6SKt4af2IfaZVDVviwaS8eU1n53svdbBF4gnNsFMhKEyYigaCT26R8
0un7BEG5zp6advEx4PCkPan/vtqIK6km0bwSdgFx7w+NxIVhQEq1i7KAbluFUcFlY9nSsM9pIYU7
+US92TCOkBYHLJLzZJgeNYsLRItKR0XS7+mDQSQDWCGgT5+YN0790PBMx4PRRSJaT4bdGx3CaIjx
4WslMgPgCHyDhJ63UwGkQadkyUegIZEQw1NfKBn9JY/V9sh2QnxuljWhONVo0MQ0KxLC0hL5ZfsG
vNb3a69OWlIqhbVBZgEM1OPYTwVWtxmRAMK0qkYPVWnpAqnlmZkoDvcqaxNyayH+5zNDpkYTDJpE
B2w7hw21KqUFmI36AcC/un4MBHXZ/Pg0j5hxQqbP4YVXXFpca+VxuA7rlfKaruX5nFthQGNFYXxX
KEfBV+2Q/Hj0T5zOhp1/AqQVf7psvjNA0UczNprUVhf09JtG16xmgQj2ZwM+nXbPPV2aqScqtArF
53WGnlBUKi39Hz7623+K+fFhZ1A9CRXKpReG4lUr4OvT3NmXh9ekyVIC47NydUFg8/0S6lsWFUw3
12bD+TCJGveD9+l17YuuKQw5aLjvUE9S46gYYsu4MkFmJPSItRxH3fREoQ4DdGdXGf0dWJzHkq6M
DutHBgUhQUquoqPTlEnqsYzDJB8GZ0cy57KXXPELzdy7dq0PRlSIgEBJVE2mIk+1thnYJJwfkW2l
g8idfyzORH9Ir3t2pS5ARoiKUl3nhclSdT2dYSStUCf2UJFflYHO6Xm5mtdu7jWy5QGzNEfmrHlI
LQDplmeRd5zLXUxu15vPdGTB5uzwgzZeHDwgYgqgeILvT2njs+K9fkPIPItEQi+edSlqZdBkFWXw
GLu+BcUvmlwtjSfF7lO6mWy3yOTPENr11IftRXwscXSFeM/aXJX71Hb3nA1XDaTOGWYh/J270ju7
yhQ92IB6yJIvqUmDDPAoZUuVs9a1VEb4L0oX2KHeLzyzmCPQ+UvIn2GIrs0w2y6KAOulvHjVPLTy
yq6JC+367lrLtlO2HvVkA1hWMkHyTGoLyjctw9aqIEMTA2xZ9Efikqrdcz6fcet4B3qduNr6hmVW
oqBUT1M0w9TSOqEf3eFqbMPvZIkPiWJ9dPMAgGi5yEtjTy/DtAHe7OyJEPl+2K0+r1YYYNWFaw4t
zc11TMYospRoCyNCFI076+oOc4FeA0UtfT7aOoUucaGEsehDY/Uq95CCLLgF7up/8rWf1zrjs5dC
3pzZyMyYsOSrD8Q0jJq0fTVgN/twZiPEx40SYkapVZi0fyAMxiC26X8hVO2Vkn68ktcszbBA7YK1
AQLVOswbkA5PbvfT/JJyqBcRw7PeBHlvGX5a5uB24FzrRul7KEBPMonukVgLSX3tqtHi4Ij5WiLo
XIMTgZHQQ4n3g8Id9Zt0jMvo8sSxYDdWg0wVwGXMNSi5AW/RQTLm9QWUYzHE/IXs1C3eACz3gyqr
kD/CXrN+OvNtAetwGUYNRj7jQFNsH5H9xFo0mCj3K67xSE7+SLG/7C7iC4kNFkj2ajRwZ0PF7j8S
R9D4p3a8njvkHkzt/+jtX7JgpyMC5OvmTp/urGl0/Uh3GrtD8GJ9YGPc+sNUoq4evFBltAQD2QAf
t7457SJ9jLxST0PcEMFzwLX5teIhmLkDt/GWjP1Y3/zQ86TkPPvyJHd5GP2crgV10AT9V10MK5hH
oCgf9vwWQ9mhrvU0lYPUJzaDYVdKibYMRMdTxsubnsO93F/1N7FLJIsQ8/v4NWP9Q/7oj+CN5i+/
vpaaeGVT5jBsdHCaV3cVxIjC512oURfHbNdoj4A5RDtAhkrTHCzxRThRy7JFwdAWi9+d5dX80Qhj
X0o5UudrLFLqIWu6ya6lThdbt2zWHyZuhRgXJ9lE8+EdnrOSI8/ofc/mrG2Qy4xwP4lV4MPHKnEJ
zrJLvu2SssT08ttl9wlhldbNkEArZb8R5yaD4D7dRnw1WAox51rbCrvWn0pwwOwwaYds6MjTKenz
BGSKkJ7Tgj2xPqN9bT+qIa8w+8fYjEax6/6GdkFXDN0aOItPPvuTIYomWi2wJ/OC7YmlWiEo9K37
KLa/JdADl4L0PSLPxCNR4kZHw8BiaLTvhgMV4jfXqPMCMOQDxvhWhB0snFgRg1fbhuw2AT82zTaR
eSpT18OtATOB+1Lr4+trBBPCYDdLVRit1WoHkR7OBbGiOP0KbEZRl3F5r9fh/fOOdNSygp1MacY9
Djbwt7BjosS8QMWKv4Gb9YGpBJ3LrQGuvYP0sZBwM55rFHf3jPoWJOoOQHL1KuW2pFfNdbUirCoJ
lonFqyV7ciFBQbSDxUwlmjaHUoitxTr7hevTaOWjps793hmW/+HklJYnXm7d+aO5bHmSMJZbDc7u
P1/OFItSS968ivmuamr7WX/O5IxWxiyZxmvQEobdsy/a7IKLlYkKo4G8uOwR5M4QERhnwEBScSA1
c2LKBjNcOFQyWvTsDWFCNCGkaNXZtMjASTg+5Xe8nxA9nLJcJOzEPby7RlmQqppWn7nv05PrDpRr
VtgQS4yh0pMIYgfOdJQsPJ7aQwf686Ipl7zrHTKsTnKfBD/ZLS5ALGmp93P0AciEqxkrBYBbLEQT
fZBi8HAB/dzfpKhe6zsYqxgg8oxZHs+pPJx6oQNdGGSoy2BFpL4ERaK7iI0c7S5EbRwf8dxqqgIZ
FiutoxQ8lcSdL12cFc8AgyvirQcy08P3WfdraNb60lpneQHGiEzbPQPlu0UO/HpDIG+bb42i3hyg
ZrqwTW19diKnPyvhn7NbJpo2EOY984UEcf5qIKxWWuoLrooGtVnx/39v9zXdiCpd7JphoGQB/J9o
u8kS4cOD4q2+OcVC2RAEyizTaGUTdE0ClV2HdxN7NpKD2L8GAaiPFi86jc5V7osO5w2VxbpXOmcV
lnCyYt7Ng8c/0cAA6DHRtWvzSA5aq8X6V3rIAxt+QEEhzAwDN94toke/CovQS8SdEW686oKdN8Mp
sapXsZg6yQTHAvls/t+36gKbi+LVFGsDDwwlb/0OKDs4aCVy2KBqHkCMNHWXTumQDHgACdWPuilr
dfD5lpNIUP32EYtsR8nS5fW5oNkGmdLVW5klWZJuKFhcB6XNLevugImbs67ztpnl28drr48CDv7s
DUbgbnoyb8lU4yV8HCo+kgdcM+0mSttgBzVqPoBL9i7RH6qe4wohteNngsj2OYPGBIxvtnJbbJyF
WKF3et8OWWjei1+xOxdGzAUUqs1WElDZ0QywlXYW/g1cwT+8ICdxrOW8zqo/yyeeXTursvNMyl+2
OqaYMirciTWd36nH7cpcWHJzjVwKELFvyMAVAgD+z3+e+gRD8SohPCh7jYfrL+y3gobIvRPmCigv
QIlkgLSu7130JApFDEslFIOTf4DUbqPeWU2Vtt2VjrhQDcrZPp63XP0LmGbLFhvGtRY6wgfe0HZi
8Ni0up30kGGkzC5XA1Ob0t4AvSAlAKufRMByhavL1gX1/0r+QMhPnRfzZMv556UgnHmPgo0X8M8j
XD37CInpRn9YjVRwADn3jB7kFWHxBlvZKu2JxypnFk5h4bylCk/QEWMRty0kB326U3gBjeOxebqa
o8ewpZxCNym9qjXJTOgAwYvz27KmtPHSIPaM09MM6LELR3628GlQCKZnIIiKoqfwyfmnyFbitRmD
4+aCAG+cabr/N0AXcodYs0jtvta+9KhJR8KuF/hlmfDtPjNo/B7T2xap2F/cTKcybFz5KTyByHJr
nGIP+XxYIrahwVtDUzIYNgja7ZqvWBlwYhdwZIyyYRNt42DitILLGGzTv9z7OFQ0pyDnLfyZS9Go
8U068qdos9Bku2w8rqkXaXSCuBO2Jtu2P17vA/lHaq9rt4ptpqf+brGJvC3c4J5c532UFy5mlW05
fErtkLRbwH09Rv4meFApLjY5Q3Fg2gufXF32UYaGpWRnmQ4zyGbYPVSWyioTRub1ySkC9AqDef1l
XFuF1O8j+IB+GOPW9RHbScqclzc6foG4rJk/RmZ+wmhXBZipWs5Jq/PZbSMTfwxq809MsHgTHlxV
/ucNbecJOuFxVjpp5gELKt3BDuuNS6JwS17ckSs9GhySvm1wExrNRbnjHSQFvs8rU/MEqdgUGNHK
7VbGxV3PlhL6h9NNQksal992WiEPyHRuxEqTK8G/1WnB6Mk3nSh4BlI9grmLRM1SJJVxb6QMSjmZ
XbjQFqH92VeWbP/vgpniOcTEabWHYcJmkiAW4+68RxEa9rHTIwtwttEhHDoGAUVBqfk1nWjHZuA9
WMH1z45g8KJRaqeVV5Os9p4nilHWMRqXyS82eXwlA7Kj9WJXnS2YwcL1R1V9RxHO2iFkjgVE/iCN
Kvw6EZkcoe1lCa3cmWXdrlxsOjDZIV+JhatT5uqxVR/D4H5EHj4T0tF5FpnHwEI2znm+ttUDoZLq
iBWAS6OkgNslroXKL5G7g7zccQHuANEbm4rbExZyDmILnFjRQ73JnQ72j/Gk6cQX4Hj7c2t8ulP4
V5ybOGJUCkHILNEkQNjWh3SBpCfAmf+OHobDVf9Lsk21oPeyIkyCeyhoY208taV+DYkNW/9wTuht
PLo5CobBSlpWiHtkyspsMG4q26xeU1peJ+AIx+4PF5uZD8SFgpj9iPbsv3EufA8/OQRch+6A8ige
M/Ixq+yQfL+mTc3zHPkFF686eRoUEDd8KSjZEZVsX+8EZXl3GpxWLuVwP42LWAU/U1xGjmxpnGRn
8boqeKiQePf5PVrHfYoNz8qkYuOxKEpOHoH06GV6dTp0V2Nl77vYUIzLMsJfofDt+r9w9/dWpbEb
krhHvJhdHalt5LLon5yEWJO1F6m9wydk6SB55vsJqNpjC7fRxKIzh+HDH6AMB5gVAeQ2a+tXAi0/
ZjQLmncnleOFOfD4st/0xmLIm4bFNRji2MV0DYmpbd+Jc8GolQZwZRswQN9acZye+72RT2Xz3Wjm
yvALlGqHEDWNMzpBnK3j6vySOoH9HhkyFjDvj1GfqCsK30hxAXIkl693zZHamOh0P5nXNK7X/EYE
1grMqLQ3CciZqljUIfGH67Q/rf/TAdlIebUaTprpYqaQU6KZ1H0bV/0t1VewdL3HlAMx/AWrKhUH
wQye0jSBoD/UZ1ivG7fcnjiG20n7jQLIsTzpru20Xo69ZLVVNU31iTpLzr2FzsPoOq2zQ4+a6Cfn
5OKV2qFimEEltGbQIWLdbcXxZJ8trilIZvP+HTIFdc278rj54GfIiwuqSBGUAhYaCyWv77U6i/xs
RC1e2yLrsTdcRAn0kAcyVNvWMNXRUO5H8brJG2xIADFDjpSeB5PbZp0FfJgM2KVOwYy5shoW9GOz
A1vBscJg5rqQ+VCmJErM5W5s5ay7lt/azgQslhjBmnJ3WffA91BKpgGhyp9EEq+Xa6byvxxaNMmL
FiiBT8BMspi9eA9S3Ims7OLyx3TjgIZ9KB5TSia4KrEUiqGsIfgzv6FPe5WBsKCEXzcFliN7uFjf
U3agfF4QEOeS/r9U9fR07GkB/jnQYiGXLx7jHSqpkuswmVZbzsTun0TviCdzqzOi8jHla72X7xsD
ZfoIP7+qlbrAAglRvIjIMMCWzFQULjzpRYq/y7Cski+youIbV3BEUP8xC2GvWS1FfFvtkVlAuvm5
b+HIfwhWw3Subvuw5nO26bpOU6B+2+pANtqRSTTCh807dihAi3GDJlBghEJM9VlRp56vzsvzcfo2
vq9rFE12yvGRrWYcaI+Iz04CVqykkTWt8O4pGQpxFBsODKH5nj5d4MMt8shsGwxh3FcYL6pC+6y4
UJYeCFQpuB/DAlb6NlxBeeqUFByrbIzMXabO8O7GMGFd3VZc2zJ/1Dt/QUPDPRhfpxHpZSZrtrS4
oreOf5aNYBTUZj9ELS+QVgSXrLwn0j4Ip33E453X5x+XyicOgu83sf6h8CY2h2CiDqca8qkWSfQd
FKcumCNLUtWQiCYLNPi2yG9vXHNa+YaeleQTxwE+w21DwUgsUnbA+xendlNncpjofQrrupvpwL67
SvGZOcm8oDDEux7WakqXHBGDNjfq2jfGvqmTY8sTnXL6czzH2vfZWtBJO6aQ3kCWxP3nEIm3lZXs
9Od/qgO3WoWr9MIEqkDtl+Egr7MjJJstTShjR5n3fulELM28Nmcf7HDEXsdSTm2YSXFlr/N6ww46
I+s3TQbHnR0NoF1N1R6jF+nAAE2CjD+rz1pzWd7HQtW/pv91HuRD2PJAqUxmTL78xELEt3xYpywJ
8v98tEYGXsjCPQExbv7WPte0US8dkCDP2Qrb2ZGP6J+7o419MhpvCA+ZUyqaoUYpymZHd4pD1Y16
tTg9P217NTUsq8GPEyj5y28l2YtZYv++2LCK9ltz9Ym4Lu89NFmzlnnUMT7v5YnT6DLjtOQVSMNM
ZQcXh6CoGJz3juGHyhBpUSEoVXC7fPNc8+bdWBjzF8iY0m2ZmfQebV4aL0jm8ewvdT6ubAHqgHma
KTHNKQ+UzBoPR3VevOtKhQ0AmxtQXVA8v3T3oxG003xJ5b2CHy9zpi/G0jqCHCcLLpbmROTHhIBR
CQU6p+GSCXEbTQUP9Wntykgoxfxm6jwqi0Q9AXyrIiE41u0UFrL/xI6mAkll/GvSC9klOWZqE4fR
K4i3FsllFmz6tqcCeyCq6x2BznEcxX0AxONIGLbof5ZxNAXYyxRYz2xk7BS29g4QAF7LuVgn8XNH
VFpSxmAx2sgSLDdCB2KefUJbYvuyAffMf58iEkflh6zTuHtAXifI8a09T94OhDEaoKnz86Pm6EFw
yvS/V8urZUjeh1fNJ4ATGiE5+Ywz9Ch375AdL9N86x6c9Femica9ieU8kjVzHPO/S0ySpGj3UiAa
pBOTqzA3ENIFv/oxJwFS9/SB6BXjRDoAaFS3mMjSygEMhX2ADQDtBl728A5yTH82gcu4+TnuTc3O
dj6pn4+9/KxXZwJvkLx+EFEl3dlR5tv/524++Fv1UUleZuJniN0UkCgOdHJKDrkIZg1BZPnK+067
wo2BwKze0TrV3fuW7MCMZkBUaiPvKpuzK38rggXImDg4Fqw3LBY3rIxv01PxyGdB4BuIfvJDMgO4
Ea2g3aXkA0GhI7zcurQK52iMyzLizYIyiw8wqRslcvlxkuw2p+NNuxtewArOmE/lLs4+R4QqZq3c
lNA7y8/slFcjNTCWooovnqlqbDsDpW2Ed56fUlwA+mP7SE8XPi8Gfl6Jf/THCOxISq9MwWsAciFs
gPcFP4zfp6QBxsi59SrL3A8XIJDtD7YMFEZthIHd/BFEWbghKlceR9yVyWVbhxG/8Ms5zw1czlTb
nt9XXFwVGLhSW9kdx47kKYMguQR3IUi7050R1vhCykG4rGqh8lAcTXFudWvkAmRaMe0KXYXCv9RS
S+7o79Jc6MKKHZj2UImZNX/FzBjLChs5/xzga3OsYZfL2x1txsD9iOgdRKsn5XYAijaWGHesdiSO
Ux//wSHCusPV5nlWmvROC9MbPsj6YphktR0TvrCGOFml5ELZKTsQtbXhNBD3g6RwfgHTBW/W5SoR
z4TQmEBHuYEx5LAvwnraaTnOMTsO8YfXeNVnO3NyrhtBMMA/GBO8rgtZpapyOlVxrl4t/LiGROXi
SBRXmWv6x62r8fr9lBKE5uI7f364DJ0dLapmJ4QaOSW27NUAbydYMwDimdCNNSo/luxU/38VFCZn
NudwZ4/lloSTQgLbo3L3XxM0W6dIy3iRD/NQiv84AzSiuTzy00Em+BFtoOBJoZ99CQfz45N1dVqZ
HRnGxrdTF+w0Vwbr4/eoXrKD23N1qNofkZ3gwjIdkZgt83YCdB9CdTCZpPqvBfTYyrI8uJSmrz2C
xs8h+37glr6QcnxHkNrn4IW+Fr530mWD85encaGAcaHaps9nZsC2KsFrzASA8SpKK8j9X3y2kH3r
caLsvIunYDm8QZXA4UXO++SzGId8e+eGghaIEcDsG3n0qL+FNl3vbLsJ1qiQObfC17RwFmdawJEA
iJ2vasb2RsPBzQvaGFJ3i8qSLyGRlKEn6TS33j9bi6nlhGWthnSTPGpiM6gSL/1Pi4Hr2W3B5X03
m/jFZtId3l659v3mIKXPIJi8p7DRhu3G7J6IoO5Cyyo3jT8zx0Zy+BYqVqilCm8j0LpwPoyzEP6M
lFRJuETyO5668C9SWO6LX2sZ7WI+ceLFK5KqncM6zIrEMtcsl4CTHJKnzuz/l0TCAON/MVub5M3u
KPjWAV6YBi3LRsji3bZO9ptQtZOKxPzv1wrR6ELn2ceKSIxlQ/btoiv+tQMClPHtGzciDuxyicvs
Zrw6pBEUjgw1DZRws/M1i6GSMolwakt7iRBQCNxjmMyfLmz8r/ahWAOuK5GxMGbub+RFMajRMUyY
Pro3o3GgDmQtniyEfSUE+bWrjXHa9pXrB8zZB3JfmXg6yKHqwsjmZlY4u0ysJ8mCFEV80LmH93Sc
qFcPFpVREztJ+gZ1jUx8rTblo3PFJWT/acyic2K7sAj6QbK2gagkLj/J92LJTD8W4y9gT+jDFeRV
M54d5QJr16zR63qL+h/PO2woxT1/h6WCH8MSFByXs/FsF6cDvuP80Y3RTT8ZQzi/MQnROTUyT5bj
CcaDJwT+z9LZdK/cAysjdeoTPcV+q5eCpVlr0vu09GzY8KHQKKpHtOel/ovPu/OTTL4ZtyH+k6KU
K9WbOufv4T9tpoA0HqTxiAhyvJh5TDrI/dyYEtN1AFs9kMzVKk3ND4Be0BGIAjQFoK424z20npTr
swr3ORlk3UaNRi3D2oWbpA/xVp4u67O/hsham/OEBXQbqfoUF4nggIjoJmlqXvwIPkAEL3rlURa+
yh3FqgexPDVr0W+TAYjowseNk9ZZC+bAyjlle2598PlL3jmECgZwvywa9IjG7eCyV2IUwIzngVjM
UTuDpEOvhzLql9zinoVd95HGgVgG1itnigdM9ZqxWbPougsldWXWSZy4DwtzrQyvkZ+KxLviaxuo
/LlbO38R9nPoGgwn3BDjyZFQ+bCeHzqSOHrTi7x3eHn1YZ8U+BjdRTtO0bEKgu/QkSUQhjmR93SS
jLF0AOoRjqeybv/kE9/IxN/Rmhnc6zc6a05H9a7kWGABVlwj9lX2KTb+vJJmWd/lg+XqV9k6BGkV
VameS/Mebca7TUmiGAK49Sj8AlnuSfrPd+HGkur4bfec3C6wD2gwoKPwkye7VyJTuJsq/qgHbqVH
opS+RzhzpeH9pax/S+zW5TVuk26jiJ3Gp2knDkxSZ3EvXEhr+SzHYFu7jAdSYrYii4tsBJdovNoz
bV6tui4aI0naIP7K7GYrUMo4soZWQs/r1ziI9QJtkESRKF7jev1gKX2oQRoVYc/VgF8UtAnUkItt
XtbAH9l+YT6Bhd3hUiygrgOF+psLIxhg9YmaEXFSWiTgdxqd4WjqMwWKUNwbAigM4J+L1T0NnLGt
Q5zBOKZMYPAcSOu/kHk3nEbgwbwa8y7gWMRT/0E9L+761RHZWj83yB+PvTZmr4iNtSqhNh/WXqA0
47rriY6+frnVRGiJfrWkYu0zMx18GJtLaz1nsk+mw0V6dwrjRSkT/q1GsUM7C8P06C1LEeCdC252
9bgxREFXZcG5sjwAhgMsKW5TzhCtg+xJ38qQyJy+a7iSRoAbaXLdUC9LIU+I3x49n348cD4olGEC
UWpH2O86L7bm/yzJsq22uAyMYvVLOTgi7GiCJzIqgZloIRm2wOj2B4GqOfdJTLX+0OQrUhp11gyz
zt6IBPAWHp1o/C3sNB42GDB4z1RtwlClAN++cpjoFSfY39dZSG7lMiq4OUOqVftJO5TBUl+9fm5p
HQJ3sqvLH1QDEHW35dNa/a0wJ5IFHP9zozgdnFkVb5zt7EEBq2IgYc1TLDPx4AeyWI2YZ8rhMXqd
95Qa2ugWxRMxjE9VhDCXrTaZ6VkEmSUu130lF+lYfx3yDU+/ga9wUXMS6SYaUvF/VWWZpcqyrcBd
ZJ9f457dRng0ivB7N7UMtHrDMGRZ9+CJypPRtG/vdXmxJQls94J7EmlKMUAaLEWksQsRr/1KsLQl
/UR98wn/MRJX6AobjORRh/NnffdY4CaOVuu6NMRKeyP/tK8N478JbP4nXzpFgFYAPyuTVHc35Wtx
5yoy4iLswEO4UT6kbRLiqscYCPEK69ixb/FBAW9nPbZgQrYWtpyzE5/hc6s/wFwfzBLFdW+cNrpU
OHJ5SEfn2Adq4ijts936KldwIR8CJ+33Gh2/flDbGnTPDzZVq02cKzhsjkAqOhex3kVactD8FoUB
E5TMgR2JEEASOwys8r4BNpJ78Bnp5psQ6+2DLu2gKUaUp05KQkMwnUWcX6w0rkslD7++/lBe1CBx
/teEhM5IVeEswCDsyzPyGeNh13qlGdT2HNmZsUiCB427NCu4BXB3TFbWBcahmtIffRrUsY20cVOU
fCLq9w/g8U4iiSd8Pf8F5s1CBN4wvAIdZF3/GN53unOnPPjtPLdENxLRSvtleBKy+mA2iyeKV4Tv
MWOaHS0SrWa9dji6+Oa9B+ktzP+JDWWH5KdktVeKCcrrJY0lU98d0RNYaDxmH5CTJAj3NSHur54G
1nbD/XS3dMulzBTcZr7T2Y1R6Xp1/LIDdwFAvVjeZ64S4mdEfdztu7QP+IAfHlXBfBV/gHS+ozku
Eyee/BwgTpvtlngyMJdCx9A8v85PDGT2WLnLskALVL6fN9b2J0mLh6JpN7+LK+Dw6bmpMtAF+5tI
rbIfVYAobqYLZ76hTTfLjK+6a5kVevEVVgRxpdvSEWB1+wFHgqvLLhstlsVfMAXFxDtdLKGrfLq1
GyvJOuinLesnYwoS0AyioeNrCF5y41++1WzgefeZb//N7AS/MTWPkqCtfR2gp3NorZq7RXZpjZTF
qs0ftWT8zWMakHmQM39QqiNjSCWmt0jXqNtZGjJp/GPAKqiFvTjoNxAQsG5p6Uq/GFA80vIAYyVi
TqiHaG0NSJ05tBW6i+v78sNTuoX4bUP+KfRxsBBH6rjrZZA0NUbytKmgMUmdPclZhSN4cFfI4r3G
jEiaUp7nMmSe3l0f1zo14cHk27dGIkHoShfRjJrkASbTOMymhhJW14TG49mwHUWELlHdKxI2mhJC
I3iZAd58FkgV4XKgiam6sTuBAA5y+7d5TsZJS/KMIBnR+YS0RjQi+slk0ohXoIvohWDffoPYBVcF
lnKWvQ65X6IbfB74wEnXXEaz2EaYPttRyFMf86J9Ly9I5W4xA+8pVsFeg5JS7jnVjaJ2Bgfyw7rv
X1UZBn+MQCLli/tTwVwty1Pyn/mu1iJ1rfYKyA7FxeyFaGVr9hKMCebZS8aY7G7rOXRDTmGy0Sw8
wjM2lIyGedbfscXbW5/oRKn083iXRFJoLy4VbX8MzMyfdyFCVviiLj1hd/Bi/Ho8+bI31mYjI1mn
jEM0mB26GaNsAtZAXuhEu07t+wiO+QnJHUw/sfnblcCPy9T640MBswV9gKIDbhknbCcEV8hWUl58
NWiwXgksNAQvrmMXXGtccJVI87vFcK1+X+MjFT0kMc6yGPhOpxlYlGDLD4KEQwexH4gV8b0AS0NY
T+KUwylrn86Mxh6Iw6OIRhkgzFGsbE9idfCMuSwyqkZtx5PNZ0eqSY0aOlywvTlxeb51AZhSnCT6
UzZrwaPwHzmkB5XkHlwaH8fzfCJAOqByLUBSCPpkJObGhh54Q08QLn6XC73KA2BQagg8B57lotEj
cw3Ow8WeXKd7oqm5NtqfzYQsiY8nztIZzRCV3JOdBvgIfOngDIGrwqwHCx3YJPWkWhZmCweC6H33
QKNCwisZC4vI6bhCBC17zVHnqM7o3WKYcn+svcsqvhzQXS54oGBuFlOx6GdIz+VlRd2KLgRkZDr/
QtOvK1su2nlKbkGt6q1z/W7805uw6r5aV5eogub2b+AUjchfzycMHnQpXYL4rY6XNq6tI5xSmgzs
vSJPQRbr1+e39S+lJJlvdpl4ho5ETE2p/FgrEACSnlMLGL4It32w2IxXEhOvkqtXC5i/ZbgUQfFf
gShdslxEj60sHkG20RKQaSbYR8aZNaKs9gSNV7rbDtove83eJWl6MksUu/MmxYMmMWwE6E1UlBqr
DYOBqIx4P3VTZ2SKbXIsFtBnwN/cI1F6QlqoAp5zqpCtg2oVidapXD8Ff4zYItyy0jB/3U+oAjeZ
ipak62o5WesmV5haJIeUHWZB+Xmvwln7kJ504N3cKodsBmMSMPG9xkTJrH1j+0BgF2+1tHgCtIw5
Sj/yrvR2hVD9IY82E/pQxP69kPht5RVbRI6hy+7WBDak+DyIkb/hR2+Ld6BdhqdZyJq3RvHyd8Ga
aZYvkKBtZtS3Ten6UFUXaBJRwroPu7bQYfkwDqMtg3WYzbnILMgAeWM22AhhOVIPS/mf15iF+KFt
xaPgdJ4uevOl0vJl1W1bVDRzfEFBC8T6XZ4kIfo65PQ/WneN21UQcs5kqnogbf5hxHPlrHDpaBwP
51cBLnASqmQmbw7FXoVBYSTGaiBf/GEYUodt7fAra/2qXWIGVIqW+q1566igWuxFOtCE6/6L46Gn
b1TZ3WrkAjrWeFP30LZDkjhr6FA7rQHvbH/4rzeWZTN4WEtqt0PrBi8PD2c/zOMrxtWLN5u2SN/Q
OQVZvsRRlkfZkJ48UKAZNmMoTrXhNFM/TgKVjSdEkwDg4WebProVxuqHevkbTFP4b0dDyFCH/z1C
bpgUeyeXUIDFmg/NMLoCllgIMJTMGDneIBPV0eYnXKc3TbeIJ0xf/KOjNIEFh7DUuCQZcRQqX+Po
NYty2u1nUHYAzojt6dS75oNpA9+p6wuR2+N+UkVUcurGO7KAr99UlUDWZj14dC3ICDzPGsP5a7+w
jY34GoXTNH9RDk0se5rwv8ZKFglcxjYbDFe67hmuuoeeIh3HNSGB+/tl7tyh+yXf0hyXE6rWOkeL
6f9pF52Abq1JexUAXIUdi0POmTW6uyUYP7kTKMfzWhAMIIuH/NMQy1VX7JfYf2WK9riDvshhI356
5HK/V/uN3vFeVq9H2ZxmbcixskRMIwKKzUWcyri6qNM9fqUtbq4QqH/ZGXCLWXW+VCSJloilWzcH
3PcNJkiiZgv9nusLWgD9i58gK8TNWOJ46B5dV38Drm9brKdX/QowkAsubBOkr9Mywe3KrAggo+EF
c+Hj/UaEI31CGlwHQrD92UIQmD2Se0iljy63LoRIJkjOQeKJKJNuPZIgaL/5SohY9vOcPFEcLTjR
4QUgmigt5SnfkJjuc3df3gxuMEg1zc95+emDldUHk3ZkZBF4mQNEUM02hCrOphxA4zpE2R10E8Yd
MhSL2Vc4Onb7+DPTaTURjpyqO32jeUTnbeU8hI6O1FEkocTjdvNko9ozVBCjliOCnMs8QMkJZj1w
4pkT9+D4epw+Ds9g6jgZbvE/4+d32h5riwfHxrEZ7o1Gc9KY/txyiqyGbgKnd65ttbJBs569B2v7
BiHGppVQ+PLMYqRpMBMq+1rUDlNVt8vWI9vnOgyN5Io4Mo+a2XoACsQU3j9Vqp0H2p171M2N1Qbu
hU0qQdEGHcW+dmPNwTMpMzFmB3dF3FvomS77HVRDh0XKkOGhOyDRgLMyR1TROY+dYHJ4caSzyCik
e6YYOCKuxecTx4guHx0HUY2zeBcE4zU0tXidyftaFEzbufjYqyVhvqk84FAb6i6yXLZAeHLsNMpJ
n6mTpwcQkPnt3odDgchtI6MafSavwBDlDeXKMSZGpgDXSp7ZoQfiDuDH4Dtz4Ymd+wxO6BpEXNkM
zPlCskq+Av+BVqr3LqTAHbD4KJwlDeh2x4xSJCAKsenR3rzunv77YVd1wCfE3qm9QZTZf4zUoJbW
eZD11iWg/9irZ3M3hdupxCVgMzWFdOeUMcxrE8EjPREUSCsQA1Aj4ZOMmGa4gKZhalhG1IRtjYTb
CZSh1Mqka0/7Z8u1Lg+WnsPUlUT1qceIdlEAE0tK/vTZ1bd5L+cOY8iuJj0Y7JjL/pB5CLVR3r/N
oZDPziXuQpophC6m5e7OpRTD/CZrnbMgnd+Dnlzfh5/k9xyOE2gNrcc6HpgkLcD0SDCpGdNSWOO+
kYyzH6WeXU9r6kZLrZcQ7JC9j39t8FUg/9Tmw15uVjIxpJMWC7HmgGLvhf2oQGd1sgFXUL4GtLtn
/1TJTG8ObzH9aPaBdfYvDaa03iZ893SkUItMs+xFSIiNahtEAN2N9vPi6j5/qRQ217sN9ctUxvCz
Kmz8d8CKhCwDkJVgr7/IDejGpDX94rVkNiEQduAIWpq1DkWmAiLXL0KisrRAi8J6fdewcEwgPQMo
DOUskehzmeGQItNdrzUfkfHH2AxNVT644ho/phkWXBdv1rsMS1sHYY1lBePqf3UdEX+6t0DesIn7
4MtWkxQbwj7i4jFDPNBIIJgJgQQiGBG1jGBbDvozhJ+ndxrodYkvNTa2TkFykz+SjtC+senxR9TL
Rzf6gcrnRCNDPDobTv9oXT7AQ09aBxfPUAxEGonKKaoJtv+GelKr2RK/3TGJpnRuf6ZhIiOP/h51
zDR7TAL2N0b+59Tv+38Cg9Oc16EuIB77RY7tVg+CImVGOQ0M77wms2sjiL9A/WXLOnPNWBnLZv/w
3zCZ6xrXX+hmx91HH05B/cBAVXMH4ercLNB5U+4iUmiVYtFiGYj5XzLezYFBBvVWPwp1F/lCXgjR
7FmadnVxvDO+ZE69Qfqqd4EN/90B5N7uGx+Ie+i35NSFFqkHi+65MGa2BmN4MWff0enEO2nn66aP
RM94XMmOKQXpgXUvDdTeEaD19JckG5i11YAE8+BgkgcvZQ3Q+47evsip28V36701B1gPKx5OAgTM
pFK9cUi4XLy5Dbp7vfQHeHVlQT8Tl/QeoD+iH187Xze+OIbJfGGewr4CPlkGFzKcsVBrbrhnRsH2
RCML19DVcritRwmivFP3aPy49cDNv62P0rqrFW90qrx2mcyec6vw8uRUktHAi08wbPDFehzD70UO
lZIHVfouUYL3Iy6JqY8K2gfPfjD9vj6iCjxPSU2QgArZLA/8fDnZAJtyLZ8CUl5nC2WQsMnzcl/v
ZZ9RSkYC8/O+qSPWwIrg8XKvFON607pRfBjSP62zCcODu0d4MxzONT80W8hm7z1mmLvqNxFoDdZP
dpWWuopN+LLQZDmajEROJgZjlwOSX59ld+VipclC3NEHNp2hrNzX4VblbQJ7stLJUAkB1t/BtPdy
HjSCLMriD1pS69j9CLLRDa8Ji7FpHbDceTuh9HtT/xFBTitZaXJns1u6/I+oHnrDdOBPe91E5aVZ
1dgmjsheEfp9we/LfIqU/X49HgSOjapwmqr5LJAb84781ViZvWDjhjz+EdzQIYISffwelDzJ2nWI
YGcFm3uYICHezcImhedXT9fymr3bbwUewIRuKZnx5hE58wDos0XgsbRTBJ+8Vf9nPFEba4H677YJ
IQr+wtWy57wI9ZKG2cGXBm8JRCTtm1b+WEfDR+x/EMY47cK6o3EZ1EUbS8ehXyaGGwwq8SZb6Y7O
FphYQwHprwo9U6lUgPKg0hHm/+RhaJwDb5UtEUnB84MtXQ1gIxUFSfPpK+mYS46pWqPsHCR2oQIb
kYwTcnopTtoXdpIsUNPWA2nZHwTgcf3dW4g3MIQPMKTkaIb9ILtepbb21Qj3NqlGUDa8btl+kKCD
4CUEsyre6bgzZhwz2/yMQWqlPSkmM/JcOgpcT5ee7r+DW0osveqUNvPHL6yqR0trh8tV0dUyFiMT
eV795CDCgDRtcfPo5Tj4BKjCvNrUMVcP5jMyf9VZAvmMArvLsmAzwYM9s32Av1XpGEliP5bB2kd7
r+6GLGIBU8HwzEJYII4mblYxd2MKQkxE+eshQWzbli8aKWr0LXdFzAYaHxr54OH0rV8e+mSZZxfu
8VkXSTV0a0b4u/mi0BoIEjoS6w742zoPcL69Ftk9w4iZKA0NbmN5/Gf+xxV81nOun66gE4aQ0YkT
/eO64e6PhiBHbfY0CY5bBy8fFWWCQFzsec4uSnyV5O/GuAe0jJ2kexH7DTN+wftihRkBBoPWaTnZ
wyh8IXGlcQTL+D35PN0jSVHT2h6OMRnecSREyD8sayqYKfa1MGHSds0sY/DdqyvIayiLSQxpHis2
b2ztkwWq4ccIfOrfAdtJWl4RIJP+NWKkpJcyZGi9CnydZrid/qRPklOiHMgGpiBkwD6qZoSS/83k
4RWXIWTflLRw5BxHIPa3bzKpYe7VrUd4KjdSjQFJpEKeOQ6TavZPRKhdZ2Uo8UhFnYGrAYOzzopo
+PEcOQUZCY6HN46lcpWT0EniW2VKgLiTSZkNwnNwozKkXkFM/UVpRxPh+Dseql+SXc2/+NiXx+Nx
bhlB6SEC6Tv0o8vPVLLg8JYzCwTGccSRch8xRdqIA96nTi8XlfVn9D8AazNR2fnFdOBBqJP30FGw
Tx+nktMEKyopK3Di830vOLXmbPtf9dQ0sYINfq/1qBF9cSYKOoQrmzGh6wpXsFzH1TdaaBFFD6dB
Bd6wKohO46eCnMxYMQOwBEQ2UESWhf/HtkApcvRjhYQkY2vY0QRfuDSqPhrnhrL1TXonAGZ3B91W
8849L626qZKrQjeNk5aXmDeePWGCzh04u9HFoQUq1Dm2tXDOD57B/Z09nsgDDL0PEJEtRunu8SBy
/Sf9D6vCKcZa+Kl4sVhg7/65jAeU6dt3mNDTmhgBuVyU9j9zqTDsKLt+/P45TJb3F6P7KSDHEukC
0d8tLMk28x/+8ZV6o2IRFvT34ZLYJdp/tEqNsgWxyXoLt30i1UlWi3P2HQMXzV1zqePgYQvRclfu
o74LBNmJKcZ1yytfGdax67hcBqg2CyS3PNwAhlgw7Fvg1zxp6UEkDppSVGH77JbcnsuMa+yvP3ty
18MWGa+/cWQc6XDoMKsulnAAVxZ+iY4QPGSbUKmw56LkPzCFKiokCTRkB3LV1xR/0Av/DqeP9PtN
l7tpbkqs+AxtxP5kvF+5EWQIWVBtDAZFzob+h+Hq4nLA8EqMV2XruP2lb/OmqpimQKaMLcrPL/23
BPCGvbRcfAGsTBbFAr8TX3r20ZBm+bHTStVkggogTESQuKJ0yrL2YV8WjA6DxB2IaK1wZeLSCHti
m5OFRCADdKTDGRA9ncEW5BrOJ7O2t0y/IJq3M4WEgRs958ATwEKw1xHl6ISSKD11DQFAuHbfxMsR
QAglCCOmNtI75z2WJ+D2GGLc/gPgDzCaTLH5/ERfRFYrXkR7xMgd8JMUtogDnKW8HPdRePt4VXWZ
/2RFXYbgJKuiF4bSmD9M9R/cjx4AertmCa31PGC7KrUC0sUSWDaCGbNbeR21suNaiKnVtI68EEtV
lFL2lNVsLvXMjcpUAbm2eVWPsUWzwClF1oQhbHmNsv7Dt+QEivrPJJp1ko5XG61I6IkI6PEpbbfe
pLINa6qwlbTtf6OMjmJr5Rgvr58sniZmjtjWRlFGeNebOtRma0puvFF5KTBLJvzUsDXkyyaQL17j
EW+sQ2mHN15icA9CxxXy5Jcg/PGeI1X/pPWMVLIqtrlLMUse/c/Flf8NfmKpY8ICQ2iOXC9F7Wdp
WXkH1FYaguiOC1kgpF4dwfuCC7O16ukwV7bMH2vtRZI8BnRDO9k8uzSXaLokkLWty6/7gRNIuqrG
zdK1eBBa+Mt1WbdKOy23sIN7HcJHDCqnUW2YyL2hb+bwpjm9N7hssvBXreY9UpUeibK3pLPGghjV
qyXNE1bzinGhSDJmp9+MiCXozlKZITTJITmH6+G4ZIvvl3Ay+ZVj5QjJu5/ZIxMEUgDSIzoXcDJ/
vp/KBpDX/qwoZ2836i1Z8iPROZ/hm0UByj4PT0W64UkMRW/S1SBU9/V8m7pZOerTvx701V84pf3v
s83895lmcI5Qqylx3zqJyRu/TryppzFwvxdHYrFrOJoV5YFwhvmCZQ844t2lUVF+iJ2NOt1eLE0Q
zKfk9WFRDxKfU3uhQliFwUK1dOKj3oPgdUf5uqitdfIqYPwNfW/a6nibBMe0471AmKE4Fn7yyLdt
pGFLr8drfKvZIA7gaGyZmL/GQq6Zteo5UGHzZ+9URF614oxDm8GREgi9ymPmUz/oysckSsZrmHY3
/bgz+RQCFmKgdWv6zojfmXj8jlSfJQQfEfEsjyNl/DXK5bWdQEX+Zo0MXMkLmdNtMKkFdM376/zX
5Xu7MbXzbld6PU7O5KZ9f2Siz8nnU8Y8o+khJwk0Q/5mZ0H1NQ6KGVqhc2qnp65V+MDcrLyTFJoj
e1v5BHp7rS0JXmJp6lyh35ifvZwCAMMqvG9ZThmxTu6izhT6FAxNpXxOCcw/MA+AstA8XFrGcWAR
dcyb6urVsNyrOAGQAHgDZNJgLTUq3kXbPTZxpOOL86qd6CWl8BzMP1B+I2Cy7qmyjnh7h2vGWzYo
EXqopjSSNvRfDrmWjW5Fzui3k3dQ2OBJhWxlBJSQOPWufM2e4411KSosGCWXM3jDRomgCmYic2sg
1z5tCgxRMneoTv8ALVOLeT9SJU+X/7OMIGTMLDAqMwXMxsA/lkktOh/6iv9aG5NNpXhKnPFWfzoD
O150d54CqxXcWPawpM+kpZwWXYjbTnXu6Bdfox5zdpK6vcjFZdt7lR1HEQfqpb6WF5xR180z6hR+
mYaQH/NkOCZQe57RRqXVsra5IUZ22i38uUfnM/ySnodd5awpSpJuq86CQqWRCY1anIUjAeGETNVj
ntZ99wbbrC7BSCchqGSXzKOdL6w3GbM7DgJiAkRbHwDKujxeiy9onYQRS9A44geb014hzqCW4NDq
IN4E8Vt4851ks9XXk7N1lXXGsYswh4tlzcm9ItwnXrLvVqYmi/hpYhUr1PJXphy6KOvYy9SOVrtX
zIhQKucTqUkR2C21YeoHgwXoKoYbxzZ7aVAvcmZu+J/MvHGxqUahpOKowpQh1EhticW5ZuOegBWK
r2vCOvdwZgd9IDZmhWyhB/QovCPqwJGNhyDjp2FGLgOxDQxQELBNlcPbpW7CwogmYzO1JWYEdsas
kvZvhyvIAad4LTmcPeWvdD7HIveylQIa4V2ln+IGSlYxY/LcMLdG/ygLvz4nDKvtTRYmkX6VHk8r
nLHBzuQ8JdunPCcFnwNDFjxoNGQwW9J4rG75WvombW/Xi8aCxK1J+E+yE8Hzy+IMpeli+Vs2UA0Q
idPfK/fKP9QRqlulo/IfkFAKERv6owVe7huwqMZXJUqKvs1aC/Nn2DCz4mRPd/6hXoYzsOuQDP6x
5ldugBtMbSvqbYXC6VhJcuVXAjMKEVK8kAoglv+sd4fx0ES9abCELJpDcCIY3GYBj/He1fKN2z2E
AMph4ZHuY782PAn9fcLKR4lFF+nva2P0NgCL/NBIWb+kf/55Sl1xwndkxrEBCm7U+seF8wzs1QAC
YP6kztQGlHLAmNXA4Y1/WPJR3ssZaOzLyZFAQgi9031qfgjjVkKj+OfhWOxE7lzRYqoZa4c6BGZH
Ul804lHmzxLzGatuSfGeuCN33b+dKO926KvW6m0nK9xe48wYgjt/IoCikTj5x+o51NmgS+tHNnCT
V28M9ty3l5bhoIGjHwE3r2LC6s2ZUxVAViNqK/vbZQ2wqz7xXelukz/clQzmt+cLp62ExGxFz49z
3wvHbZ25An2H9mTYh6rrOasDX6tcCapYYiUsDjXHNPkDkSE2mTEvEO3ttwJO4T0r9CQQKc14pQUs
2W1rbFCIEFfuctzinpMgEE7tE0yUP2CWx4evpnh4FeL4jdSMNyJNmhsAXecpc/EP/IakPpIauQTV
CUCSA8C2z9WeE66TJMrORXD8eHu1zlcNZkOBUGj98XeQFUMj2cz0aUJtWUjciiUNllaV2mfBB3E+
Jax3V6gsTOi85Jp0mhGvzqhoqGimtlueczZ90Ilaob7zO0+FXPuHXTvm+H7UAmMD3HIjZEOrrD1Z
iT2BnUZqDNrdDm5PV3JDClr+zTnJ9Ku6QKuVmggG0/gd62PSMaRdw+xawqvvQMQ2sw/lfsjRmKO8
vbYWBbvTm2wOvb/n2OZ+Q45VNVPJi6Zlvn6dzydd7/YyQHojvAzK9oOeoiJfwMC1MXlS6u/YfTyt
anWkdgxwts9C46OhL6ZdpOJr4ZE03qhkbLbjuZXmJ9mpu7ebjXKjjWILro8TScyRTEM32XkcV1nk
5ByGo7bWCz1GnwJjgrr3btLN/lxwgi928DfxhX0b22YY8I4zvwHCmzvRw4lr6Ofj50SYsgResSgQ
5/7jUyGnw8Ewjy2xffAqAoy1NqElkTEtH4Xep1tg+W9nB/0jXzA1+vLBCB3PDlIK9D2uKEakHxNc
a5pB4trpkE2jW+9d8ZFMso9R3Jsiz/QReUp9tZB24f8nOpRysQlAC8ooKQs5ZjIvG36jt80eqoSa
tkjYSMn+cs6SJNYeTWS2r18uzC6d38vX2sQIDHTLc/u688OKgzpn9JUHC0GryLCWiL+BPQ9Z3fI4
bopApYHnfvKkaOdKqdmKM+v2x/XaaAxg2h2u9RbK6Piag61486N/XJ+Pwt9p7Gaet3g1RRZ+PpPX
mhQw4i6QQyf4zmKol8rroa1WdPd6L2d7O/zJTAekyZCIurRiV6imctjf0y4BdXGD1FXxGeGa1MCo
akoIT2Ucc2gCl6NU4qhtUCtgrD4a8YzJh5oTt8yoOkBvP9whOutfyqo/uF8FO6XPNxBAbZaLn1uY
y/514IW5t6glo8N7/riEGqMjhCha0mpn5p8bVIwMIMNH/oYlX5Q6M4rurWNFgt4K9rbMkL81tEOu
6XBe36gcTKMJ8Y+yCoi52J5UJy6k1uPAQ95Mc0AgCUA2J0P4inHCMnzUq3WMFvcs9aM8+/RbPVyR
EX5BMj0HfOMJdf8cvJCXJcGp+VZjiRmK5PUtjO3MhZsabxFJlotp8UCPK/1tDw3oQsF9HWqEpV8n
3dVKaxPep0z3Lx9X+rLeELc4fbyg9fwpBJO4bSC7wrz45sl85Ec+sErkzThIME/jifkktBp+/d49
iGNbfBwTPWhHnPy5eNBqXKCOHliiQHQISL7kJmMfH2xYNbnb8lZp9+fZ9OWghWF+vhu4t0EbaKdm
4GEHv2wY/A0tamWhScUY9CmB4ar7wgu8qkCxPE9KCEEVdElV56KKxvD+d0zzzrEPYTEAFzDJ9zV9
wOX650Gr6OsJ1CwY6O5kGvaNjAxX5PKWbNdwdS5HGQSkAsIvHUCw8I84NQuMAWJdQWRvJBeeuJQd
F+wmsTcy+l/RjhCvR1ydwlZwzC1zRsoSgbMd7HDbvjsfdW9zxA9WptziHFhaQc0yBmVS7cnCTSiU
SS29884qO3mDv8Fwdze4e7U3N5GtgRyfnqEF0BZS0V0Xqn0MgnuQ4ni1P/NQMDF7MoVOs7/Qi9bS
vxY/wpS/mTmsxQ+6j8tY4FC1L7iSf4db9PNSBK4jUMAtO/PZq4Twc9IcOOwluoErbxqi7SQG90fS
/uvYKG+ZkDZnCwlzw/xmue4871QUGui6sa/wYHSOtXOjExiQ/2CT04cm9JcUF8Up1EW+JpEVB/Nd
qXS6XlDxfTx78EDMjqsppThihPF7EAklU8OWGzD3D0Q0J3Zwn3TIOohDL8TaOOhG161J6Z6FCmq+
uk6v5QDvEJTV40qlptCygy39eKax1u6Mm4tKRW0I4X7NQ57YSETk13xbzGgdTtb5gvOnak+sZloa
+ZTCuEVA1OoFBLSyFlIdM0/DzORTtYyC7vDqvqXHztJFYBoWMkGlxDORWv14TX0shYjtIMaNy2Kz
wnDXi7Xr1EWoHFP2xxGiRk1u65n/F4T3XKEKcQORmsorQpz6fLteMm1vmbmrK1CEuAdvum0HeLTd
14UgHSZcoqXQc3OM4ND5hHDvnOcXZcf3FKScJKD+YpAxcJ9hFocrWZprXDjxbS+G7+G5CHeNh+51
LtITfSAiJyMOjkG23fNUV/c2oTrII33lOL85GLZ2S+f1OmNFVvX++vTjbW/vDtpT8LlEjkbUCWEe
DxldD9JLd1/QZoUNhyp4eHalvi6ljHNW/7Ad+AH3wUrVOx8PcZQN1sPbgnPr5BHY5rWsC33iNV25
HgN2OsT9nvFWp+AVWm717iVxHKsXO0YRrTM9yuRCPcAHLAUxx5FH8n/q7ISmvT+HbISRQyPQK6Ko
J0IvouTuQyi96DDfFB7o0Ft5ejSuUmV8gpsB5bQsfPaEmH8WveDzZt4bvJKZSuzyZtRVe2RIVlAQ
UvMI+MXuNr5a49+b6KbL5+TNcFFAV4YTGXDp3EzZqPc6nMI7hTlEvR05TMVRu2u4rQ+LJM0Ns3tm
t9VpPC89if6mvv8KBi0QSsTfepFGAWzgDfQudOMKGbFfnJFk/1Js/3/ZjmflhN05k2MtWrsjX2Fj
/FNi5RDb/ORrOi3dmEbXc5Ub0BVg0krRgA0C2EIDhqrt/kQ8kyJgSaaLJylYJxFpQlvh2J2paOUX
eXGTj58k0x84osIcTi3oRmeg4fCKigVBDIfOIhCMQlPnmmOE/4xYiZ4Uq1/B/fS5D/WgM0o4C0WI
USVwUZjoB8l13Kq3nIAmzYtcMuc9Md6YRhqpqytkfPAxcYCA3jJl8kN28Xk0XCiC/DOTEuj6dlmV
eNiNolEy7VJRxZQ23wppYiqmHjGSoED12iANSKtL0nek0qY9eOIGBQgjk6q2r6OvxbeSFEJXatJt
sqLjiz/Nk7HKabZlU8slZPQxANEkAZUj/FQiFDS+Z9luMiQ0OQq4JpFELKLfI0ohSg+LJBDR9OLE
HOYxspPSVhC8eU0Tqxshb7okn9fotyaBdedo9HdWyYEkCPhYIGiir2pNJzMVwjPMfKkjctGtcJlU
Xa0XBfOBLLEt3+R2rP+4kD6TWyYWSJhKXzbOJ147YL/DYYNJmYm5s6otjwkBd+NSANc7Qa6/LPKI
yTn0ozmByxxwK240NewS+ZhusDH2TMNvcm6/bhDzHN2c/tiX1FVxBKLspK7fk5sM5c9jm/L29yOz
f+QkC8dNctE1cDECL4OkXOmcy21GQl5LzSaxP56/AQAdtLR+VZ/QTQsrcTbkcXcx2mZbIS09cdgR
IjjnoL+8u9mY2Q0xXMrmjdE/Mc6JYiGRe1AhnV2e0urbEIyHZJy9rqoBqItk5e9FRw54JVj8MeUr
O0wCMwNVviGz8vnrUtbh7lCBj8kSM3hO0sx1QgSPwx8sgOAYfi7pKANZcW88cvGJLxgCS42xcOZa
oN4ecR6gkxbfWB/H2UWumsUEmk0KW8SIeq1x9ZmoA9fobA3vh06QEp7vBoqf4xwYq/osocv6X5VZ
84rwC0WJg7Pk2naIGtYn/g5fmll0/FdVyDqB5aK8wQrOMvRv4yD2vaJ0RqLz97ULKCl5NZYQvxXL
r/yAGflEMnRIRZVKzNZ6QYmC0QjNQ53Xb11gkmKA2UsB0cD+OmgDsZYvByzmE4gubXwWgeSQ5B3s
G15fgTcGs5Sm/Kw7NLKFtZSnHtVk0CYW2GsKMtDFLwuGpcJXvIBIMdbWC0deIKAihaeuFZIW/4C8
RAy5ghHelCRhBXOqhWl6RKYemDNOOrwtz81KyS5QM2V0BwtNa+9LktoIEM+tWTZ1KoRHztviHGNF
7BrZD8OafY04R5UFlkrpiUHT0IFNqbrwWq3kpcu5T6t/96Wkk0YeKTv9bIkPK92e7j+/E2vJsae/
TjtemyS/WjKF+LAcv+l9WhkZfd+Cf9f/lf0cu69wsKFGN/xUup3TNfQ5DNuP598Z86xaJtSoFhGv
rcacEQlnM6IIbdabZFrLDOAINUFi1OjWyO7Xr2KfbWW8el95HQDriiXzTViT8HJ9NkKKA0hNh7Q3
EejfEYumMwjFxVze9UuE8GCIhY7HQtrTEyMHdGxFqMKXTrub+3za79f0Lz72YrBoMa0TgFg+RRxS
7elRJbTAt9Pjjh+Mzjjyd9E9IdnneKkme81UAVo5ICu6SFpT9Tm6pHtS4hL2TdRoyVHgym0Uuaj+
lmWCXrZyUwKmuwQntqhfGdZ43Zumk+AWdGkS6P9bQxTdYIUNwJYWMt3JMmmPNjrokNNamXxu1Is8
MslwG0mr4S3Cc9yYSP5cNNjwMlTnWjJHnwt8TwdP3GowRTfTRExlbYOXZa/x1FY0+l6My/fSjcF8
TB5z8NNnp3ULooxHdCdP75db2mLM2TmEnsadQGHOCfdzoAv9bE/8BwqRhWizo+MI51w0MJ9tBFQA
xOIVseJZtRbjtrFwfQP/Zh1wNhzbQ2AvDoK9lfeB3bsduidFNEglBEEK7V6WoBzpN1MmmqK+21VK
EYsW2n7mkXOAgPqM80FePpeoOi+6LOQIgZoceoldtK5uvoopyTDdvSQLVBA1LjXjvwaOKZytyiSi
edayyzbuMQJZTZJdfMSjkx1eysAZxVJMeJV6mpVRQlulPzc1ZK2K/CoxfPq924KCUmJkeW8DQURq
gLD38vpNKT8D6YsCx6AAqwQZWvAy+K6xiAiSazTeFN2H7oi81jNmLGuLWnlbvfuhKIerbdGgmoJx
LgXYECvkeQNOWA/eHdzMgxvSnMMH0u/5/oa8XJVliWHfbENf00Zr2/lphlVOoIFIM4DRC/O6toqu
lyIXrcpLG4SetvZ4bDkkvEHzgZ1mxG4PBh5hlGIDdDNMghCmSrTREdIINpBOzPyiHVP4IsUm92zj
q6E6swWLaLMM+GOT/ZMW10h54yR77AUo7/Kjk3V+YYue43UZtkPePS3svBJvyyyo7y3mMFoqkwRQ
yujJ6oxth5daLWocJzkK6m1S5FXhPsFZEjR/DHShtJtnKGShlZ3ipWNYPmJXVpXHpCbPMFxAvs+T
F/FzIYQ4rgSPn4azTUZUd7NOGf4s5BoVOR1pxGufLlJDirfPsmiVHILnsE5q6pCKGYXzFVxmIcgC
8rzoMsrn8i/dqvYCZpNtgubGWdPvV/86U2j2OLC40UILq9IKV+E6SyK2bmngKKMq5CHT9iSgg1dT
lQtVYWqWpU+6p25oxP/BniniXENDQ1/ZKXLyJcsuZHC9OLJ8pXOp0RRS92CMupn/5AeIAOS+X10t
anZUw6uNi5PX8jnZxb2l3aTX1S/Li5ryl7MVDmZGYv63pR42+3D5lUHzXHC8gEBBW7sElsti9Fcr
j6PbvVTz3HNfBlYDUggisk/REP7yP0QX81F0ScOiPUlL2K6m+abEEDmO1WUvHtNXD6bjFsZv0oNi
/Ufa1ciBgGNHVOPLQI2IEzd+esHsm0Gvz/P7ptNBgHlwUf6yH0O2hqcPE590ozP2mhBgdIIIXnJC
hdLRpz0HIoYwOpFc9YHQRsi0rbojT1QtULDADbge8mpQk7PQS84Zl8fpDa1ZYLKVr/AJZgwHpcwR
GAs6sR2R7fcBJAjfhOPDphgh/RNSAtmWu3stTwk1UEMvhmugHyTiK9SDQY6Kpgp+4uk3VK5jNqlq
wCYu84EpFxZm3PDNFi7QoH4CBhZ4oAY3qdi90EQSUQiNPn8jGAYW8PHkIfK9wDBf5NGkUueSEzCD
16gWpe45VwOKNz4/e+f+fpx3fRe6u8SJTMomte23iDK/B0kFnudPLxHyf/At/7TDV2+/ba51jJem
R+YEcuxDeCJCSG9QJ43FKdq8ZGjiJWjNP9hvNCrGqHwBsyQLly1ONniCKC7wU389vzczrxewJPCJ
setBipRuMwaLOJ0u93bFpG5XykdbODFd3OCJayCvb0GJeezetQgT6sHJSKgdh34S+amgvQoaiHfS
JTbrCboDtg8j9i/2MsOJ1N65JjHOk2iM3rOSnT/5C6Bv4WCPeiuZqpsrJMG9h3K2o+Gc9TvyBpor
vqLWk9XQd9LM1tw5C3bLEADPA2ccpOGXqmB/Yd0bde71Z7Riwzh7Ql/iacayOGPXFwgj/N93aU7F
mIBZhd2JwiT0MxY3t+7ejHpRymnaFbZiOgp3ahuOzwH8F6YznQNeAFCvZ69SqgFgaY3WL/pECuZi
J/ikcxA13yKHNyX/B0y4NTnwKOg97xYv2C2QhMugeaClC6McwxCe1BdwO4ibLDRvQ/MRoMLqZakm
mGm2D7p4yBSyN23uoEJBh/KiebWyYlAFmNzamCh+nQjhWKrSuftQz3DZQ/Lv+qxkjaISgrnmk6sE
C3HUgLvOY9JfA9ahUIHbBRY03qnlvozIIBIuKIu1mDhQZQ4TwL4ytQZWT8XgHetftE2b5sn+GeeF
AxFFiGgf+Wqpw0XOaHXmuKyvATFWOK6D/Ug1L8+yZ173kWrnCHJ0qBA6VMDKzqns3vW3VybEbItC
euKSIWulHnvugaG5nDbm+NkZIUw16XQh1pUbVM1bP6F+2Qi6thkSVG6kiKO26IpvUUeZVPXZ+M1Y
jXCEuxm/x5Ib6wYOESYPloIyKomb800NV2voFj2wEAkHqvO7y1OBAq9ipSGSd8kRdjlceRQ9xXAb
wK4ZY2efqAMA3nRyLQak8RS4f+lmxLfm6codDNUv87N0hmZtPY7f8oJcHqqttrG4OMv7d1SZZqOg
bvs9kscNV/oR+b/MousCVn2Rwm0QDrgWkaWTBjUw+qC52EVePIGFUyhOE4VH3Eu77MYuNPDmNIHn
pnazSULifa9yfu6H7SrB9XoCnveo9b/zf6MjtBf+RNk+wmU03hwhnlk2XrTROrE5y6Y7XlYC+3lQ
UAMrXF/51UYtXhZeRkv09nlA0w7Cn/BF5gR2JeEiO/yncmy2TAi6OKwZe3OwvoC8wcLy6zrN8+HF
nR5o4qYlSO/Ie1mumgAI5h3XczL7+OuZdYuXm4GUU54HMhRyK9b1F5YN6/DE+pycPg5g9bOZib+v
CLuTvxJAFwzuViru8vxhky3T6miMLXoVQ7ZVYIAyz88BgMgYO1aS3FJG8H7F+esnPuen7nbLekbf
DSnhTwS9hPAthN9Xntxs+Acz2SiT2mtAMoJFvOqtfWzUVygzxvz2r+wKq0rVfHOw0w6U277ibKjT
I3N8vnLCt+eavr8Zkysu/87o4GszCOaVa0QZBVOnkAbGdthrMYlZLxhPMP1CVTgsF+E/xbV1tAbO
BKsa9B1QvGvzJo/6BUdK596q0nBqiugbvXUbVygD4E1koP/1jZkAnwheZ9Pa9e5gjeJXdi32WHNq
tmIVCjlgp4tbnaDAsWwfcziCe9iFMlwSBJqxKe28FjyMAmUWx0A/Uz3+YlwE6cHyVJsl38sGROw8
JW6OqZ3B133VaPOiKWdQQS+CW41sNGZOGu6FdG4E5Ky1cnGIbMBtMNTCU7JbGQVonwxV3w2pCF+N
4kRNm1fNGK394pp+2JFurtm8J7XBkzuXZfRueN9KII4ZdYNaum69+f7FHzT+VBZf97JWW9fH4ApJ
GaApPSfN2akmUMlJLkGj4iNVvaRKcYVtCnTpNJJwVaMwYQrCpfI/w7CVMKmoPYv/ftqxIUkfxQ2j
LIGGux/cB9fnfS/WwsCzgSa54eNi5Ha7vwf9Bd3BwMSHbwHfpEQLNpuLo7AG++CK6Y/GTjJIOMAk
5Z5iumC6WJWDz8IuV1GT0Vxu7Yqv0O5H5/yPvMPy0tPs4FeCfzZ3Wj9P+GJporZXz0/QTU1QaFGF
K6dgJd5TW3D2ID7nPSpApHl3D/lvbnTSNk4dhmccwaVMxTQm8+EUO9SpSan7fLlyaQ/7eVZ4+dRT
KGRgU44ss/wrn3dKoSs5lodCpYfjTs0Js4lms6DyHK5HHyIzZqzDuKBetoaGYToArTdCJKj1VpsZ
/RygASIR8GBGB6arOfs2OeQvuZ2eaJjQPdfTSaBT8sussgCWtRMCffqEh1qJFkumikTSOA/IXgVZ
xiTtAg2ss+bJjo3/gRaUg/fU89Sbn24/TBTnVk2WHdm1qrBQx4k5Tab+OpD+eXNCSNLoz4dj5BGl
ebxTs8a+0CazRLuJ3qdqJnCdgr5Vme0CkIYht+UmiOzbI3G7LmH7XdVhzBZa2alP2LcFLxxjT1QJ
4kK5tWlKzKP+3QVTW9C3TJ8bj+GfnaFZfKBsfUA9Xtj9Kyts1xlB/G+94XiwIGpVGwoPPpY1yn/A
LgupHsWHt+6eYHMRHUS1s8zu1Eag69pMrroZ7ECCC1V5t0CiLlucOc6TRDJKExaPwAIX1oexPhIX
5byIF4ufiTKENS3mDu1KpLPRyyrz49V3S7Ue0571PXikPC5Sr/rbcwypgAiPjQcd1jV3qEsSz4eC
9JtwOJ7+D4KzO1YRHb0AZc/JzwznAc/n8UucrcIOE4ic46XLR2RWyd2BLnnHSyrccO9dWPNcMhfe
j4minRcbyWkS51IJkagtwUUB39/kDk6m9a8fKldH5Rp8jlgvkuWtbm8mlYb5pnlVyMErDMVEJFoV
D6j8vDxYmIMMdWrcBnh+kM+v3Es7AKjrK192y4Ip0asizNZZG8dBUewMZp7g0UiPnVnmla1Ep4/G
93Ee7vpyivrFSxDQ3xsfqboRRWhQYcBZbxK0rBF0s6CJu7Jz6u9MlZAIeeUeKqzb2ktSjBm3Nrzs
mhCGS43J8dec+zd0XAsYMyBF6ZuvWAWFPz426LhEIa+ad6pBYHonCAtfzPeABA3/73gEkylE66Jz
3DVe0vzWJu75qEh800TCLk8EY8Q9MI9d2U1hb4Pqyt1z2Aii7FYjT5IGIS/I4cY9bxw7MWqbkB4n
lMHJcNQnxlxPq5gB77xaoWzewyjPOJozH/mLN1aLCVfIgW1Z2OTTgfJPlkJFIhUhxwiPzhBdGdiP
sUuI5joXh6yB863M5hQXCxwpI8CNAqq7VJaw6p860BPCowlk9TS1EHuT9Mk3iDt/ossIRxGCI5+Y
jsP90xPJXScKJfL9dqzAOKjqzp4obZqxk7/QCAMnOA5g/fHX5BZH5Si5VvaQ6j78T+lgW2ULaRwQ
kP+39zj5chTBhT6fQiFOW96RmrDGTu9NEuhHFb55fk0MtC9efuj+b55SvLvvCFNbKAhrfrmPmAeY
t/dFRG2zQc8AL2hHQx9Xz5WqYlISU4ahsPZF6rdcYz6wZ7m/F/xdA4AzXCCuss9RrTQu5Je2k6Iv
ZQ4d4WMJYXBNyrE/sbrd7GF4/RZ6szkYU5V53xjnRuJ+jP2vjmebNw4IQY8+eMqS59P0ejb7QlWh
mitOwxiNJeZTLWr/YLVn0O+p2KANXHbyqhRfnzkBnWVWSxZ3C8UJmQlRLQBHKqbhDdN6V91pnU1M
bNznCYAcFRNwwAn0hO1Q8EIqHs9K+2UxfYLhA76lPBpW+pdcILhtCvlxUnh9SYNiTbps3P13ruRy
mWFUG80Wof+SY9HsATiH2W5FNgyxUwgnO1eS9Kv6O52wy52H0CUoe7z5zE+GsV5M6lZbitvZ/daF
NsVPnalkZ+AtUrEEFRtqif8f07bgzBfWocF2MtbVV2RDVFGydo1oSomEXdRwBoaittQ39JwImQvB
0MHp5XUqprjD8D5RdcjMOmpdao33tkkqWiIBcbqgpbgzCkrhkshkrbU+wQLYUwaJ6CN1rnKkjBqk
HBgTgmLkiJFSXXoc1ILA7ZBVLcl1o9NFEAlmDEYCjnnMmUpFmvcW/0h1TbAjDXnm1bnenookIT3t
yPWLPNXImya55l935xp/wQWevt6uyI8ELr4ruBTyceiALERcAlmJJYNNxiqe47tOw0hLqmHgalKI
J6hIImEcfT1o+ieK6ehJjldi+6JD7rMitYadFCHjII4Gmy9X1xReyRccjCzOZBhzHVyF4AF+JuD8
sXe+/BNpnZPMYwsviGCBEt8//dccPLVei2Viax6ByKuu2jSQypdmtmfVwDb5JyxfYlvnasOJWeeB
BVLegXgH3obkz/Jtg5woRWBNtBkCWqiMcwZ/bW5hI6Zlm5psXW6k0p/yACVV2uxLUZQxwTaG4ZOL
+FzANVIpHvhRxMF8NQPk7ILw/Y8zraF09rq33Y63OpCTTEJYzktbhmCwhHma8QdsjodpQXbkbNfX
R5MiV8CwC3Bb4DO9nbrDnOGEVZzSDdjjqrAp4qVpWkqzq+meYRf5/1DdVH8Fql3sljpdRDqI5Bnn
loX3L2zZaXA3L0ChJjwOgJdaSYKeQjwmZq8UoU1oTFbkC9Dvp2LNQ59ZqWp5LP8C+jI9ANtc/i7S
ln3U1S5IDAHJzULmASTD8ka30Pq/UKLLeKcKUN7BdxvG+iVm9lelegK/vI0Kxv0wF+QLn5wH4GQr
g36r0KoWxAtbZ7fo1p8INtE1dFn4iyWXIsnadPqTJzaEO42He5zt387uj+v1+3PyTZw0MHwoXTxi
yUMxgRGvfbHeM6SxhmPPHtFoGy6PmsePuzl2FnrwtLMP22fn29oikBfPTOLx0028k6wY4KsybMEn
Ob3sQP5NohPeUqBa78GUc6UB+M7fzxm5BcgZat+Y5ZNhXbS1wiJUZLpUSlXCkj7VLmzAJZB0QOic
3JDuWjy4Ndx2KW/sjoUYU/PK+Qfpw3gh5B9186OPNO6BaKbAosO9dX2ken8673Zs0YmC7Ki6EHzg
XOxrBgbJZ/SSxhqfvAorxerncUAj27nEUF18yaiP/8qdCFWXVfEdGq02dr8tUtKBpiUaYL0onKg2
7YE00wKPON9nBgrLF32gThKTIzS8TeL+ul/l9MN+3X+ej93tKtOyfPbm0igahhW58oaP0IruPc3t
aS966Zx6b+LJ9RWbNzoM0KdJ/LW99MvD2Jv3bU06F1CiAmTNK9K8Z34mn0KyCw9upDoTov4+eOtw
+aG5XTb0gyK1hIBskzko3PE6efosP/9KiAGI97bD2b0Uqbp0e6jYgoGlMZz+EWlvBe4m7wVLhKMt
Ud5BXRpYQ3xdG4rfiJ5PallQ4HzV2SadNwOF2y6GCS0j3PWQyhnMng9Z6nmIXP+obnIq1MaexB/X
cBwr4qztUVAaLB25RDO83CZELupeavzXV0qOf8A7IF+XcdKWNYXnNBgERujeQTPxAosO/bIJiC8b
XqC7KVSxeYWcU21B0VGsJtZ8CaXj5NnTOVV/SZ5KmQlgfo3GfTr940wI0+2PXCnp0vh+YQXRiFNY
Mc/oJE/rSNaE0BSLdY0JkiKuXfVMEjD243y6VTmY2eO1LeNn3dyE9ifTP71DVzSqKQwPujfXXKmq
ts05m7u/pE3nmlKOBAY0WW7nrbF+cLRE9JUqZ8j36xsOevmdJMLkSfoJNCGYUVMqg8WOoqmUyrvB
7iNsiPFZ1rUl83ruD1nW8aAoquvgVRc9q7WMVxj/XtUZlbh0IXn2YtXy7zrWFdvrE6x720MjhPGa
D75S3fE0WQE4Ypv0sAuycJ5ybG0gm8902h0AY3HnC78sdiaEQ73waYN6S6Vqb5NAR64hMH71J68y
Z/TYhy/e88L/P7vZVLmvKm5wHu5Y9ljTtjR8NZGdt6dUMmDHbhgsY3kMmF4oqpMBiXrGoKw9borX
zJ2aB6/kl1Zzr+U7b4oq70HNh5ArbB0GVESc7/XA/uAMYpKOw6Y9LXn1aW4zlwtsvy3TBkPAxX14
NUEKh+aO2BCLKq3JdL/yYMpY/oCgzefX474wTWHJFslgMy1YsSxgwIKKXAxjNyE1Cn7f3T2O+jp/
YUPYTlxTyYXTtnAd9YuDwfFDB7l9HnWf6RmVMCiHZhuh8m8UyBYBhDlcD+GbHy4uFSIRYK/u63Dg
z/ysZMSZfctbQxKdaP+HEZ6odIiHRgkK9X0vt3RXnr/yWKvak+sYJXsKVVhRLqU1V5ghrXyOfOtf
96gmm6UFBchDrN3wGhQ7/M3rixJ2KUo4uClxphwXMAeOkCd95TYPGT+hkvU/nw9BDSklDsYeOqSx
4+UIYGP4nWgrwTEl6mfuQsveRQJKrZvysoyWGSlxrMsS992eQFBkCjLr+3G43N1copiA3JcWjRTZ
IEROr0OvaKm8RiwYY0OrESFk6CuOtFXr1WKDUYPODAxNToiGdybR7lf8bYzE6bRHnfWt39f1l+yX
8or9xyTv6t5CEXi0xIR1uKTnXxjfNlykJX6y9JfC1W4wdGbO5dkYisRM64mDvev0Lq/dNsPg6l8S
LQVfUv2CAZeqGyxJHe2q3FlSTNAAhFFUY/JQ6F0LE7edtva0teX149kYBktOvl3Ucio4D5+1Suty
CAcM77BAkPPKr/WmEF1Y0CNk6JZLNpAUh45Qi3iMMI/8QLcJIwnV5VmF+NwzifAmvFybWiuLqpi8
wul4ZRFgu4nXZ7TI8+vyI1yT7ZupZ3UsKcFDJ4caJexnNlAvAuMlA3Zmr4vKsnRli+/XRTpbEhtI
wudAzpOUy03BSbMnM65j2tOsFvn+E0BmzKafboi7zjHPQbD8HGTm/O8jvg3v0JkDXnRjtfb8hGAD
szVL1cSjCRVI3yg5X+8PjmrKMQge4VMMHVwAt8aCC00Q10LwVff9EsuSX8wah4i+bP/DHEVM44Bb
yxI0mWCDD7ExZ0FOKDAc7EfKU812KYrqw0o6mrINU0fDUjLEMBwponoern1bLnAvPB64qpUDgLW+
L9iVioVcL9xoFYACAXZaqd4MiwOgdGNydIF+M0eJYxwM5qA42zmOPumR8z2CPCQP7WlAilUeQKyl
SsluocbKM/mNK2rueKFj68Gm9kKrR/jEVAPnaGfMAYnyoGPmmjBRA61TnpJsekfmKe7y2mJ9I6pM
/B2o67fJNKc8FuU4vehkex1BnhIm+/DCW/0M5rukXMkl+7V7mtMuhwuQibv4WwmDz+FHR1XjfDM2
SjZFldDvQUdrf0iPC2CbwhR56oZ+J1sLrTzzRCOuo6ZnHQQ0ToKyRKTzW9Wbe2Gu0CyOH4Smdo9Y
d5baDZLefTKhKbAaWACJ+84CpwV30I/5GBmLrdYgygX6FAkY22kfcqZTPTSyqjiDX16R85liyjab
fUcNsikcBknVhbzpbjq6u6WsK2yQudKhc5CqXDPQVowsjbAw4bu7QQMo/3/cRK025921ooWgw+VT
34ng5Goa4SeGRq/bOXJbQ/q5COdwBY4UhHZSeoqzTR4kvGMGsEi2YAoLy3l4mt8i5j+UOVhpLs75
Z2Zqv/9OBlG8J1VboercB8sZgsHIwmlHtAzzsOBYgvizoJqVsqYeBtcHMAw0Wg9UqBcBS+s0cGqg
KeApRlEs26rvOOXb3/0K8OeJPP1U/7uBQZ1BNoOsIZFcBJcii6Ra94BccfjNRMPYs6iqFlDMLs+x
Y69b8nvNJWxTlHbHovR58ZRZFhfl/23CNrJFEfLJovm67FVGVPbDMAAu8XyL7dztYH3h9/3hmFa5
x3vL9y38pb20dRYN59prJB/hHOnAuK3+7LpZxt90CzbLGpWMJczfE3o96JT3VUPyYPD+BGdsuruQ
pC64XZNBvz5hzg371CMbFKTqZGzgMZp1FhgexqydX5/YTLFkaIiKXcBMUjDqorpwlHepWj3gWrXa
NRjCGoQjw6SLxiIMW75jLPtYIL6/BI+eTfAopXN7TDDtDUd9kiu4UWXzL6gomII1XLD1zTc3rHMj
2ZcDyfz4OASRbqWrDJ1V+o+RdfAb3t35unJng3LbmF0MzfW1Nq76PI3aFyflf1IdLO6OiKDcKAqp
VEahSmJKxQ7BvN7RShdLbcgi1fie4U7TSBVnWk30dqMlK96seWPQBoN+fPRRoAN28GlSXDVs58gR
p4aon/RUMGIDExe6JJHjkNTQcsYyu/lV6hvqfvf9rQKp186w47RpdQ79EE7Zs3Pw7hzbQSY3kq3p
zmiqQk+D8vIUtX/Q7/eZxIHmKW3lEBMvx3FweH+5fN+5EHeuukP9LMI+T8cmxEVSHaK/EhGimTWG
dNiqpHhuLVU7lYRkWmjL1Bf000eRYJiN73T1e4odTMB6lXe+Qtb/SvtO1sgtf0VybEeXWV32v9n3
ga74kMliVcvJbaJsIMCpzmVJ2VLIPbpfHUiojjemBsuh8Vc0q0PctPt44Npx04HPrCVwTJ48j73k
X2k2n3d3P/fFj1hnm6Ubm0QgOLE0O0o6DuUK3w6EzAE7ZoKCAG0pF1fO/d2owXH5a/2j8GedNpQu
hEHbEGqmnQLDcpMirLSfWs9jcZV2cMxWz1LR54eH4Lyo9QEpUGW7B6JQAHriaqBq9ew0rrr7thev
pgku2xI0e/USNaHZOqdJe8P/elkF/04y709sRe/p3m33xr4lD/mi+kGsoJPSY93bTKixOxgNvlXT
W+V8JkQbkA74/rqdIN3mvva6yqVleoEUux/qnUcDoCRid+09u/+CiQJM4p2xkfbIh4YKazeIDzTS
2IDhKQKl+PuyfosNbcn2EYcGJbunkg4EQYh7L+YuZ0aiV3KQyKQCbEKRFkJA4gFSYH3oRCmn/BWt
CXVo0ULcKeGn4w9N2dB0eWzhSOV+dQ1oUz4j2Ch7CJcx/GSicWlVPCPHPQwFjoMCHh6eswGSDB0P
TCfBbhiqV/Npin67oq8L/kBloQhRahZ4J2vbXtcI4LN1VCWazaMQJPeNAnPHa3rEoIqKqeImgyaV
K/IoPKEnpvTggqUXVoR58Xwi9r2Ll7UYMhOv7L6aMV8ZdjvUG62TDlU/ytcVruu9ZxkQ7C4l+iR2
aDU1ymFg+2f/AZNw4ax0H/G1WV+L/Yay7Aarmn5Cp1Zu5EFFJIv7TNyjazi7WfpvOB7cph7Lyb3e
lRcOQ+Lw3hdIpVblNjCpS1SOP9EmAerp39cpH6wLKDGkSSjZusmMqHbHpHAnI8+wLO/SBIOhjY8n
Kcs9lb1SHqDCQzKcK2gE+t1HFNXJLqejohgmwT+LcG0xXvfS2aNumMQC0KIYTBP1EdGypWyOIioW
YwnW074Qa32wZAx7OQL3874W346dogsfv129HlEZp+nP4btLcJnznzUAlZaI1QNtMs1/OmWM9axE
es4U02OFO7Cotw1BmQsghEsYkaUsBjLY9+wgZRcN7TNEkmivrABR2EEE1jmiYVJzFxqO5Pj2WDXX
wPjxydPgTMs1pFfAMhHaKZYJmXnXr3WwgR24iP3Mhje57XffOzqZC43deFegIpio1uxsChfy6jXb
92rHv0zr9fJ1hkWWNV1c+mjjVj8v5s6DMPfrpUiTQ2c2z4z7XphnCpF6Se8PQxqdaxZzJSpgEgdz
Na+iEUcZNMf/d7+gteYcuiPT3CO0T+X4aXsSJRHnQ842DJaw2W8oSwJUWyMFPo8SnqbJZV/7YOBb
5H8cxtDnSQ3Sz5wheQ2t1ZJ5j/f9DHUVGJA96HQt0xxCh06tZZ3Y/szfRKZm3iEYTrtKrJXNv5YW
AFpi6/0cJFYprfymZcbL60kspWCBOC3vX+FqGa9fku3WW65YmdZzHc/fiD6W6DO3xkrrWgXcxAhM
Rw+eO/WXudfUuUFR7bqvbZh7bpl140AE+PgMqJaaeIpG13XqmZpbv03UaZWq6pdutsvtkwDeGhep
Yi/Ee2+0D21E4DStBUmYOqvysqyaJWnx4WZitYMgi4siC7/vrvs5e237wty3UrNKNucXBxF/jiSe
IrDE3WTNfnPZ6hqNC835Ez2LBFFppEJGxEBPY3n6AbVIrJcW6OQFVghfDNdisN7ZZ1p/fKciIwid
o0TThLUSqM0TTa8gs5PxnvjprxTcLVZ/wjsZAHS+E8K+xvZ8voZ7+H8Kb8XRTMVGnr1ijEOe96+U
Ip5Q7CdkwNF9EHts8KYHUDJpgazLQwUJ88VoCC1dLtam/br7RlpOkN9OqczS2xOg1dDdW1IhxnV6
0qiFjV/DmViVYXfesddiJU+frr/I3RMWTOIABwlBLasP7mcyTEbRiJzjUCmIlw1LcXHEjsbVq6kJ
JvX6Cx7l3Ab9fSWJx6YTxycDCg/IdDBR3nkQcTFqVxlyxZGwY8ponPRzN757Ux71b8Dvu/1y60Hh
U1gKwEffjisUwum9OcDZiGuZjGVTeUd5qZYrPRTE9N3owVKTw7UGpVxyfKkvL5DwD6JzgGGE1BK+
MBGcPFdrxj29b8o1mYExSDdOYO9aWWQ2IsZ7j0ipUv+5amhMSzgp3T1RDPzv6MiyKoBR7FICxYth
gJAB4RuzTmLqoBL3VHZWbtGEL0YZ2vEN465S9GqOhb5IWKg8nevlUwXvPgw8beUOn5Fi3yLdukjk
JnSmSEbdi/vBfobn03FpuN40XfqhpA1lP69cO3kwpCG4H9YTAbUxtCFBtpbp14sZP7hnnYUSWTjA
87oIbKhUQZUJjFrToO/Es7/djWn0V4/1Mh3m1cms5x9Pp3K8me+mbkmPR/o6VGeaXqYVtatIt2ta
4nLDitb1vV8RdRlnIzhozvQCLhOrPNwx/ophp+Q2GA337pZyKNNFqvXwvvg/4kBBvuM3OpQNc09u
HZlQvjULOrihRXmngkRS2+AmPdGnp4k7e4rawTT6fLAogJQZALg4+ElIjUnIEhgSZydyJMLiUMxg
1symNO45UbAu1LDMuBMpSannU7CuGVSirrpJ7uXsBFiOICus9BPP/2ZmvD1zsQHOVnMI5HP7SHrA
ox0FTUfpXlUwIKuSIPZDbtzQ21a+QW5YlClYub0Fyk257nlv0OMOPeo3KF/hW92qvBfJs8A8Ma2V
aHwOcLz6m78sMmCgTDghrn/npkhE326dh7Gy6dFRlLS2N9ANxJ7pMXkkV9BS12JOSoYuydKubInH
ZmB1XIFQsI1evQo3wbgK2c76RBHiGT7RAm0a0CvvLlGUOwRYQ/Qi79o0hlGpqp6lwEsjEB132IFo
fsPoF6jcbLFtkmARG8wBbq+YfmUU4ZiE6zCCTptytGYK+KileV5NvoxoHtv3oAIEseO/Am4CzU6o
VCrRNJXoIbyblPv7zUo8TJvUWz8NOpdWTXREyIco01ISLWtFN1lcGUmgSDkI4N5zKgGjwYkktrkJ
01CqDg4dcTUZ9pmcq+LtznZGCv2RLh1gss0gFLQarVLvY0gqe45VIDAVcCVVnKmL2icPgiMc3fc0
j3h3xmbuW4yhpq+F3k8sh/HMSXFs27DX6VaI+nVyFZHpRnIlyLpw3A1RRmkSi8LtIVr2fYVJEm50
qooiFMTDSIYODtdAzDTGrV2J0u6GPvJRt71Bra5TaqryPNI+5uf8whZymJvszUKvNld32QePeoSx
iAHdeDOmVwqm0LLsp6kXu5oJp17t5y9nwHxmldTWHSSe/W1GNjaUGfaq6ncYk0LtnqqWewTz4SlE
CzAhjwlQj9We68DkjJqF5wN7Hl3Xch4gWK+92dkPi/vpHooQNieVYNL2Y/v2Pg3XFp2oKF113PBh
hdAtDRHIPTSPuVfp2nHozcNBcJM+Ae+MbrePYTazV7SyRFMcgF7nm+Q0lnmVN8SUi3vx3b+EqfWp
LIlVpLRi/mhHDl7DSGbdOoSaHqmEpf2R3qBVMdFtod+2RpMM90wgSM/CCSvHJLGmVWAlsC3JeODl
7cMYE7pPagkD5eSTcZGZeeFgw28cwIwn6n+V+9n1tQzu815nWbsYnXtGFSeEphh+0lPiHJ8nupLN
WgBLC+PFBMrWy7Fyi7ddGg3vs5v51RfgipdhAh0Uqq8nDDtKdHIBAPDlRQ4MwJAsDBIgSS1Pyh15
8vOt0g3vikWfXBsORfgsmrTFpKrgeb49wvhdWQiyUAbyV/0rE6S9Hex+heN/zae0NxU1bTT7fYZp
V9eMhk2ivPT2xvp5AaZRoxL9BtqaoVwPoiyU7/jnH+Cl2ualrr6gpN1CLghTitKJXpOrIAM7arRb
WrVBTz4iSHiMXX7UTq/vDE17n7TuWIAIfIpcIlpPbUaFEVd0mtrzhxCrgmNSaMN+BysK4xGuWTW1
1PunXTBEqY127yR74yqrZZZOH4jK9L6BtayH2FWMw+qIhM3HRv6N7XiBX4zqRBMONKLAaPzLTTni
uNhWwkRyfE1+kkwnHE8I6q24C0xmeGpav/7z6akP2SZHZ7SDhdE1lqgn6RvUaHWH8p+5MKYx5c/1
TyiFW5x1ePoP0HnImFV6ooRc86pb9/etzWVre4dM16ro95sfYmZgf1glvKJO4XAYM+k8/7f88lKY
oHv0hbEwgsTLz/neuhT/4NGf9R1XrDcC+EYvuax90aZTKILFT4U+hD+HBeYRy/9lTGWT9wm7rL9M
Fgg8c2LCVidY0lq3CzYUHEyz05K3lSlUH7Rr14xrm7nfF87dBaU1usN2FNDgmz64Pb1VqPsKFVNB
KtPOpD/3bFtI871SXbpOWCkgswdYbtZKCSMRE698NNbIpGZAVjmEa3gOeRyy3KenLYqWZk8ah+m/
nRTczZosdM9yzQcq5Vm6droDHmrN/xez4/6gzT6Xj4xH+XLXe6VyHc3+ajjT7NCiFvuN1pTtrfY7
iaorTaw7jetO4qZ5SJQGwhb4fWyLc1XtKXD8TgW8gdZqAPBuloaVVp5qoPy71kJGk4jhzuHU2sfu
aNtwSD0RZ531dv5Lk6ndo+gPrp3JItkDnBpMlpU09Sxj1Ghkb6UKLbbPP/UisEnRXF4/41IiARru
UGzrAMoIhISgXt1GiI0gMHTI77lahUBPqkX0UmJhg25JJwHrvAuRdfc5Yk5avCRIKwjETqldN1a/
G+hZ1/It1slPwFxQZmm+DhAfrKkkudhClG2ofj80eZr0pytrnlXpW7gGD67XOrdwZWvxgxINVneF
owr+U0+iD7sfI3J+B+44LdrXwv0qjZGXFnxH5hZXQ24dv1Nx6hvu33djxSpvNfUNJBTS2zwHG7sL
KeXSQVDp4pIWj12JQ3leMQ1UKxdEoKH/3IIXK8+iZ7NKmLjUd0y+ZJ4z5eMEbtu59m3M1zOUIME6
UgpWyEo6AkZHdaLajyWLpbl0RRsa1Iwh/2wHof32u/P8pHkZYkfkJGn3CNawT03ZqXqxAYTJY659
3t59BqLeRB51Pz2ugjv89soQi/F1WL5Tq9e1mUHN9+Ly/MZq4ku+/fpDxYkUfZfyJf+F0B7NpWa+
sBKCScocn/+Eu1lJfG1Si1t/xtugnaLON68uc9/9iOXp48fISuAcwDDIBMYjfpVf+zgor0rh1FPP
E4/0UZ/Rudcicoowe9lleAZrb3jE34jzeYu6a/fvEixgFkS+7+KCLFXckkmlzFw8lGAsYsMEeX1u
2SyqshPHzjLZno048XJPRoDhl5C5ttjWTE3e9i3dDLDeCpvy5NPO4cC91wN5qTDa7GF2vIiuPe+l
GNpm2GtMIPXAy+GNpW10E9cBEPDdMVeSRS1gVtEl/AZxBD4zgDzcjeNCGU3TgtQ0VntOzj92dpq/
ero6gMesL7gWMZJyw5cSJhLwsAQ2AfZXluHDTKGfcoDV1WPTRO2LLt/ozMpHbIf2hx4hGtUY9/6/
r4YJbOcG2ugFt1N27zLBvn+eUk+4kPEkpUzqKbuxeNGs1/X0dM1p0IfVMmPuk0bCtDB/glNHWTDS
niSspn8CtnK2PD7+nFM/CWE/4TWbzy1R/9iE+d0VfSOwtUyWGZmEmEFLlgW1gbihNOWStZEnCUMK
EssggLb0JBN62HepZfRM6eMAINpdBjkux3V9JO9PD54nuBi0R/uVcDBrx+r6GxThmiLDI40xsJRa
4wsMsfnsG0/QvkpZBKfT7DwdudZzp1YaSqb7280hRXBtoqHEhJra9z+PWSIqjxh59ytvDh7fKmC1
N0sGwxbyfaAT2ZQFaQ8gGQisy2rqyVSnUzYbxwSngdeObw28GQluYttvw+iW4yunYqEP6UTuLT1W
ihHhRKK4nBReCEJggVKw6/AtltUzP1HE2Ir0cuTGFk+qk6bTBnot6ANJt7C1f8ILJHg9FX3eUm5n
6arp6nszDzhCDp+vx+yX7oQhcWRgxX2s0WOi3/8Co4W/ZK9MiPrRVc7EHIhFRQLBc8Zy5PrZg/5h
ZRlny0DQFT26YM1IagIIoQpIGOHpFTKJsNoitvpPBQWLfKl4yuJkzMTpis+XVsL4jZyrZqZCfy0r
Usy2V2c8ZvqdjzWn5/iFbQ3WALtWPdhIBtFEtLimo0o9upnCt5dBL22r5vvDYTLBZLMdtYUS7bvH
AaXzmmx0AqEbZzRLAxq3s0LHuCUruS92M6jkI4cqQEmnKnC1zpgq8HQoljZfyAwj1bjfw2zuww9P
InT8XHcYI4mZE+i40wLCLWGe8iFcKYSOKWf7kZfDDaZiCBq1t9UT2G2eSyFmw6XpnuPIZIdWm9+Z
kZnOPFBvDNvkrR6PE6uLOsqzSTk6QCODtMrLoTMB7DZzkWI4cWCI3OLWcNI7ZyQD5xV/vk/TG1yL
PwldkFYT24bZYhzcI3WSlPS0n5k6uS8Lv8eoRXrwxPXp/VoN17ijUCIv1f0dhR+df/H//5S4iNP4
H+hdV2m3bAiqAE2C2rSmiArGJnXKpi95giUI21hB76jOvn5FU7FQoA6SGdiZRGMYhv+Ih+Wcw7JM
o821wzzu7m3ZhWCFeNSfaFCk1dMaXpUToJmFJfk6/AGrwHuuDz5ahKBHKRgrusrw/2MhuVX/Y5kH
ss97CWKBRXh6wlSql9ouZExsfxlv4wYneJ2fcngOpblt3i7i2wZCLeHuprLKrhXl+hRClohdXl0g
2M9QtBghvjFFPfesnIxE3rzIDd+zjxSZ1+vzda15VdeGdLS8DiX/A8OJsOvU5swFvfIQ3HPgoiLu
RGUVUxiXWtdKdsi7DJPRzkw242ORsghVCQm/jVCXYta1S1QluZGNXpZ/H4Yp7yZrZxmarAg4kBkA
ZYQnr6NIY2OlmCO4/cNtClMoo+K8gfr9GplZyc2C3ujdaBkO0i03cBj4csLMWmSIvo3fyqqGo5Vx
nFnQCaxZBLKXXyZXSHtbmvi2oSO9NNarSKXftG9aZgKkSlD0/blH4xDTaNRTWxMuBl1qmtTZOBAJ
BiDLjQt9W4FGswaLiX/DB3zGMBy2MO41LRRtxKr0jHqKHPM28FdprjBygAWLMEvv3vWqwAYEVNmh
fVmFYSUafJkvxbyTtDfhJ479vn5fju/TuCJTfatsK5J0k5swlTfH1hxKEhWwyyRejDYDwvYvUs7N
mqtQYtE9MA0V3cK1HTO2tbRDmbiE2/jIqQvHv/B+7iTOzvak8XiFLwgGnkN1+tXDi5ncR2lLgJPK
2m58UMomACwaJBeVidAUsaWlxAHfuD1eHIX6WWTszqXM1i76+bYie0pE2pOoZ9Ss1m9ryA/dWZQl
E/WxpWhucDgyncMoQ0cHe6HOazvtlGKWOnME+jjubU/F6UcGS+xWagXU0cG5GKPnyoc4VV6ZCc+R
zDtNzizyksIww5d/0yN7k+SOGHpwlyHaqWsrlrSmeYv5DsGubmWCLV1q+aON9H38XOFVfS0R2nwc
drLVWEjQ2rtnkiemX9cK2XUiOPsjIYeF8D3zU5zUtXwUh7W52bnc3vZKkuwBerx4tJiaE4fVTjlA
t2s6ONBlBmVsfLFHsHCVQ37hjSuk6TlZG/jLVTQuZvOmLkrUeRDHanSQuoPio2XkSCn360tBVrSi
+M3YMRIlLMg2Q8GTB3Eyq981Kp++zaGz9KRZmnZViM0pPW6hOXcaseTmud36DNOcH5xap6aGBHSI
Ce5ykwFNXKopC7+kBrvHZj0D+3KYUibhz4Bln5aiM5ZNJnACruybufzJnXislgO3qVZyY55UZpDf
oD6E3/s+u9Iscfl9PtDhusMp70RtG7THO8syBDSf0lWzv2uT8QrGVpzgHve048vkIrJlI63Op1hU
EPY7G4zNYV4z//AyVLRSssujAFOKpx7+/OmAUHORGt1NB6BKp+EKROhEJqF92IVhszIbgu5na4pi
xvcSawJCDL7TB+N08Nf27twA/c90tIQdXVB90bCaGTlF4EcUuOYNJZmum38Uv5zb8Jzbaj7RWvGs
EgKr0/pxVs4HLHQ5wYb/veiHjU4SNu9xNiSzYHLD7Ajv8LFABAKlhBz9DuQiKIPNhH1TCgAHVTF7
Xi57TQa+2WFYrInAxHcv5NtwxyojIBIn319BavGv9AahO38qd67ZbX+Fy+YG3Y2/zIeri+kK89Cg
E7qzwEdIsxOHfQGBKwYJS6kzszNUZce6gfVrv5DX/6CcjeptZVmA2FqjVMzzEIfxA4xy8NxWjz1v
XY+nmtJ4W05eLHuorXdL6ps1FicdiYsoHxMiIXdjTOQbNYaFqRAKpIVD0+LRK54EA03lar2CGU2E
FSYmOP+do8nPo0MoLfCVh/5JE9T5g37geKPCfSnlEkI0LMw/fB9iShNvSrOfTNF4dGvlfAv1ViJp
oDfqqfaL+lXcv09B8rOrR3FR1u+b1aBrIkyh4WSu8/y3SjAasos6qxQxXtrXigHHuiRXBo6gc4D1
kcB3wsGVhyo8IrwoBk7jdLiaYDUoQ0Lvazk6er/gJjcSv+NG8/SaaBcMxdgNxELJBXoYx7LlbZ/f
Smmn76GQYOBMJ+d4nEVusiJPBhYQRCwFEmAmEIi/JBNfcaof4ski6tVPfa5Gg8FrbOhvfAyMzV+Q
aB+m5O352RlQyEwfzEfbL8B0D9Kq+GceX4nDbkASwhWJTrjAm5uzZxwcXbcTwaYlXsMeg/k0Qkiw
LL1TQC55vlkKmSfD8SWXPxWpr7J1iwgGMrvrC4Il/juSzeoJQNKmicwvPY6f9sCMFEutj+r7lOaA
3MFXe5qOkkBSV97o5W2DSYkdsvAFuexamCOtGL1sdkXV/mJ5w4h8QEUGLglKblA/ENQV1o2JgrPm
vQf2MQ/2J3o0OaYg5ULdwWKUPAX3u33476qVDa3JRAYyD3tojfpZPOJS0KGvvW9MlVPgP5yFLfBg
NOBCTu5Gmr1ObnwXiE7FY9CrXQJelEBJoyp/HRyPeOyzU2pE431y1SWzaNynH79zebqZbAh47ZoL
k4coeZoI/yn5n01m7EWAt4HIWQ489xEYg6dabTCaG6eOLmQ2WMb4n4ndjEV6KnUG4/LjhWhvP7pk
so6ZQFf04W9U2fCltmYJzaYDvoj3/uPpBRYm//+aKy0xrESDTG5v2m/iZp+Yw0ZZwIB/zwUu1Fxo
ddKxASqfcPV29pqYKWX74rXm3MWo//whwSGawcgfyM5dPDmmXzC+W5BDvf9iNFaYxhPnyZVZNHlZ
PetG67B6G1/X7NXS8ERGjgzxg9OfpKSr3ix93OKqT3R8zyOHNHURHoo8scuymIN3ElQK7jdsacw2
6uV18jPWRRf8v6QcyDg+YDf6hx/sXMNt3s2S4e5NXnd+W4q9vRqEB8pCHW2/DuWHQfQ04uFCkReM
nznDoVYNhghQSJxQQvkmTQNleCage6FROdPFxRXIc458IsBmAfJScRh5m/g9EgYMfdtDCrxMt0bt
VqHBYQlpsyaVypw1oSNV/yPdH6oSxfzphz+/WCfl7PXzUFLcaj1VArvx4VELD3rE9PdFoFkaFR+/
RdU5VFmZXz8d0HteaixORFAPlDWY8xszsmlBj71Evtqq8WnUvagv92Nnr7X28KEmWGA1mOXmvIyI
SSNfkL9C/xWyngT5KIlLEdfL1MevR2rRvQPPrQv58ZvKhXResmIPES2E71M6TkO0ZhQL0kswM684
HtQ7ZQq8bf+HiWgjd6YKT7uxcSxoN0IKnA5Ox98QPm5c9UBVnMiIgQLl+sj8UzpyyrZBP2VoaD7g
r2c76XZ9CcqFwzfZr2Ti+l5oQHJTXZhPJz88ZSNrzwCPC8v/wQS89j5zwuzl76km5Z7qhioh+X4G
HzsfoJirxeCJds2XJAxwsIss2hurGM0wdieoomx1mk0ao2kXkXRbOw3syP5n7VqRq6wJTPDonU7w
qFBWnBp3+jHLU5T6LaoNFI+aL4ny1B5gcfXHDUHzLm+drZ+/qYSgD5pVKUMjJCutd+7JcDdGEYXJ
+Hrmt6nSgyV/5G6KqCtVDUridMRl0VeVao2i78YXEbgjd9c7yINT3F1VxQdyK8ANF4tog9GY0HXw
AlCCCeD+fkMYbyZWbglT2omUJx3zMod7KHtn3eJ8LWIgz9JvOvqGCMwir0eIT8r66FrYZqqoF6zu
MCxpjVpzJSSMX6e5Eb27ItFUu0bIPfUp84j8rRaE9DaeuMb2DUPGcsEBWN29zsjB9cndYsl20djW
WTeKFpB/uLbvNGM2mOl0AlnoQoYmoV7cpoEw/29uh8zexGd20YpN8/lk3zIOltswUlxHcYxJRI0o
b17YXLoTabwZJCsN6rS4u4UaVxGo7FT/yPaZPMqA2UBn3ZLa6UwfHtoiUdJeQlrD6/qAUJbnQ2O0
E1LsY1KSnai6h5lyBOeCezQSjrUP4AxG6Eai+Mx/AIjtuwX0JVR2gY9hAq2sPrOKnZ6dnA70DpEb
80VeJisUGpahqh4If5Nvpq4t0r+NifOpFw5teKrx0CWd1orDjLXy39OCWOBe6CE8qi8dJ0I0/qKx
sQ/KLBpoN0HeJhaHi4R92sl7HVGxJYmI0xqs/hv7SqoAh8L67xJLhFHdqFT0N8zqVrxEe0h7uiRY
iLuyFvON91BkxAkAnsgbEqPYkDhdeiOdRIf+RQDYGBWvKR9+5Vos7YVsnMSoPNj4jCQlIm1mXihs
L/FjLXEN7+5FE7b9xthdhNeD38IncVhnrcbvRTHY8j+KRiZb/SOudKmgwsFMeSQr9ESHCbrBPVat
eyAnifpi1FAt05rG8pKh8KX5r4hBStWht5/PeqqqfeDcpWcJ3JXD9viozVYx7D5zZXLy6INJ1E1v
stokZzrdgEnGZ68wyggqDTKWpRsutB8OhHsSIQeiH3CO+697oDOO6i+nbu+GoNOeLj3nfIaQOFFI
m02mC0u7HCQI2WJ5cSUAiZh9lUxlMVTCQG6ifjET8lnj5wMTwvyeT84OM8/qmEPjAVqGjCp0LT0d
4AMk6T0Nxd0QiHM8v1zhUACtmGcdhBHKU8VB8NWcQJBnZo19yGSEb4za2I7xVSltWznQsZCOJ37Q
v1CI7KDq82bBQMHRNbPnPWjrpJQhYZwR23YvqkjM6NVvtIVc8SGpkI4Lf+Qzk0vcE6OOPgjxS/Fc
NEHCErRm/ElZ5PqWzAif9dARCN/vLVOf2jtynzgzw2nC154c2cN73MRtKlXBWwKrjuLtuuGVsNH3
g3+nJXXyCkk5+TNqUShAsu37kcCSJYI/qd56rw2upLMoT7Hjeg7oX/1ath8rZe/Xs3UxKocYdxeQ
Jpt9ShYpeM2kWqq8Q6OV5S6oUarKLin5RQDb7eX74eGi/5WabxMufxS326hi7EaTaVMNeI0/ffG6
eJTxOLWOP4g3pCXs1BZyBuE+193H02jcwrdEV6t6i1MUawoKuDHU2g19+DYRJUycE5M8rlemcunR
jNK9qkD6k/rd+q+aBzXvdd9A/apdmvz6rMagayh4mB38ldtDfCOgQUHn8m4CYzkm5M+bf+tEcyLN
0godAYBk9BAFX1vb+pteCQFPFr9Jud+xXl3+aIV03YLg66kgKH/4ZPgdJSX47ollyQdzZJcxveGh
ABss8pfvRvxBzZgxub7SLUFZVUxYQnM2uPpCWEheYBu+9Sd67lvsNBare7oqLQbE188KAX6i0O2G
UjHEJPz6RsFmf1Dq9aXthzkHuOfVGBURMAagJmO7kSMlWePLiIIBH+wsi7HHy7zpYXNxOCZeBf04
i5XDG9zetP4c/WT3VHDyjCznUSqS/QxYc6ZqnMRnQ+o3Os0+UyrDqoi6l9y4QGDuC9vgTan6pMQc
Dt5akoNkMx9lAdyVsZTgUiDjmcOJ6iL8SCJ4uBuJHbgehvr/KXctowp09mj5rQHjKdNjHJpgJYTH
Ke16DkEI8+halvC8B9t3ytwH/ZpFOEZ5bcJ1SRQC60vBBtjPcSsrDvNp4am643A1t8kRx3Bi8KIW
yOmjCkKJd5eJiari9qUOVoYq+1vTlKGg0kX3tNGEG1nyp5ef6Jp4VziTJV+n1znNXlKY1L9yi2Xo
ET/1T47B4Z62cu/R+wk9mk1sD8mitp2YTY8dirrcXAEgHekheTgCwEreHtwn2CaRPGVurGChcL7M
Kxgi1+/IwNPHJZjCotR5TCZ41GaiBiHM3RENCsdAZWjVHxQL7BVAya6RuRYkJrto6CdEcGi1UkUF
1iKPqkO7iSR8A7YpoK3WiBIMCg/tYoCDBHAYryQv9VySoeKgDg0CClMNisx+2HLov7qZkQV7SnRX
zZtkf8R3ja4mB2Vr3MHptCpN9gHqA9h7ioxLmyRQeK3G++kFFEA+hUDiwyESvkLwDgikedEmefoj
qEggdJWizbXzPcf5boDBPRP09qZp1SiQZgX8PSXktxR/2vacpnx214h1TZv5TmRsgt9bptoy1vCX
z4Y+8/GY1so8xNP8idxgt5X6PlwkGsWFwkJbSr5WdY6r+9OlEfbljRCk0Yem8nSSwlYtHhR750yM
pBxyIgKCc1E1DuJPLxy8QB6EwzCvmtzaTI7ZxP3eJ1nhkIp8gHv2a9DQWOYbS9Yh/yRBhepbdd2L
XWnJVf4yl0WErh21zQdJUzgOqHqYgin6VTD+juOcySc6XA6btSDCCaYmBTRorEcEUFheBeBxNX8C
v6x8+ZUYhzmuGoLSI3De0v/D3QVRCV8U7/To2l1wFUrvW3VoFaBT2m09L0IGU818ccX7vYt6lo32
0M11FXfZ6OcfZWyPZOu/pFfQ3mydhmH+kmEK+Mp5vMqsK7tfs7my4kBJ0wAnPFVMBUpXFCGXQxBC
sjoG5SsZFHtfzn/4cFnp/ce9PlI8JiRI0UIyYKGK5NsmVsCxuehbi2YeZp3ZTsSlY+kbCNkT9+8s
Qh0pfn4uCZ1Z2tB6PI8r504XiVvIftRInjCHcsp+uDl3Y13QZeTVIkAguLMKFq8O1XcOXkInz/Dv
RJapbTv2VDgGsr88GnYcgkkrGhjj4afEJSIB9kN4xu/u1kprxSPq7NKtNgGDT6ZNt6PVyVUkxjD3
+9HPdhI9/ar3dP4n78qLxGHxNW98zCdGeOYU/zgEotvPiWED+FAJ7SDBoXiXJHiV5TSRVPZ16HnI
v1Q94yLGYVdMVNSPXRQeFvR94VZKq2TBUEmqSswLsltaKDmd/56Pt0JebrJGPmAjBLYuzYbiTdNo
OpvtQ8RllcblaEF2as4N+suUG+AZV9i0SlSMqEFpNFMe8U4aUUCJl5QHtnRVHHeh+ENhpr7G4G4I
clqN76PmUEVNzgyyQKdFTVJoTuDOGLDSNoR6f/xx7igPtRJBNTK2qDFQgIzhMgF19DZwjVq+/xTE
nTVheQaWhB4SNh/W9q1mAGRDmsqFtgg99Ks9Yq1l4rATerGnBzx7lA7XQcyfttqt7LOgzNV0i/vJ
/cY1yJ+/FyEfMFZHbkzWJRqCP2oql47NwPnG0QR9ScyR8X5eyg87fVFoODtQAu4DV2fJH+5CPCjT
mC1SH1TQGD3PSppzUVfoD54Rhic97SUnHCKrht01fWdyY/A1s/yXjROv0uIKPY+oHoqauxpjk50s
kiKFMg9h61Y7n5HrW52UV9vl7/0CuwSN1AbY9mKWfH1Vb1zxRj1z0cqu5YoZKkaZFwkTL5ipzwoS
bLc6eZKQkvK6sIVBUrMDuDp+Ogc8b4u0UmJg1/CU121aUrEAZn8kf9LP88l7xXt8O00zuK31uD8L
iJsCjLAHVh4FPduXGwd8XbghtRJGm2S3ShNUNXV2UbEW5nhcFlAqoDqtKJAYN8EqbDx+X3J/9cne
1inTeISdzMhhXdAP37rdpizwGb6cpFdiBoAGA2BhFNH4oRyAyfGrUizsz2lT4wPiqCD5JpUpV2Wy
qHdBU4FwWpXtckyGtJON7nGJfGbRFELJyqQyHg6+SDN8JxoC/UfCr/4dOzPy4AaBLXxuAVgUVTMK
miBclGvF4P5HzzHUkvkZMizaWk8MAIVwpq8ZlhD24RajEn9jalDv3yBPn2yM9Dc8nknQP0e6en42
tnHbdVgVtuCuhJGixt6a+FJvqNB9dHIkiCtRLzk9JrZU9mRlVVPmfLTIa/6A/sCY4WsiNtciyZ4K
JZrPyRrOv0DfWASQBEGIjiHzyuiQfopgWjg7zO8qyGicEuuGZz4SmsZjyX+yEs0gyP7zetJ6yoT/
hu1LGviP1fftnWVNFhvF0s94Jms5rkmkZfTzVOlksPQnLr98ZT1F7HIR94cWjldy1KeIbjyP/Gw+
UEIbdg8uQa7m2BOVAHebD2dd5sgsC8XmaCbAdT47/71vq855b8+7WqwY9EJZXJdJPekU6v/voK0f
NOsLAlpVpKBY+G94vn8mXrTAvsXXB/kQtf6Xl3TuFbAMIt+wTlylvYUneBlnwEiLCGHtTmJHm19j
UMOYzaojpGQgfS6sGsHdBP/3F669+s6/1yduP+FQDgyKn2rrxT0agh+CEIvHz87TOHBz5BlWm55Z
h73E3vU3oSIHQTN5LFINj7uBmsTgWbdgRRSoTqXJeLg/piB2rdpz9CRZEelsPddKsOyppKoaCCml
OO01R7zmNFQRdJsNkeuiKG4Y8oCr7D45h0E5+RvgwbWbmDYQ1Qolz8CgYb+sUMzhDDutVEOSFMMg
AGQc6OzArUN2k1ZgFoqIHhQki8sba7VLMDSCd4DDNmmnC3LTxcNs1EsfW7WBM+LdHjDXLULWVU/u
bm8UXK+OtJX6PanPnmrqz7OSYcmnaSjxidF5yN5nfsnVeEEARfUbbEWcBBrS6Ab2Gbz1Cb1sG9iZ
MQiKIpg20JtEcrNeegt8NpULIheLNlpJmdHs/jInwI7hRu7kQolxBB8L5+8ZNcjj5ACVF/fJSztt
Oh/FD2as0ErvK190qeyTvk7Lm8aVT91PsSrziXfmFeo8v6jOPxRL76/3Ypnj5HW2mmVOWxPGnn8x
72NUJunjFyXkqg4D1HNygLDechbp0sap3O+OLBzThEYUeCIZCtoUV4Nj1BG7GCQNcXGwbCsOmBN2
uU5Rt6qwWPZlUg0KZ6jJB9+/Ps8+E15mfJBrKUHr7mAk9bnDtR2tMZbzAJISOrNSA/6o4sc86BoA
c2FakDlMaXi2jQ25FvbPwn53NJYYedcrR0mROseEPgaF8nvW5Eju0uhJuJCJLEUvnMM+Xrc7dpRC
RuL53KPW/HzE3hfg19CsDiB6hz9fssiIvEaGsl6Nv8sQMzA370Mh6vdMNGM9hAvMdSpH3p3d0c3j
uq0EA55ta3Zpa7Ca3a7RpJZfqu2UQh18+Wpkr795BlpsjQ6JW71pTjBPBk/q4bjrbZHeQdIrGkHB
OyRmUn4JvsWH5D6gCwxZNXow9+B84njsK4ebCdKV28dEJI5Lb/V51Mg2NTqeyzYOZkDI1yT7i+vI
7QIZnD55gijO8KC2BpsWF9bAbsPBmQ9scVwoPBm6OA7eO2vAJy0K4FJIxlGzFUObTMuR8mBsakka
odJ8ZYMxGMX4pSORtN90ifQJzIKDPIGmRkpBSN6HRVnlwYJNZn/LEEJJ5vz/cXhpX9LHASpKB9LN
sy0MdptemhFxZz2HsY4GZZLl7rmIy+FuunkiNG9XhGJbR1yl1c59kW15zncM3A2jrT/MJ2ADHt4X
0Muf5cWfiWkn6OnFC8M2F6/aeKxq9ghXRaxqvn19uT0Zw9MzJEeMekFNIfLEIChrULBIHrxoVTkM
1lN3UJdQDg5bAqL5mh3QMdJMjNOxtc+0uFMSmPrjgUjv6N7VSMiHiklMcHYonXn5xoardugQDKme
ewQEC/ZVcOx70d0PRB23YxZa6H7LGI5cEn3jyuoX3+x+do/2h8O1ExWR9VfkERgoy/R3spuQ/ala
huKq7WqMDT4P3lPVPVdb9MOFHbEZMcKFPFPdgHKsmpqfvVq3YH9UPn1bciZmVQxwcX83O3qMfeaL
Ig9bxZ19hJRPoVIedyalP9AR7kmbI6g4Si3VVKjT35r0T4CEromxzZygDJSvtZzDKoLXA79LTlpZ
5HAKulirEwojiTpfrSJxBtTBCnuqOC/1FRMh5Rl8+gKsBBMAoZlvtChWtwtudyAfurpjuooVJQii
Ki1WaORXmBfVxvQEv2RrtzcleHSunex7gv52iuQJv39acAUXmAfgrN2rXRwdI20SujwqBIqT97CK
to8v9SCZWfMkHwHDu2WYT9/TrpVJADowESvHG2WDftbLcnFFJfmcmU9AW2kvmnU93DOW/CWUquzk
eAWpoIfcRkrTk1VGzk27Ck9POuVRpb6RsD4BMkKTlie3qhqLEwIkaFn4kg9Fi5LbzeTtVzobewOY
Dn/fiprW2Ea0LiwEYpd3L+HCXmOUDTMoht7UQ2QJkppk1IAnDi/ScpvJkBjltmdNIGhbsVQZLsWn
8GbmDqGJT7NCJecfB9kDYQNTCaG6ikuzepnamKqCfzCtIu0USd0HCO+M7ZN/GJo/cmiRBct9G1GN
abaP9UZJnqp4dn502TlmWEwiTOeLpC70plLOvcb1/GslqsckCw0sfaYtNcH4hZ4JjGAcj5mwNSgD
X8xyRAc4uY3WSqWGTM4ay3u+4jaaFwfvt3IuolP0wEPeeCN2nc99e+VwybIJHVfe0DaSFwkloPm3
b1J0cydkmcTNlraq/MC0YgZC/fUU1TTpIH82GaeZYqsZhn7ck2NaoQpBLqEDjmAFr0dCJOk1bJbr
5TV+nkZd9+80bqdX/fa6K+ab14aBPtl5t1fvbIx4VJ14Cz+A5C//93UDJbnRohzgFpfcINfiVHDg
mjTyxqn6eiHfC04hdB92qUSIZYn6ZlzA9Yh1/qH0hOG2orsJ7EjcCJFSuAE7iYavTtHVqcjkQZyY
UkvRwzK5npd/WeSsoSGNFBQvBcNuzfdKhl1jjLO3f6ftMgjw5jsrTqomHHVaOuMimjlIaeZTT2qa
pPEaNXdHl1+J6qPa4JHV2iyoI7jfyD1PzsAhOX2XGkNF0BYfUi2jv9XqyWFcSmULMMqrfEc75ps7
j4JPqtvCH3hnk8M2BgnTmkKnLzutTgysh4IBO6sjQjoUl8CpLW4OsERqHJHC9a0XuDZTzkIzFjmZ
M433Ss2z2P+g+s+0tt5tR+biMmCS77RR0bBz38bH2GfPEGyaQpn1HALfChTUzC1qhOuE5TEZKQkB
GvN4qte6TWGhOmJ3GlrY06BkjzBu9J7VsjkrAf9iCkfQFBTdK3iolSzL12FrhzziuhgadYksvk1I
QXA7ocXTBHPOrP9WqDXO+0d4dB3esILhbuE7aKdU3N6TNY5LcY+Agg9v9YzYGaXt6uCsJnmeNT6s
N/nx4fcz49eeY14F01UrPayJZQ61IYCnrYb102x9n27Yh0r7lzIz/a3BtlIlcu35gVQT6ABbR/5C
I2ke6SwhasWgHL8UABhnpWANAZXUVoTyqNsJovdzZMicXgDl3jOT/6KJABISUgaZvAYV1Od0Axr3
/4Kwqfaeh/jsHKFxD9HmQhCshkLWkBHMliK/f2NwGrZovlXLJzqIQbP/1gonqD90CtADvrBMRs0c
YGvQk0G1QZ53ukW+UyQgxywDqunyE0/L3NuHsyA8yTXnGyHKEaEc+56EkfkffCdmHUAPAxZzThZc
TEBrTdHNbgRqJKz1ngnyqc7hAouyhIOshnlKGdmF9twWtSCTn0ZH9hK14QYl9K8NZrkzrz2iDDNO
I1nWmBkNWnyRkqiUt0bt/0RQ9DZOl3ET3vLVp3I2xQDgHY1MF+aNhUWhEYvUqTEvlnqtwoRTKSS+
dhsil/EvfeP0N+Ufa7YpZRDZf7sphULXIxkvLglVwA9uV4EuwWANegk0yBWjsUf6VEjB4iC5BZXE
JvBaujSgtX6je/156H3lEXmwhh7CfATXKND16tj++77LtxZWVvcx+NhBGX90Z8G2iuQG6Hxzj5Aq
r+psFCHEpaMMd+pOJ+PVKRFBMTeFT2K+oc5Y2QHkVnIBrffVUJm4ITtq/cTGtbhEAAYs7ltdimUU
Ib/yA3Jl0fgMRwpVSdhlRcDwXx2SwJyltBMa3tBgO3B+w1aLDpP9BinhtnbHEckurjvCIWU8Irq/
GoMKfXwA1hASgK2dAWSUKK3s4kLHt+V/tSC/BlbqUUQ2I83J4sTSyl5WW7Awen4qeraXSbTdzkTh
yRaC6I22Cy9GZCbcUphq7IZrqro5XSeNfCRnHlqD8tRhtdBTpzYIlUV+JIg+77FZ+ti7BFb/QwX/
Zx8CklV3otCfWA3lvzwU2tPl/ji+QpxGI5BgGG+Bt6VOFKLnuCO2cjZktWMpSFU1WyIvwXhrwxhu
1M5Io4Fo/zotgKKSB9gzsFcm1UPDJvTrOGr9K77fAWoFpKxVByZ33bkIH2s++K1qv0HFcDQDpUcX
8AU3qgAMG3zAwSWiLXk+lqE+9vX+viBJqN6lwWyP+l6Xu9hn+kkuUhulWKMWD/eVUXtEv7mrscCt
IpWnhAKKx5e3vM/FOrmYS+LQm4xJPxN46KpP5WiMW4qZTHp77zMEzRzr4dqtU8zSgb4N1kHOse8b
rI9uYRT6US1sWDdpW3IV5PWPSVuHsUmMSfurkwktpSUCWpyRI2dk9w8KxXtYcLZUlmCAWNOR8V91
9oYrtWhdZiJM3uRLmLXUy/BmkfgQ8AA/WCKg0Mr/MOClDsMVrNbIXKkydJhbgXbafNroo9G81u0z
vlPXz8lCXuvu2fCLohcZ4UaqTxIecgxRbcPdzmXoQy7lOZt2Pu09KKaP+LiP54J4fCQKEoMfer59
Q3hEWgGaOLIxUE+JM/6FKJnLga7cKZ5Miihq9VqzJwyFF6nNcdqV1KS+fpqFYZWnGNNHQTPO1TMc
5aXcSv29qpidUbq7SlxJrV1qWRyTj9E1jKvNFOEwbOuvgiW+GY9gc9wA65lJkYdlRAeFiZfN3XsE
XM+9OQ+WJdE+7D9kpx4fHO6aI5czUHj7epW9PPrp8dAPtYds2pAjNsPnC17c5EUjECOjy3P5AX0w
8xFyjaBcCBl/W71C1tKnJPKHkfBySGnRsGAGQ+GZocJMd9gYo6OtP7RFTBl8TTGkLvw+7juC/IvI
hdXYTMpUxa4O6WK1XKA7n0rBZ2GIkIs8XJr82F4JniKddNi4ory4tmGTAk7dX58A0x6ShfekVbZz
NVQn3UU/r9ADFoPtxykRe1pRvbOHJiAucgsSGSW9lWOKgHielKKCIHI0EwlKpyINAYkMrpfPdRNv
56+Ay1d1lcCL1NRg6+/DN949a5kMyNCqkuTJEWh0JCDZvAlc7Gm9K2iwRj7nrWWn6jqOOvqF6Bit
ihvFKUWZsMVLtD1zhzBKWcH1jEA3MxmquxpCZn4hvJqUzxMoyWHJq2szDpFxKZDM949HZHODs+75
Mg+Pddl/WwPkhqP8q14Tlpwn0UdHv+0P4bHk9zIggeRa0XPduSCLjRVyBOp+mm40cpIrJE59+quH
e/orIecd0dsEt1xHHm1TROjwADiE39NYSJfINcV4hSczkgwfPJKGoLVevauV+61qpqWh5YP817js
3Rx1cwQ516qIah6BL9PTK+OEMCyu12AIa3EJndxElNtrZ2+x4TzFZSvzItXSdX/VL5hoFroSVknt
o91Tc8sAeQkleCU1wXLtuOO2Rc9RxxkYJOOm/wJKDJkgJRPBnB67FGSUeYwtCyvxVTLjYVW50UxZ
QKGC56UTBX4gSu6+tV2dnRBM5fTJxPhKlcP3HJQlRgaqHojBne0WSq+ccsrDwqKbPdkqQwgTQNtx
IfH3cVgpcJpwX5abSuoPDRnTWxU8qrtMICtI9SYxvlnTd7aZm/Sr35bmXz1zwG1J/eNe2L4k6gEh
APDD9usiYfCkIDod4XVPinYLVRp5NDX4KJO9JYcSxrAhx0muFaLFNyGYgrU35O27u2D/d6TLirJd
XIV6JOsT/HSP3fqo5q+7Vgq99WsXU21myLZX69VcbWJnoG6zeqpYGfREkleYZnUUmFJMqPnZ0D2n
eY7ksqM61mcVVizXANmlrLlEvMB20kjihEJbhiQ17iZ2vZSbL73v2LR1Kj9E4YrBZtUvTSSlHnxe
bbSTOs29Iq8UFd+qNkfa5qe7pa/jMnYRyxIb18HvX/mLrEdKRe8dd3i27kx1xY2aYvO9QHh/QcM4
Uu3QBarR+aVGtLtYmuv/oPRMCFM0W/2BGG82rc9HotngM+965MKTWpgc/KxXudOrnEIulxY9mnuW
xrRVOZkiPsOX2ie2z1qIDxWBMsC6oGso5HZuK6Vg5Ibbk4XFm0/JbJjetL2S/W5ME47u3YSYZ6xq
vvJOhMFaNeuMHKReQUUbGF4/VvgkqQMlMssmxUVYR8nAKo9bHlEyQZe0OdN7UjG9mZKV2OQ8HWj6
dwf+rSeX5pfZqrFZw3JBBK53gHepIR1iScz3H3XjqFa8vNoFQJhnGpxlEZk/P3GhkocmziwvxtJz
Ys3Kurx4tsmpZlK6xRlEmQn1QoeLarh8uiDyOsTShbQWYb7fwgAbsCMHPhHYQCfEiPElK1Q+TSzX
MpRS8ZPCjqXdXDRKzOCbSUzt66hjAlkxfbkHv3R7ZY9CEc+RQJoDzBT/VB4yKQ5W+BPEU1bHnpx7
JNSAt0+8cxMZMwsh7cb9ifqRXR5ZXD7CAclI9fxE84gbNDZAklBuqbSyrj0Su2rJOjAyZZZGR3Nk
O5Pru8BWkdqDVo8JKbInFn9V6xH64V9zCqmwbUs8rmq0z4LoB44CxLMVqINpqH2pk1D418HHml+8
g/sMlYKS/zpszfVXXtUNmuS5B09rfIAU5MgVGjY9fJ8WQG3K/vAxZxJTWP/LvE8FTLS8IjQfrVMs
8qc+ftHrS7+dcAOJ9z80FJET1crH6LZ5D68brzcgsFs8s3gnWaKreaGaeBZI3AjeiwDXuJx0IAs8
yYk0l8oVS4halJiGiDuiAliiefE784uhSyWhRKS1w0qoVD5AkhUtD3sKNGHQf+inELCzvYejrJ5D
LfPZRy4/ksAHtlYh+oqBLkeXzrgLbyhOKAvO46Tmw3R07mSJ0YW2cwNHYR/LX4+VTGIccoduZmxu
CE+dzrhcID7OsT+qacAE11CvMFnBvp4+S4Lir7Tc+j5ot6yvaA4LA/PxGk1xWlPVBie/OgemqwMm
fR/CA9zLBW3C8ASwcpKOKMlQRqApWbojkLxR1MRhbH3X2C7o0YLvS7vYyNwKbTHIsGxJYHrBoUbQ
ycP9R9KEDmy4vIJgEHR4jON6ByrdG0B9uYzHhbays06CtGhymwb2Azen+gVLveKjGZSSxJerZHek
5RW/v+E55/gRL1uLeGcR9kWaJ2b+T5KiL2m+Sy4/2vfUWEZR9nreN15/FPM9gfIccqzKvAN9WxVd
IgwwBUkRVvlszTV5yX+fl3FiQ33UBTzfWXA/CdmdpTmOXyBS9VM5Dollsp82Uh01OhRBNE6WPCvh
e24cV9YahSsrq/G66yJ5lOgCOlFMGlO5z4HKKIO98WVtxgg1xSFrISFGoDxQWZs4Ka+gpKoRDvFU
G8iuMdmu/R/oHjMpKKkzK/f1P1hwLW8ER151txgRpoLvfcoZfurzTKeuB37JLoJDhZrMXNvxaP5t
C4nvrqBJWZNzjtGJ3hs9TzOqHdkOkL7bO0sx2TCOAypbw9Bb0VM+ORDjU14/mX8YOBG2OWl7oCN2
NHBKdUlwj+PP63+jg6vcTRLrOXIWtoLJyHKs36XwOem2NvN2pJJKyA1y2tViTv0fOavKveLuquCb
xzibwaxno7zKcgFFK66OuHBDr9TDDpABbhMLqZM0euldeGc1MCstcbVZWK5VdD4EQaRM/8mRwbNr
A/XbOvbBR3RSqicy8h9P0XGrbStuFVtgzV5w3Jgme6qDG39O6xXoAEnZEnXgHYmp1oEBjEMkUljv
b7QFcLxqUDWEa0ZVmhyaO6g9L1r9gaOdF4pCMdX3+qxx7sUI2v/TI4Ccrx4MOhrvlVINITqMb9fn
dXBimmMzr+zjTv5OoluhkeFfqCuf1qvyEUFtGmMDIC0irzqj8p7/hUwaHODgWcTwiRoAejkb3Vao
dxjyL8jMbL1ATIyhpgSWMlWa1gx2snzTSZJ/gnrB+fkyI0s658YOSYyLvJSRhcb3rbKHEkEr4YnP
bIppzEzU/e1RPGeVgV4cUWuKpnYGIhyUMx/diggXLR6yUpLODV5J1AC/IsyG/IKqZdSrdnhPiDju
oMOEcNA2Rq6+mrGXaSgWoBvclRvccqhiPxCIIMPT1LoMytMOXeVNC6+YdJdXMOPKnp5Ams2tgarH
25R6vduxnsPsOqhd3QFZ4PkhygedNNXtJNN68n8PYHTnSQKp9Abu4QEyFNhMf5Hz5kkzq0kaJENr
c7TGDLlBB6sB0dUwIjouZ1kno4HGQB8ycfY00EihuBKi9RVJy2Oy5a2cSMsvgevdD6RbaGTmtvNZ
+w3FHbMN6/Z38HvwFn8GvsLYh107HEJqGD5xA7RrWI3H0IzwY0NAWj7DVDASGlUY0HyqmgChHcYb
+cbbweIMq3uVDFJhBihhHGzh45pQjHjPDGOemwTgzWSXh13lw4WeNAqp+XJ6SGueI3Aw16+v4dTe
+HFx1VrNh3js80azB6C2fKYQEQBmgOTMqySFcwJvQyMOlJMvvYzd28NLQrnszj5NOBl+i4T530YP
P1sxUWd0NU0JbcTs+9EipkkaPJC+RRhPUs2cK3v6Toy+dRfq9sKRQikjVXCRTqf64/R19S2shBeu
mvdVHRACDqrtjTg2eYdWuZWJ4CHNXtWpZuj4JeWA65CAXU8A9ogRtqzOg40HrOenjdP/vc+ZIyQI
Csp6yvlXbfes4CVLKg4Aq+CkLvk3t8D15ACuqBOn6m/6l1vXIayTkjknkBzhegLe5H9d2B9Q1xZl
VXMJVvnhMkGE0tJm4yhDftOQf5pPGPZMRMtmzQfhFBQwkWNaBRax9Cmt8nMqD3pgCcEDkSp3KhbQ
6HuBaGCfNQKyHuy+lowX6z+Ib/dXXVjuR71xOJk3QBlJ5tJOpF0V0SCheXx2H9w43jqkihQthzEa
4WOXd+PYHtThsEf4PjDrssWHUOA5xwBzMy8hNJn2cFqBW+SPQnC+7E6ZDBQvrfC6S87WM6xCbrZ3
2rWGNJcpvH2kuBxIXsxav9IqwAhc/JyHRRkebtHMEVT67topEUjRsMErYDQzXHxJu6A6mPoLS8UK
s7gRDsboj8vQ9yD30qlKbhWwpt1qigveYj7MuEC0lKZiuDIjPEIrWOWTyFKa88xs27MgwJYG3Ves
fTFJrPdzaKrFe4n/bvbMQD9CbLwg61z2/tFqtOwHgxt9WoGZN3/EcPGcbHefvl1ZvCBqbr9Y61AC
BPvhEXiRBCuOuvhadhT1LTkwhBnceg1sVKlih8P68oBJ8vipFwS+R+pZob+vDhzZ+YQb/Huby9cW
XbiqHtOPQtZOlS/yLrPqe2uo8WvotdhnRb1b302TD52HbJomDGBosJna8j1kWm1NMcCz6emMucGo
jju8jZs2dTMFJhJfow8lIzdhCLNJpcEYZ6liX7ZKbm4VMJGhoRCJ2X5qY5UXJ7lEFg64Go37HF6N
tMPid3dpYe8KyV1c+vg5ykcEnyd8FbDrpkaH/0MwelyPftMMQZZwu6L5VYMOyK1wyMF/tMgRcjew
W0njqZDScBBdcgBSrqQ/Ehnjfglr3h7Tqt/IVymconfT/VLJx/iHPXN4PMGEKLNW32t43W7c1Hii
cvqxGWyfGbUCvSYXvQD3crTka1Q8hwYyEdXlILfcOGV4FDrnFrzUr1RuNAg/rDtRtGJ9pJG0EA4Y
gRC1mVUxOeg1KwOIVoWuFnYPDJ4BZhHVcnUbZewxeoO5CXJgLipBB6j1lD3VMUr2eh5HI9sJrLyC
JS2RrXBrojsJXcjwc/E8MFzOT5aZkujJunVeqPqvF7xi1tpI8P+0gGfsyha63p9b3xiwirb03MZI
o6VCDk1P4ncOufTYS1AhvNz1Oe8jUtS18VVkl/JkyNdqFfoZ0jzfSXN2YEv5u9V84KdgXqCk2SqO
Xyr/VOlmzc/S4fFKDaL9wmYIh7mkmv20jxpEkfo/u5mKQTytJ3sQAkopA+e3ZNZvOm3fpz5GLVaA
4ATId2lQnmfj/YQOL1Hh/gqpCIXnlSZwtKcg6uC8XAxo/sAdlxC0zlcAXlH+bJ4BI7AJXrPdXpDM
B7N40Y0ALzpV7bMyG2u38psgKeIqgzBq6UlthEaf0H5MTaPU5zYA2JFMUFfwYpiGVtqdEHlLeQdU
mVw9gQJDCVaI4BhMvMRzfxW+Kqc4gXuP4Czfb9KOEMqBoQkJPJszdMlSuLTgGqXcsPNoYcoBYcMl
f59sRGupWSfl3C5fn/t7j4Nw86imAJxUHQ9aSlypW1bVnOMiTZFdWh/ud8JqT5K7Vj3bntrHLH8V
6TpO60vt6n2+hrD/xiTuQMqQIQZGP2+QRDF3WgCdMp/AZisbqyMZhNoeU0mMt8iw/sHKxxLFKwPl
sJBLH7iBuHumpn/tUP7np4d0s0bGWSMyT+JDylEM8HPChMVNlrdISLjlVRCnGSEjwCyTGf4Q6E+9
u+J1Z9eWluOUYiDQ95JKSLOYMeiW08pUCltLM03vCi1JfvU4aBiAFPlhCZgauQssfcxuDEKVGtce
85aTJpBrsbzDN2vkIt1wkZxLGzX33OZ56S6YMO6ObghCkLl87ta6KFs3+oZ+JtEmY7G/TFBrEEWB
6Gv0qdzRmOft7LVrUhVbvlia673Me2x+99XmyD1qXz4AQFhw7uoWpqKRMvHUHTTUdOI6Qmut3sT6
Gd+ya/sodyq8Ynd5vq4dnaRXOPIgmgy9sxWKMFMEoumtg1xBTvfe9LqsUXb58aO+ae/ijm8k/0J0
C1E78ua6/mO+a1fBT4dtYQxaNNvJ7mbXyI2RVVAuGRu7tbk4oCBglubA3UFpvfMqVtx6/DPYxw4v
N9hAKMhkDKQouc/XDfSYPN/I5gZ7ZiUk1UkMVK4qpwgMc3qhLJDF/fdziS6ql3OmGIN5U7r3Wp+s
6THTZQdurd3f9han1OuQFaHTfbz9AyBuz9hE2g24DBAw2CB872unaQATIKFTIqQYDMvlHeAJDPk6
LVt9ifSmDTx29P6RCfJ2MfmA9A+ZzLzuR1Eontz+qC3+izqliQOJ60qOhhJbtzI11GSIYqPrAFu8
mCt89gdvx18Qxi4n/BjMOe483D4Z/hTL4iYvvLjcUUas0+TxVqYnA/26wYWfcSLRdxbYqhzP/u0v
CV5kgt03md8Fx91uw2NKGhGOc1gnuElaz+YJceRDOhc98EmowNUxH/EdlNgAep78f9Tw5O0TIzaf
Cqb1fqoM3EWNGaRdJsUsCa45ct0w5E2QIzBxywKkt8PuvW5ZLaT7tYBEJ8L/1kN/dA24IoA+SLeP
CnLj2WgUrQhWd4Uoe6hrCTiwqNfPMgqngMV0V9mSkyODZqcVqFXdAQyuF3M7BGrWX/cSQYDFsIMD
0AC5qph39V0piHIj6LxXqAtnm3wdxXCyke+5RWor4pzSnij6GKiCE5BE9vtXEhiFvlkf7+RbSAWH
ITty1DZ0EIbyibWTpvjgpXxH6S1NTwXDmC8M7xc3TwGZ/H2M7tANEgeFEnVqZfeUFsZwLQu7ZVNi
qOKPkDFPmUHVmpslF1iV2xSqGUsX+JQsK9boZ8oFWvMbKzAllNjIgmyrSj5IJ7iTT+8eryW8cH5l
C79ZQ229NOrpvpRBkSnGDGbz9R4MKpjO3p44xteaj7TRlr9MiR0O0T1z1PnhNIIS4yeXoBAjsSBm
wqD9wqxN9IH4VJzUyGP1Q4SkvN77pagMK+lSHu4cF1Qr1B2MEXGVfR5iEBcUqWhXk1+3RTYBGq6J
Yru4wgUyn/c8JUS6DvJFi9OinC6X6NtLwOsr595Eg5cWNsPC+zDO1qSdlQSyyOtZInFNcBaCbaW3
BhCW9rYCJTg1jJK4AByG9GXnHtCbG7dsCT6se0a14lPhbF2i4ZSVaUvA4iA1yMGy0T59Dhd3wb73
4CKZXbPn8ZbULzjWObTTjovBHiRIP2BFDvwLsM0ZmMeJECOERR9IMgkSgmOOZu4gIXxBoeo69VE1
hxK3DtosnpLU4QUy/RK/whOVenrpHZz9BThfwYGtH3d+IXUT41u01sTFZDNJbOumZv3AMIys7W+b
Qcep3SHuVLWRULVItfa00cHak5ED7XVFCTHZ1SDS7s6bFTK+teeIJfcbt0dlRy7Av/5pfCqaDHf2
mNy46gDQmCZ+Q4X4jPw24xRm73dPPA/3IoTcVeolIVzLl0maFBsAg9nCluFsDuclwHKQeLgrH4vQ
YsOX4A7KV6Kfbu74eL3t6dTs/2l9Xm9nl3AlEdOY4sFjUJyRTPoUpLm0PJxtGH23aQ37WRAd73rU
gOPaFczwGCN3Kvr/4ggyXxQpPs17bQGIY8/0d07k0CXK6GlNo9nQ/p4B6g399bSbMy82naGbYuKq
qobR6N+S6yWEMTBKs26DlyezOGQt9BzL3Sv1RspR9pJgk4PYWrD9D5J+53eb2vzCxWqkrl/dmiC5
iNrJoJBI+oG1xh4lRR0YGUDohKy1oK0Vc7yDaMkDX8u3MH7Yq+ZGAYz54XsxoEXaecLNiPWAXD2m
LaDJZjwflZNNE9sg7XO5IMOPivnzEVMSdzpfdEEyxl7DWHbfaMUvp8blOlsOQqiXzogQZNlgSbAq
XgivyY2FLPrKX/3JGzAlWQR0HfPI6mKcpIDXWGKU3AdoYHna39WjZPYkotZs2Nl6Ip0A9Z7eor6g
CVRcF7pvGki6uKwbjhTSmaELWCH8laUpZMN2XRpsT4v/jHd9IqWWImcSfzNN5q1l6xXXhUE6C4ZL
Dxf//4XpexOicNYwCmRjaI36t2Xw1X6eNlztdNWyHQlGaUZXK1G9pVeVg2iRHQSIFbCjxIe03oRZ
tS9sg120+BYNl7daV/Rer40FxdBLBjth3yECYEjTIqdADCNbZRUqUjsYTff59tzodDJp1WCBpQaV
AxujQ21Jf/5cij/zetpc4kmfrWoznzHuUPrxJe3IPlvqrBtCM9jta8kjYJyiDNITgYKDVRlAj5j0
glHIoIsLjUlHwNDjB83jhkHDGCFsHsKscR64AG/J1gJ4EbIYglR/+kw1EHHVVFibgsR2QlFLORJc
uu8pVf1h2kv0AVMYw93uSp/Hb1v86lLfl3B5Zas47eCqw2Yzjlif9nPVxCuSYaDxskFfBqgES2YJ
5MF0jVIL09gahNskQ7/TLXHU6cj2JGcn22nHazNDY/EMkQxrqYl8NCodohuhvf1K59rCrOFeslAT
CmrfPg5izHwfIraaLT+ibG7Au3dfdcA26/ugtHB8g4VvfeVuiJWTluooQKp52MB/cZHSZXnyTce4
xRLpmyG0oTZPJCq8nAFQkcPUXI11UJX1rWKe6YmGWyjWEAhqctImI4DnoiydCOVR0G5g3PkjDFBh
789H4p228PUgreZJj0m89yBzEjpM9qx5Dgf6uWTlbUocLLb5uOa5gUhTUWBXdvuv80q2zp5/wkfk
q9B3Vtdc60zr5jAXeK3uFD4WsFNnBwx4A8WkFTwC84NUtZFMEXCIbSmdoM73QCCnZN23x8ITGZQj
F18/chABXxTBg9TXom6Hr9vJKEAnVaTq2M7mxER1uCu3GR5grQyhgkkTmvNh3IRz9qMcBcccrEiG
v602eRv9pWA2dMdqHd9y1lYfqkTm6iOlXAzfTsFqngMOa9hF8gcNqvEPIXN6on3EWVYCzvsSXBM6
xodxoDWdmq+wvaxWqQDB17Qo0qOHc0ym8056upUn7PheCHD20Chzi1Doih+1aoYkdlTnYSwdgMfo
zpGqOGxsy7Wp73pWvR+iKyuTooKxHzjpFYlreZdDuHAVj90amK0EkrZZLzZnyMmXCqosfAFJWGrB
5dE0UMQC7JwLRBuCcY8pQXbXb5GgsvNrqp7xFigJ+MjXvyzEUtfdD6LZpEQJaoy7jMC8zouF0nCT
moJOy/zPh5Tjxtknfy8mSLw1NgUcObHDcHNHcdcHVEEhG9edIXQK4Owar5xNX16lsUgorCWjX3BK
yKbZRoFObL/gAGOGPg+D8tI76RFWU+f92F7+MxJTDI26WdqyFfkvZnmVqTC1l2NJkygmw+01joEG
lRCnQoJgu0wMu1KiKN0jmiW2K2AvZqVyWNf10mUPHUdPudALZ5oA/KReI6Vuy+CkXykfJMAdH9mR
bL22OXRscEoc097m7lIvo0HkSOrIg+rp9VdVJIHxcxqkDxJ7tRKc8EXKgBPCpdu3Zmd1PKioIpco
9cAe37Afk6JNs/0NfvYKzS4DYjdSDD8/pvM3NBe3V3Or9PfxMNluoqbIkKXhCPcOy+L75yG44tQK
7VTFbt11rTBtP+5f9pxVQJNEciLFjKwAAVr9cnZutF060u2+aJ5CxDJU2/TTUSkRY9pHbuB3xwsD
WZdLwkXXnv8LomGt0CgwXzk3S/md5pxvXWmGH9+7qpmFTPWJ/QkOYthkKVjyQkdGJ6kgjbU0sp6J
UmRHKratoFG6ohzL4EJ3o98YSLLly0IEEBptVzr8M8u3NSaPPFReOHq3cwJPY8TD9vaaNRHcP7uR
9SvChoKkvPsu2zADD+H7RTOXblcz6OQRlGEyDuC36+MH/4GV9tLETAUrhZeSaE8XfeRS5iVI/CFN
PK5HhSUvK63kevqZWul6HE2CreO9awKsFXAg1vRpeU1AyrGw7JmUijG5hWhWQFQwcZLHJ22gnCHJ
QBvg4aqY7zN4o+4bRTmIJdT4Ip5v0MP4cf4zXwoLB+wgoOJwSM3E5+oGr4aS6hsOlQBC0pYZgCjb
qrESzUqYFC/BCUHu1MkdnpHQcWuv1JgmiNTMEL5MO14XQpg0CZqF9UJMALLer0Xm/+0FuU9L41FC
U20ui9kRBY0uvL0KEagAwgTjaZ4vk2FOmj+8WLhzCGzDQ93LYr54mL7DxmKuVaNqPnU48OAliCrZ
+C6ADYutc6v/XSDjRLa1Tz9XgT2H3subEl3StTqGRYotDMV/dbPgiXybynB47hVg40EuuGq/ysrB
fXBckMsnkRtY0RbZv2i3YTC1fjkmJBzmytGftYGvxKHpI33xf69qZ3ChYkOu5AzcpkDhSK3aV5b2
ez4T0JObJlK5Tx3tfAWpzLM2OuAB1SV8+bSnD4f8OgdjC2RpTtny1g8mYp87EnbktmsI6BtmeHLf
atd5TXFQ5V+5HsKeAGwTvMFqCJL/hrLU8mfkfL/2JsHtpzCg5bAavgdCtSsEoGtmo8hOMd8o0dGL
owMJXxHXYHUv9l7e0wFXzws5TnwQVGbOGCeIcRFwbakLeTWBgjO86W6nPWjPPjojKSZgy3NH4MqX
OCACIUHeY8PJXTMUPyuyVTQBc/tyOdcRvJWDwKg9Bkyy6ZgKxUMCmg8DkVt+Tb8WP2d35KXat1MJ
lgm3sOBqwWQHuteAAHkLKepKZCy+tPFV+9AnzrKGLvvbFEhg2aZ44U8bup7s5LzIBTCFlaiJjCfk
Ane/Gmr9xOvm4ZXfa2p+w612RTK9iLw7FaF7fmjNM03l5Z55cCGWJJhsJNo9s+OQkF0VrTdctij2
ZWkotgCTxzC7x8Gf6jwjDY3mRZq/QdVWUKwXkB/Al1M9YBxnZ3vZT2oAdJL9E1rbx7KQ7G2mcXPx
uFCur65pPoj1UpBBFiXwvqwtAw3QD+GuwXy5j6viwUaP6emG25IQulXB/zMNjxsXji9NjmqmyewE
9HhB6xZd5YxQGnJaWuPCHduBaVXuW4Slj31zempQ7URGNuiy0yt3doSiGE10/oaAWx40cZGnsOU+
ruuto5JnNY2o92rnH90ybAfI72kgPMyFrSbttH56uw6drV8yCu+1AUd3qvkZv43yiaiDSNM+IQGn
cKLksaacoHaDbCoJyPVc5OOcJwCW9wxMMTuejiMzCcDIWdngY/UQPPdU3I8xIfHwHFfzdaTNBHod
ZoaOUXcr6kKkQeK8f+HBjwyOsa9E6BFjkgbdap0jRQxITi6bVFWf4zjmiDYdQdPSzrQ5jPQiKXXB
eMoKJpCYnVXySyU2xiLhIlqkfKTdylmIy+MqR8UUVIMOoi/Htq4/rc8/YbusDV3Vgz2s/lE6Gr8/
5e9Zj94nioQ8dAY2fgWOV2MLbc0AlhoAuamJ6Nb4FF7j6aH7WQzkdPNmQ7g9hYnTgRrDzJqtDY4o
vyJtzR14GGZ2bP5legpHJanTnqW979U+XE8db3ds39TWIZ4ndio4Vj7mC+SoADRyHNQHS8ReEIoL
b+lrstE33a1Cb895XxSzKZ1S2zZQTFggR22rJeK6722gL0YjkaOu0uQcCXt4v+P/CBb9OlI6t0s8
gdeDWxeJumO4JZaVPWenDAt3JY33aUv5/MTRaMhlH2GndK3Dm/4oV314QxbK3LrYYKnJ40q2bPYk
P+1nXy9nBGfjqrR0TFil//4aWXcD6+QaDU9sOk0NERP1O4kV8Ty9FJvgcFvimHepidjv/0dXb78J
s+n0ufy3o7H38q9xB7NTfNFNULb69U0bPEUoBSosdnej+grZ+xm3gB4MkSIvuV048rl5POFVF6Ko
UeK0VD0GkvJNFlca03jDzeiPKiUZtIW3zb07QrUwKJGzxx+BBeKi1nISorBvTTnW9bk3kVxOrLBT
Vf6iHBrBhuU7z3G0umsT4nhg/HgNB/9xTv9mCAvwdDAmavt51KiK/jefh6Ki6z5eYzZ+PG1J7YRn
3sZIpRALxXysd7sUYZeyeWWTT1rlkXGTMcPGoy/eg11gywqLCt7e8FjOx/NH91AqCMFl1poGYIFJ
oAzjh/Os4DcjEf8L3y/oval0USeGawXCqkr0+a2RsOZ5t82CF0y9/xkC1ENAF0d6OxYXFPAv/FbX
g0QXUgdYHerZ4NKJnofOwMCU1bRQ0Zw2t2RYa0Rt6ZLFfMlBkmDKcjQ2qvNtM5xid4nC0ynx1/bg
RhCKvZhZ2TP6FYlhfHRiyj29epbsgxNHEJJx3Ox1iow56GJrJHyZx9rdFoL7ZHzBphA93HeyiEEa
cvhZbkxld3MCHms7Bdel8jfpHWux/5XvHNUOiAWk5FHXVO1Y/PgPvkB8aOE2zfdKQsputsrVdL0r
MkaS5wANJF/GpWe9LI0jI67xTmhhzY/3n2w/46ZhKCa5QVpXcf1U8iBvkrvMgTG0LxwP7kRgq5CY
S+3MWV6WRew5ae0PmkqAipASpVwkw5Rhd/rtQCQsLCsG1nmTOs+UmrQE4BVnFGR1a2hLLXn0zLMi
qcixBX5PLkS/40ZLT22ePsV6mjKiH3DdqSvb/HD0h7NtRYBsgZY5M/uwJ+mYPfKntZ9/lAX/yyuW
VB2hLo3gkbnE4YZqHz+XStOoJSJ+lQroC3vJ2DGsvvl6nV1eEs/iizYhv0+3BE6K9WWJ4gSDXiNK
Bdtuv0Jwtml49vq0+VAFRS83aq5ufxAjq/7tWlC+1eV6tvqDL3qa0uXCUJ178zebaEHb2zPsviqq
Jynb+QBNInAXoGXL6HN6EaoGDnmNWWEpSfQYEIl7RmgA5+RA7A3/iU+xmYjZDvlZkitcz3qjLBMN
DaZZE405+wGpY0TZUdW5kXMvy9Hmy4VsHsAPeiH2X9aTBIuo85KsYXx6Qr/Jg62MVt4UHIOA8LWw
/wdRw8DJVNFurF92pbTVs1OsqEJxsGpFExKqLNwCqjJWUaZCvAJhLh5RbmkpeJBSda+Z0HZO2f4+
AH7BJGpDE2kZrhuyAe2z5QQMPbpSEPVy6dKkKHwhB/2pmKpXXEUIeO4HnQiQo+GJDEfzSY34AVZ1
CBOWMEx8xlWQ69/2k97Lf57XCwrjpkEbhzK5jkMT54IVv9pRtl5bGRtdLWnJmS9a6YOsXBt7JqBz
9ipFsh3Kn59LrZTH6RDQQfY8ykp3SeWZjHJ7XMk24xXvAROSzohnuOJ6LwTONw8g3HG8DU5F4gl7
zN6XE8eIZ+6Ks0+t9NTfB6/FAIVi42FLx/9QJ+L7RFTHrOtlQRF3AkrRp0X5arCBKsfDvjxQA3Hc
3AzFSAITaWuzxg7JJFo2q68WZQ8W7J91KATdWyqwKUy3bmmJhamIooSd6gY6T2SFOJiHr4cdMUa2
3JJyaiXune+B4sV/JLGFZPV7b+dJ5TSYMc6nap/30daR7P/JZoCWlMfq5tXBHQPZ1KA0uGmNF5Ec
oO0iqXtZWdMSqtlJDutB/rZsJRu7+buQxpvUsEig6HuA/cD5Ys9eTaD7rqYPOCo7IefkiucKDQ07
pRLrlzWknK3Jbi/1j7Pn6kb94fh03Fo4HCihIdwo9EM98Rxe/Pcj1lCGMa+SIRFIzWOL4xx40R63
TwEAgBRhYI6Ij/Wx3uOIC9QdYv1eqZCAm+CLJuHu+krjqwohkJEDIan4+JWZJFJl5Lg3+wc1hlfF
3YOPS6aCIKejNiVWk1RFrx3WGDcgnj0Rv1UwodNqeWq+M+w87zqKrpMkLJ+HyzeZwgbV2N/Vqmm+
eVCc9byb4lEkX98lP6hrUnC2UGbVANK2Ug9Qo85ykaNQ7yTQLXZE8a5ExIiheudnmiS1MnrrU4Su
AiBHuuQi9llb4P1YgIWqkbiuGqpJkHQximIbZNFXM5mE47wqh7JYVa9Mxtd3eIug3oZejSNArq1d
qjzDEVZZR04m2CnS2CARIQR/N3+nOLmtYc8v3WVOxRmrFqJZA/QpGVTwML5fXdyS7pAqI1/+MrCO
T3Obr/s8YE+DGCYs3XLNn6c2OHrzW724MmCekwrnhUJQNRAd61w9tCJCCAw3Z1fqxQo+HhIt5XuC
d971iGo+Rvj1CdHkYtXPgrzlm8qD7WiirXGgQIB2dtL8Yj8pJ6wlQjIBcdnsyCw8evZkqT/CiTZq
Fx5uf/6pHhZ05NmYeY3VcsSmVfY1tQ6Y5LodiVRGde9Puhgj57BK0VCb536p+gy+x/5KmJDWZi4t
EJ9ci/BqxVUUUnVt2CNDi7x6m1L3v9kqorByoZpTfmkgnucDR+J7xgxx+khHUkHIhqADC91XD242
m9ljZKQkO1VLSi2wj33dE3mLAyfXTzcLnYxzojHeCCGfDEHBJMNeeB/kDHW9hCva7UzBdTinOC56
MruvrWFp6dbXPuV7ryZnsKMp2nCLNDc32pbRCpd8wUaZhiwzidbFfmCTzn2aPjZVu9wc/La4O+9T
4KY9CQXDnaKEJNNB7o0cIqpY7ksKyiP/Z8ksjTJhPzDYjVpzt2AzEuvGdohbjOHLYD83CtauPpWC
GKkl6OaEyKvBwUrnGo6YYq2Ao8sh7NiXG8GnKya0QAs8xp0rmr6Ly9V3f79hTZM5za4Orh63lpY0
gU2ZKP8F2wt937Mpvdp3Vyo+QpgC+J9C7/Z4N2ydKIWn3w27PFAtvqh0rdyAl8YdoVcpuyCVQ3tH
fbCt9dgbm4cUubOvTBSd14OTET041ElPfU/aKcIHpu2W8raSpmzA+/cMDTcaiFhkSGekbWldhaDE
uD+IX0TFvg70rB91+x0JXyDKtZhf4sAyCtF4oZChhoYwV+L4WPhFx0ylBl5z0nSMikI5rwTU1//+
bPqua1YVo6Tsvx9ENVcBLyAyY/oKqw7JUG1tEyhDBMq41dyLIL+gblO51GNQp3y8JdEflBsowp1A
RbkOM3gMSn6YfLkuMIbhPvXll4RKwgt5vweWB5cnZzxhhFnJibB5z1H0SHBgGPEu7Pe7dCDXk+FZ
E5lQ1Dt7EDOH6DPpoz5zB2Tnq6oy0/JyFrazWq497aMLjzMdAbMewbNAsxwZMFWYjoaPu4KULhoC
Tf8U0raot2IwnYnbd+GtBdHzdeJyzCtD+6me5qV6BHXnSzh88WgYcgGPeAvIag25HNthcaQJMG1N
Nicf1bT8HknItT1SRI17A6RpSleAocTStPYlifro2Exp3ARIj5i53UtI3vAfgZln5/efpAPWui9d
OJJPxD3woNpTIaTYb5Mx82Rrnuc3i5u0b3xYE69pMfAfoIJJqOHPItwKVA+C70xNmT1lDtyTkDur
bi0eQzqsWDYYqFwDtGfVzzjOhNjOC8eupr8XzX2hb8SZnSnlVhYlmdBFDBQWgI0CU6jwYcGf7+PC
76wKpxpuGFmHzK6XUGVdvvKOrfVo3cEm+rojWzMjBHpCl2XHwjJxS5p1xuv5XKZjc769LR+6YUuT
lRqgmOrCBJoSstMB2g8KVWI5viKsu+7+2OiKQ87hrkcrIr6gQIneT0vsrB1PPwRvRF5+TM6fVBNU
VPj4ZuJcYRTbWumcKW2HANxT8wE3fkbmMg8zlQSKStrTX9Zcn6pKR3TPHoKlTkVJingjpInmzaV2
WnVIClCB89Rqd4YliciKlvF/C3zBPDZgq8afQjJkl0Pu5HYDgjZN5Dql2Re9vRbxEl0wDdHOUR7c
iy0TrThOWyNr1/cOHlGpNqSHfyED0cjz2m51BKCdIQuF1mkIY91LZsMoXj8IWZGqLCWbu94tTKgE
65yKHF2MUury8pj07f/HrHmBCwuKS6+LurI6peH8qmoQO/jRYsly6uT4MU8UEQ3dH8Qjr7rX2AMj
m1ZJXuoc7rea8o4WkEyPIHMNKBAUwy2yDEohu3q6zoysp/+cGTfiS2TfYm7pji7i10va1I6YvuYf
I/IfFI6+PNHrysOv7BY/0ptJ7J6mq60+73l9G0HYUNUGoMRN5vCBCnA9NhFiSkRtcwDtrEgF6/p4
trWoZ3zEZDEIcHFzgrc1WV6Tnkw/miUYcWEgvgCVlh7Aam+r3NLm5xmbQjRyGV/8wvg2W5jKomiv
fQ8+HnAxRljMcj2vwxkeN8sTIqGvS4yPyFuXODz0Pk4SyicqduDe+fxbQ3eMLYaUdYj9BxqWBPGH
MrJ9xSDUITwsxSTZ9t6ckXe8Ql5gNwP1+SqqNLiOWpXU9DnXHuNsrwD8w+6tH4CvXpLfOSr1wwbG
yvu0FMnCb1WYHloex2PhhLa4GUUtXaG9n7M7oJ2P8+w6b+Jbbbod7KKEv4W/2KQzPKXpGhM5MOag
D/ZLWTYwBnLvTjb9dR+ff3rhdg4qbV2lSOrhDMtn2fIA9fCikSC+JOPi2kFCMlZWavDiOLUjiOCK
qeIm+qCCuZqo0HpRKzeKEjgFcm8tlCB29ccbFYvhq09679xg8/LvtjDJmSdDCzfv6DKiqHUk5UJA
IFU/2WvDFWcM0JlUSOJJvMNnZXlRZyIgI+qi7rwgC4ZGERDKFPWaK49pOX0VsPvoNShXjZOdoeJY
xR5XsP2gzaxJfLmdThwahna68pXrbR2gTtSWJyr9Var2fzyyoVvIuI74iFkK8I+4d5NVWg5O10W0
HB8uF/2OwNLmeeoh9ZTc2Jcn4fyK+4YSEMdbSYZxybrqwSpX2/+eZD4Uc9z0BrPG9eIPgbpjcCmm
WawcbUCBVOqdfg4r58xAVRBtwO/4aGDQw/9tzV4p7W6CeZ+Qkw3jCVLKDb/Z8I4dMuWVMfwSc/CS
GuiC0wk1e9SY5SNUg2N4lkF/HEfoMTH0HeuBBFw6jIcQp7zJqhlfqqSLaFlD7+vWmKr1z+b96xBe
w9MtehPyn4Rm0lSbVY1hGcWzpYK7qyhV6aaLErs0rmk4xSMN0Qad625oh++SHk3D2N89ay8iRaFJ
JTe3Idfkuu5FQJVd6x3jSvK2xPfF/gGEWMfxxoWkmkW2WoPToHIM02XmxcYZyV6zmrZUUAeMOlTa
Z7910hV0Z4cIej1A7k0to2FB+mUCFvkbU+jyPqzTmVh572tc6XuXehl87hiz2JWQ9kNQK30ZChOl
6gP9+Tu4HJ8WBy2GdF2PRGwYaUaKMlCVsGsmQUJBtj0UHCshopxfTzzi64uUR4LoKshf5b0SHO0v
rxhpB6QchCye/VtCL3WLk1RG9wgMyGCV2wjDhNjEARa8dAnTSd1g3BW5yrdDU8XXsRVSDYuspLWP
fJwsBKjKlbAcXZHNAzvoZcFhjs5/0Vbe2qBXo+UtwYCM40oXD+zzcaTgCD5mK0rsKyHrPom1AtSj
YImtCHKSXdybJvQdJtUMGI25AJv6pYzZvbPKbW+hiqGVr0/IGEzTYSyF16WiKdgid39//h0FvW0J
mwglnFgGbsitQZHzaBg/6EW8JPXyfmyrhCJ3Dcwm50VFgahUH+WYy4ndzRbe6B6TeQOpc3of42NX
xQxF+auSZwuP+8EBkCw2d1n0mJ7T/sVOPPdFYNaogMfSiEmd5EwFbd3V9ZF/6X7qOYKeX/QpDuPX
iuv3sFBZgINsbaPtzYGwOx+9I26SNAKvf31wtyt/ItJS28/be11o4GBGeZLgx2NEIzocbgifJZWB
ohp5gmKG9Xbc0W5ry0Rg3he2jwDqgV2zmeLw5BM2HgGrhzpWI5j8Po/nF7tD/WoWBX2BGAEHc6Y/
I1nbMwiR3IwmzYpBS08OL0j7ojpjeT2fbp7aZ4ZYlIJlupqXkqfYBHhAPZVoLD1FBnW2nmfrICKP
0EdyoZ9BE+pqlRu4EZ+mrDJPGbhGjDryzwTdl8SuwkiMGiFv0Beik1dWLIC954XJyIH4Y6diY8n1
q5VKrLtOUxWVzP3FHdjSoT+7bHqnJ5+kp3VmDHjlVMFypE9D1NimuwRvKYAbewc72bQp/CrHsSwa
CC62LMgZHz7F7QvQDChYz+9Mt9NH/Ga2l8cQ7XWQgKYOY7v+zQko6+DiFjEGswaq8PJ+obpZF67n
CIVTn4GbGGBXersNYq8H9SJAgs88KQVPe1cQve/0q3Pn4zhA9TnpAapcFtmfpJJ6Zz5syRzcaR4/
RIso0NPSYBfGs1BEEPRh3DCcUikhDZj9soLupQYmKdM8MVf9GEaojRdae5mtKa06zh9OEvZKZyZf
E38S/t2wxsjcaGJWCH4zVuLDOzEN8ITjyjruIMIj1GffnKt6Xgn/Msj8B7ephivIcZMazGs/ZnmW
7xpSHCRHFnc9SmYrQsJVumAHCG8Dcg4QmBPPHmR0CXGVk6zPQTj7BiNakG3Yv65xLxEsRElbAAv0
jsolQljfUaNRLQhPpmt2W5uhid++eV4sWfTq92WFQ/28RTgDQMP5SCNLOHxofN+gnB578urcpYAa
bBk1ooBp7Mk7I5Sqfyw95Dg+nFuBR4j/D2vC/B/4DEk+PvtbTX1BWKQ82/Oj47+qVhvKWxWyLODR
1UBmN8ux9YDFzpSOZu3s2uPhQOf876kev2sw2YQJN6XWAGr9RpMqVu0Glx0CyZ5JN0fQHA+dmDkl
iJzypkJ7SBHHPXk0R4BejgmbNOTEGHX1vqYfSkCJg1a8s5nhm4ICu1fuwo5I5Lb/nWSQoulZ9CZF
l8AoYQXn7E/dcrYLmpn1HvjTW5e9leTLLTt53T7++UAuAHNerIboo2+JxB3nEe5BIkegtfb4Qops
g2NKUsKLOCVY/1v6O7BHBTaWe/5+TyUpJafj/cMLpisaz7JolqdSVJajiBPhVgxNG4LfT8r+Ua8U
FajHxPxYkKpHGEVgbDQ0tpNdCQ0NZ74awt1celfkfAY70yrYuJSvJtvx2B7PDY0m+JyRRnXWBw9e
V+NHaTNzCZUY4sPL212p0t3J530KXYNwyd20C/KxXgoRJluihAGHzJlLWN6ZuvDvAHhaHNufdzFQ
GWc15GNvP9g5OVf0AKEGpO+XaBOC5qB+DnKID7IeesTEyuqK6L3a5HlfYL8mjdprXHxwnTaGuSzd
5afkU0P9CIr/1IZn45hdAcXJyjXfm2wQqSbhEIEYnnu9rP0chqhGcKQj/pSFo7coXYfuIyYrTUiN
BkRWTCrTNrbhUjV0Yx9pABbX4WWETH/pij4BCk4zy9TgzLntztM16og0LtsR40hXKcm8E3z40Ue7
fxxBW3S8Ddo2lzRxD5sLDSB6MU4lJeXmnQVIc+avnCX1oAhbT7gH7HigjbDNOhiNXbZzPgea5etz
lE5KSZyxsl+L7Hq/UbclT+VMwvzHo+QM6cgLp4c4AzMLk3d1nZd6h1sSBehEtx8KG9ky3AfRMo5c
ZytUDSrEK7H74/mNycWZdLfHGFyo4Lh/IQyGs8lrK87GOc7o+7k/jXGRzM4OuJ2a+AAVBB7BhIBH
3nfqC1jBMCEFQdfb2i6uEllikjFclGXgsjuelRmRs9SPYp1APymMu6BtyyLRKjVvBA9sEsDq799B
QkrYuXcg4D8f7gq7C3otgTKzm1r8TI2eFVgcsmFMe+fl3D0S49J8ZTy4LipJN7T/J1th7JARQIxJ
xrZnDr6C3nH3941ARolvx61O9NpvrB5Xl2nqlPc5tIB1pfIUimpEofDcCiccYLGZlR9ACCrrVXS7
31S844EnEgJYptgopreByDkmHK2DdB4g92m4qp3t5ecnoKhiyW5ryaT2W9zCgstWiSR8b6b5eWGd
07ZXUX/EUhn82UBi3iX5+JQyfIAxXxGhHAm4fx1YZw92wOPBqtesEFaOG+7Rt0pJRSlDzrIqA6/p
ZIo0ueoTLGEcVWV6SnWYPgrX100jqPalfOUvRuKkOwmV4Z3mbQN0Tbp+aT+CoUk60ZIBX/qSezCO
DgkRnCjBOIstMqoVBFYDiQWbOKPVlvN7rVRet/S8sPuaF8y0OnQfoHDpaIKFV+s1FjvZHn26HX+I
t4nGiCGksOG1X169ZU1RwZrh6W2IOpMIBKuy2DYrYoHQEd/7OgYHCA+v9byZqvyOGRHvAaoduXU1
NPr6pM5u/xUb+wC27PhG0gFDG8bI5iYUrP9UrAQFbiq1vrf3UQZLKNnq2XAylJOETO6UN1jOL76N
ggcNPrGcSwo85JGGSJ1eClZnKf5KOygkn+qrzLf4wB2jgbEiRtywVYAlU6/YwS7UznHz+pigUfw6
qpeQhUkOr26P6sVo05MN/E58FPLwLEfKggM+sAdlyUpKm1doTZsRfxYxz8/zbr597hLM1+YLmXx/
dX59QSK78wprg0T0mOlGwqt81cWKsZtm6WrkAJgQFJpTZ2YLmvg9vEuW5hDPlIISjNZC0s90cfg6
G1RO4nXdU0nfQ4yRjt4hFAvpFJ1yRTSbI39/3KWaTNuLVf2zqS1q2k+xqoJeDX4NRhZ4eroDKRAS
neXI7D0POsyQHrvQm0jyUldezSntpBgpPCmrbhdSVLy0nc4Q37KBONNWSgLgB/P0wWwyPVdvkzUU
Igq1DOSbwJRNQ1a8zFFeB3Q8NtpKz2yeD8UvV3c/+WNZZf4vNsn/Gf7g3Jmhnnt7HDi04roFZPop
t6kQn25y1Xe7oGSNp46ou/1tawp2qxngz3pEXz6bII4O2PukOw8XufIkgUkfzrfKLAcwW5YD36dc
7aPiT4/NeV8pPAsYzF0ZHeHIjbYnyqDA+1H7rAw8IimmXE63+2X6p3wBH+oaMQ8oIU+n4f9iOMvf
8eu4ldmBdXwKJcli48ticaQUtRC3qeKjqyZ8rjx/F9gnYuZNntRheaCZb4JUby0t1NSoAYDST939
diZ6tknE6dtqCXlznnHRqpOg10StqYWuPLQ+OjB5dZGq1K2o5jbf2qtSelJDkgcu/3bMAJI6rA/9
E5UAcvfYJx9VAATWl3A7l1GSu1I9FIv9jtUtorOyTTjY8mJpzMhk7QgA6PXd1B/81DEw+02s5Z3V
zgwQ3qFtnt54/tjS0/y/uQwNrnog0v56BiyGYUq0W1Zija8u+l6/x+i9TKqByNTDeK+udwO0YzPn
6SlR4/IE9Fckrr/C9/baAZM+6WJbZYoc0yT0xImm+vc4pPv3y9WDn6AlLPolvHlnvWWrmJiYnUOz
mpTvpgsfkYH+xFbaoWBFDslQNt+j633cTgZW+DanjhbOGU4z0TF5VEPkjciB9yc/mrKAfbJjwiEI
TaAGXQW5fhqubWUszupNsFfqOHNjdvrcLLzthf0L3fbKcCIR/MI+x28NE2mMcN1KvvKiJe4F90VN
4PDtLe6655LVAiv18O3m79kKRsvdxhabrAOG1KLSZf0F/Z9zwlwSaJkapPhHrjyQfxaspKEl13T3
AuDZXCmKSdE3a6/uA/LvgglhqLqh+vKvoYkVyqAW2wJmwpPk1GnRA70TXFdIrv1fF0oZzf9UYOmC
fZT6iuDBwvWx7xjqPotKCz9fiJOwj0ZpIUc4b8UBkOV1RS0ixXu+pigt7qjCJWF7xLoKWhEuF8Fq
UULE2b+P2ndui/ad1p1R7Y4uHPnFVgf7AxdcKeDWgH8IdcyZj7mv5SIcVmc4AR4qT9IpGRfNTAGr
jTuT5wtP++dpQCEkyrSNiy4yqkwlzCTJBKVkZMdYRGpgxKJhuuu1BNlMUBRkpyrhsxm3qNhG1sQD
hqjI+MCDsbDqRLS1zmzK7y3niDW9tIXWTLXOcjBPOtNbDTjht/+uPXD6viIMIv6VdqFR/xBYpGaS
UVHsq111+/a7KW4OsbeWelIkSJ+b+0+HbC11r/8SLZ6HJF6FhoQOglhChdrM5gcyRAQXvf8Kz/RU
m0TiVG1KDOc1HZzAu3aVLvjcxV/6ztWNNOlQM41D2ItNBdJVmJILv59HpHukdGxZjbvUbgKlsZkD
T8qGc/RuYmXSIkKpj6PW8bKOulmFHk1LflrgMwx5+CPubFOTLesG0aESiUc+TQVacb5/qZlMlKEg
9uegFBWYgjgOVBd6+n55/eAn5kmoVGsoU8lpPj3IeHuFn0sttDlsoy2S9hHtIxpSiEGGJhMtdCUs
Uvv3GViAuaYtbevxs8S3EPV6zA/prSVHmpVSgYoBkvxDttoDss0YN3/08s/2xXaUL9zJI5BsmB3E
1yGBmX5abjtIsbJCSWnfPsGiD3GIK9YkH631nPgt5+P85vMJ9e/UTSnbgTG2NLdSt4rYZMtRm00x
kskmr4J8dM5N0TRkBJBgrBCICI0IeKt8bZzb3VPWO3lO/BN172o8Yewc//+DzirJxpF5Fo2rkYrm
siJ7KNq5fnyOqo3EMmcsUWioQbR4EQP/Z2FB1aRUSM928C7B/p+GEeIm9uu/317TYUZPUFC/LxBn
aGeOqN6jVIKrR+3HFBtDOr5xxXhkTDPCN2/tV7G1k7+b0P11BCw9QgwQxE4iyH16lr0/FOUW+bNO
9AHJtqZx90Qm1eoBgS2GB4ve8SOZQ0/CnKz3/XSXykm9a8Gwdz1OgH2ukQDnw6ZPCP61j81W1Fhl
nBM3O1vxexTgi4mc6bzwueIr89xVZ/jTHtxhcKrZswRSHumqdoQWO1CmXHnFE2xPjOj/VbEo50A2
ob0vYHEjvv53+TeYYR+Eo6TQy4NUOI/pCn33wlv8IS7AZEIKGQ+aXag7IJgkiUBWN3Yfmv/8Ea0n
gHxJC7PZYjoGJiSl3GbQ+5I50vIoyvVDwb+HS6LueRgIznlkJJDwPvIvTCqnWRg8zLeBLMusqL9n
me6DTUIZqkCL+F1/ZILg43n4CHeZGhoHFPEMt2Hmd3lUONVR7LM/vyN0h+5yXNDjdjzy52raGewi
PoZsFLn9FD6riikrqP7ezdA3qgWtiIr2bTIM0jef6xRY4aZQ3dWQY4DI31Lu2eE9Qk5NYBRjX58X
rl3Vlva9jsPPjaqvyMMGqceHkAS5bfnSaSpOlwMNiZdnipltOe/8u3zMN9w8UA73KbNyvYNQW1cX
R3eFsFhqnCTACRQx07+2dv8ddjTS7RnYsqJ5AJcvQrdCaOveM1n/9elUu9yVGGBD/6BlAjDZnQTR
EG67AO9x4+SXa+15c0euKah19/daj/lUYqcdCxqgEo3ddboWWuzRwINBvVdTa0iwiMn+rpYWUwkV
x9EAA6zUi3Rr6AxIYZbZXHMDJkpoG7NSZjKvQMQc9Uuo0TVMfVp/EkstlqfzWhbAmBDB15fZ8n9k
qN0uuUtBEx4YN844BRC+YWMKG0ONp+jNV1yPCgFlRCAxMSFp7+/NiIQqGnBUrZPF4cr80zOMwrPn
VZJsmj21WXlxDnlPzfwkLLZT1zn95KNkk4klxcykia26ArYUyNb6obgfcMbyxRnsJtaxj0U+IPZl
ZTjvtuGFUnBk+dTb91Kuz3+qLsQHBjaeypj5+5FWjBDOs8j77zEYtt/63S7kvJhdwLOtOr8X2zUM
oql0vzaOmdfOX04vad5382g0GGhfhbxUqEDP6beAbn1Gg0es9T+CwQQCka2SsCsLlYXGFKu6WFtb
bFXytrC6iWEIH94VTqtTMyud/iXw31qSJhj6wN4wVsEizfV8g24tAQLR97uMWFqIlfw1WIjf/nAv
mcNzjfe0XN2ma9UDtjwfvBHcrkqRpoJDvvOV3LDCsFmcOD4rVjutB/eyinJOTDUSb0JA/E8kjDs7
hKQJlOWE3t997zSXasvtWn07sgr0ZDOMbDtFUvR8yIBqCLulgzZhbTrVskXQ5WjfFTbwLBJ0xYAG
jYp60DG+ltlYHHTom5sShDUFEOcmBgFrziQmcFfbzKwpgbKc9gKoYJL2s03Ih/ZDadvtOi0BUzjY
RGaIyDyw572U36lUKv/0wcY15NAZY56XDlz06WNhfqoayfOkRG3uNbIsNHobZfzXUc9whQP7XnYY
QvWFDGbQOAbF9+Dit46tkiYWK8n9PL6MIcTKwKx6XIo9S1ciQ4XAkV3+mhu7P3mdH6FzJAXkj07D
pYKUihJg5BwjG20awecwHI+IZqdCabbEyiKfc3vkR6aPNA85FkMGq4oS5qd7kv0Oybn42BCzuYvR
2QiaoCtQ81L7bVQ+KnhOogX4PweiQyurNVlFaUM/vaP0didRhsoPAPtT/83V7QbhswxVRbQRWg42
cPyBd48oO+dTGCH4+efmNzxulI2/zwwMoZqti3DfVwl3ZXPVn10+WQmdDSrNSl1kDPdxkO5f/C4q
pgTvWESaUEWfbsd8Mn+br36vlUabgXGdSHYB/QIoeUWQL/u0rn/c5NNWxOJ0GAWu20kkxVP3DT9u
ZRCrrxGbdS8QPnwLoFOwFkSDY0q++cl7NixlIH5XAbkdtl0h0tH67D2HETfH3EWKGTNpptg1Fhi2
Jy+FkbzPKyoCMLOKCI+i6GQuJgf6VoO/hTk4QPMfuX3sdcMTaXtdEj+pAAkRNRyWCthntMbBBH/K
PMGUHjyVQrOR/zmp4Is7wGBFSgXrg/ojPV5DxXjgIjxTtC8q0vtXrCAiU9E/uT9TLWwGWpB04LZN
1xcVp3RzOR91S3JeD32lDH5DMC/MeuhmRIox4UIMWrvAtO73osfytQpjrK4R52tKYHiLUbma281v
Qd0rxtrljQQX/PuSeAPiyoG7zv0Rhh4YXTPI2GgNlnbbCzq+39TcjQupwHTIpcs4/fKEk2cBIiOA
wZfwbN2WFH+J6MAMStB9+MwKcXc970RshMjal0JH8dEwbqAcz8JcAy3383Cd9f2QvNwyWsWSUfxW
q+iZIpFdS1NIpyMyUg60UFDwYiJgqEAGUQvBBevMYaTnB7uluXROOfHeeom9YeIeK+9nMDRutAd7
+4yBKubixqDpaNGnkSoxP7+0FZCxlYgKEMCxo5xl1jySFX4o0z5ntZhAIbDViY1MyKTWpDOeGa9z
KKz6gVqQ3VjaeKXoVG6yHvd3sf2ilLvDYTOiuTKg5fL6706rQ7MC/IobRVx5L6354WoyGVhIOQMx
BIZfUi7u7yk4z8ROPS9eVnWAglnc1RFBtPA1VkjB97VQsy7z6pFDNCVzAVSBda4ZHm1fyFo8xXgb
iSimplg7HCI8sEe+b/NTGULVOmWC432pmVi9HmF/AgSXiJzbvCyGBCY95x16Cuth7w8TkgjkVY0D
jHNcWNgAs7CIzZFOZRzhhy9W48wD/tOmRNlqwsN935pB9aKtHKi2LX0LFgnOcHBQGyGv4yYGS6YG
uozIh+KxoDy3R0dVbMfFgs2eLqWfwFRQ9d7gUTY8dkc+6u+xkZlOp299G2Aih3ITVmsB1MHg+NQh
eU4mmZlezjbZGu/g04GqY/goV8Tt/c99U7K99sGP4ewVeY/B2cqwmlLa+ZkO56zr8y6jTBVeohIT
+3ZpvCz7O6b+82IckNiAHFvBbW5nGIjGT46Pb7RRWCP8EEwVKd7Yvmd9XC7L8isGMUpQ7DcfH+gH
Mby51vDHFKAE5mpOdlEnsrqkcku6585C+Zga/ch+eaEVA2jPDwNlojqn5hxjiZl64QVcdQA58cxB
bamN+lTGnrYt2p1LCpxqZuJbeSbitEK5b6nHrZv240MApVXYamfjXslSiLRHiXBmREIR3AWnw1IX
eOONkGr+6cImQ4Y73elt5BGWyjK20OgbS6elD4TU8aEOmtK4Idv3/S5Se1sBWeql0TOzZKl+7E98
HQ7oxLKL55ObtdmsX+jSEDaql21Y0iFTeRlxQbVaM/yT8NyplqGSaaPThQUf2HfN17J+mf/8tEdT
NLCcq7F7g9NcjYG9zVHQ7GBv2hQ2y9/MhGWgdFNQtxfNZcXAZwMtf19XK2Cvziy5m2vraQ2MlwOo
teND3+MJspDLLfRzoe86HGENe6O5c/l4sMSD/fn4gBBRvKov+vP9guQ8eBcX3gwdjguUD1vNK//9
5kcW3DcM0PrIaVuZJbiHiaWPlAk0Cifk3G0BaYztq0r+sEvV5tYkXAoEaB9bDZlkS971e67GzaR9
/kkcNRic7r9MmVM3mNtfJmvy69aBDZa+RrnIkmAk6qzvKQAQW98deHl3rQCTZ0MF/ni2s4moaNYS
bIQPmnpwWCMbCtDlyBX1qT2r3v3vIJ4hHKEjxYTzaqrbIdCzrksGuyxYyCDJH4xkpUhUG9GEf1Kq
CdN4TbNTtGTGwdU20QcJMBszWSdHgva5bOG86z2zw20zyLikI2DyQAKi35WzDxfgPiajhZIqGrF1
HQYmaoBUpZkRljD9OevdfySrDZjfvznLYgRBvb49Ni+j4DZKu5Z5nZFQR3Wa8U+KWb33UBLcDSqW
imp471QzLma+GKwSgCUSsJF/Pfw9hchSSXEjkEeqKywQqTsZi/03GE1bqo69Te4WkliNWk6XOvcj
i3xNgTn98OatfXIAvb+dsZCf00LLwMEBOrQIGNA+3Wnsw0WNaVoHVcdNrZs2z0RGFsm4VFWegwlE
aCWuPiO9VyFk5+aE0+TWxAyIkSDsQs8VQyMPusuy331vxgZh8i7pgDC3C+MZT9tsIPqwjaag5Hjy
7XquItULG3l0XC/XtGmzQhWqKXs7gB9q9WQJRO+AWy2qe63h34TSPCdusW/QSVEc62Jnsoj5Zuyx
V4ZmhxugP7HTL7n08vQx7JDNYyD2SbyOLjmsv/Y8epacZxNerdq11CCYTM1o+G4TfXUHASaAlljp
oJYuFp18e/DrQwgU39ggikLKqHth4OhaAh9akH9F15qTZ+g5cMnQUVrwIz/6Ua8juGaKvd/iYFAM
gWKWqJyvxgJ6PfbMitZjdVDrD1uEIUJ/aa6aI1iTDAtS72zILOnr/ATrjxFqX9PDAZ1bOWZoI62d
sX+zVTDZxs04qSBSd9LfCX61oq8fg1T7hJKY+WrObKOCRZWmtvkv3Rf6urMDJ4hYKAiR7nIQ+zRs
GWKub0sVjqvm6j3Xb8D12xSYtj6Fk6TlxUBZOmTn4BvMG+GzI9EYblI202KVKGaRPqLiLYsgqJPQ
FMpYddgFOyWJQvXk8ZwQ0Qs8io4gZ1JF0SCU+uOdwupwSbxbmAzj+oOiVctuAg5uORbAQozXSCVf
3UUpJlo4x/SGyvCuJY3RBY2T56l/15J8dRXAtSHwhtzAyN1TIrd8bAUtXC6BiWvgzR7iT+f+Oi15
xerl4867orKj6MJrFPVEVx3LNShjqXHQqKf1v0fVBgfCVRZii3Lv38qGog3axGFHx3PXbDih9guV
fgL1krRKxL03dvFMR5Bw5WOOiir8/stj+s6EclaHOXKWw0Nc7KFQb6oiTBfMUXyFLGDDn1Ji/Ags
6V7E8tAHeXyTNNVYq0ISqH1KS3Yg9SHJ2IdAcHRVi4d5I/fHGHnavyXVr1t5dQ5AKOVDrMCInccx
rFKDS88ciMuxt1YdBe4v9g7+J7Pz2WE6lh3LQ+elsKxR8QHq6ijvv2dwweyNiyVe85jnrr0wsqS2
+JFRH5iaedkqeIwlmKm0MnVA99trsAizzsMT9B6b3D6glZwqFzGPwT0QXeKFEFD7+cZmcDZEro0i
Ddq/MgWyvBxyJvMVHM7EHC3bPwF31hPMsXZ4jqwbNa1hJN1g9SlV9DooZC0fxNw9610yGEMhqqDg
Ydl0HiHT4sT+R0XehiuVjq6du/L5OJz+Qi1ro7v26HUY600/P6DJGodRzFgnkrX3hffpCviKxuV1
CCHGuZqnCmGJUmLzjbB4xD0Pff+5M4i9W/dmqlLleR1Kn5qSfceEkuefOIiXDzN1RsM8/mm+wz6t
WzMi7RRaGufm9UynKgnGjz4HcwE8ndLJUk8wX8zgmr5WW8qcwBz1tMGKYptOQEkd8CjqrRvU4z4A
Pg+Xx5ccuz5alsGVcmADlV4fEy8EuukRa7aRHKvybG3mIYbGauqIgZ7wn36xiQDC3Ilquiknoebd
POaqsJbJFf18w8sfLgMcGTfF9yX5YY4uOJwxb/1xh7ok0xSo8uAd+svnyZEQv8HUzq+lyrTHoe6w
UHuktADE8thvZ3UyOI2O+Rc5yK/naymQKMWTwt422eFiZOz/DEgHxyAxkw1ZjL4VGofsI2glFCV9
jPwLisuaacSawTg5pW2nVezYtym6sfd6JaBrBhgYLsII3kWsUPNo63gGa/Y9p8eO9kDkO7pE8kQI
5nEBktljxOsNsvAV+/h3KiqdrQnrfKZ+YrbL0L7Do69laOA1cBDZNH5/+2chbvrX11j69hHSl5zx
j7EZIXnr7oQACgHfkMX7ogGSLS6qrviz1+qZHg5MpTR7EV/wpoVVQT0FXZLr7vHrP8k0kjrDpxFB
DKU5ZYWvcjAU3E/Y0VOo1Chs9tmF8hxWfHkMrAt281gcRsm6l1x7fXNB9WVj+0+TUWZVARKTKWJB
yLxSN8ia/dWAkvNYcs/G6X/OwPusL5zPfibslMgZPRukmdWS2iG8kdRrY02j+Cd47GA02ocSgV0I
7tSB5n1NTX8RKftS1U41pb7n0/pEnCe6t3QCLyIHUrGbwDZUssrWJzVLqsulabf2ccLCqXNPwxUx
kzi8buXHzLTOhcv9ayeYcl1nsurUC8eomtgr8+0VaWqH03C9nvm4KZrVncnooc3FrguyehW1VxjZ
uYa5q8dCECDwCfqR050fTRePMdH6B0toy8x8etXJ1kZxpzK0LFNx4f+ETikHrEk5wIuh1GRm7Egw
ePMujP6hF61QywJfdx1v77+cnZ8q6soXHyN3QQMxQ1DcwEFp6nnczYk1s/gslDhJywzHXYmoqZyu
io3GRQhwDA4FYgDzO9fl467OiuslHD1nr/EqkwuqMEJFiyyKorjkxvru1WA/EAN4Aly/2tVYBpK1
o6N2OqW31eFS7KYLTnbpBDzcpWSaICgriDNQ+zuAMEnu0Guv1SqQ7hGV3fZpsIoapXmoW8w4Pk+G
Qo03Dl3PB0+WOB+uQxBN69Gu5mwwN5sqtu3bN/PNQi9IcwHdgZ2Ewa531XA8DVUkw1ploCIDFq/U
MvfNPb2lj8LR3raWyRSwq4fNgOMF3e7b/9mAHB0Fkk+k/12yzMee+Pf8vBBhnt7CRa45ZS2zjmV5
lq+Sb3hx4HZhUledw3SBzq21D4bsBKyRUj6Zzqs2b3hiL3eQ0EspAhlS/srkQQU6jZRmVKCSNaiu
3BBNrARbjXVDW+QXjEieumavt6By2K55sNgvs7MPXPb038gaqtWJTd3ouRF8SUNdkMWGEa4lkUx0
n6QiLqJ1k+rn03fSjhOWOn5tYg/gDIP5CChvOHa1sfytfYYV2RsvhUcgAVCZrs6xAExaiiY3yKDr
t42+rkClKxRJ1HxFOzxuInqVzWH+hnj7IO2+lz3gjhSF8Ez5AQQ0kF5NDaT/VJ1+K29oOSDdMy8d
GIw9hSoY1VPQefageCRRkTpz/frIxUAehow6Ujs2OXYbqrPCLwpb/KEITjIVDaGJH+k7HKxRHkfL
nuZiOkihj12o5M4etWF1UXRXa1FlGu53B0DyVp21SM6BujGSnSL2vHEkJoYNktbQ7CVQUDAJzOP/
mKL+Z0Zp2jRxyf2Hw8J7SLcyZej6KoszDy0yvcx+ib/zhwl9bwZ8Nuj/TNvfRZuhDGPbbkvAj7q2
5PbMEpnJQmsTqh2kRZTFmb9o/8OsQ0y4KsQxo9JQcna1/o+uTIzG27r6gISirUYv7Dc0zonOzJxM
R8cIKl3Wh5xKyLv+PS8z4oJvG0HZFqEWk/EzI+2hgDYy1gki9eou/qqaDVbS/5YIFGKe5Dc9SDGS
Nt8KiI83Z5uOejTWVo+UpWpVtqA6X9uFNIB4IwTVkp5/KTxuZvN4CgKqPBoUfbD60mAcMUyt5Xuv
TkncnuMT3tA94s8C3wJpFveKCAKODHITXODy5YPH2CMOgLk6xDQLbHCLpEwykvGd3zS3fud9v4G8
zyLtCAdYQYHo7t1SGK9dFF9UBvX7q8Q00aJ6b62FIYF+2cDlO/4LLooxrLrWCcH+fFSkx8XOxSLY
iFdJPK9VFi4DkC8PeHdi7CGwagZ3dPZbzKGR9i+W0cB/9I7S7PBM2zZLOj5GfPkDf4ntXKNI0d8h
UdJyccwC+aw9JBH3uzzeXCS3zSoG5ztZQ/EE6GniTEmIla6oPtY6LKLGPPc9U7UHwR1q8Dma2tIj
sSQVtTxQLhWqna6p7cGaidfT1ruQkA+kzxBFyz0vTxcx9ckSwOYCSXV772a53R5qGoo+l+DWXGsA
hVpSoUte2JzOD/woeQl7RhAFIzLyOwev9K7P+5uN96xfX/krWZtK2gCZdoSXDbN3LfPjYWK2QZhn
VmZjPvI0+/P/AXxv489oaSy9yrNQQn/mCQmginOCCAL9A8D5Qs0mtthZXdkRayWqyGdkEGB5lRWf
5vlkE4P3Ojpo4NI29/hxxKbLctHC3NA4EQTCyb9LYWrzo1P1+Px2yCMIV3/VSxyYSogkg1XtvYh7
3d2DpURxxfjGrtH5afsEdSjQXNmr4kbHRlO0rVErewd67iArqNIdGF8osH06gQFl/I73ZLFGORTi
nLXIx3OXVqBq7uWqiKQr/G8GZJh2SGr30zG5+Z4jtHSK/o0QZVUc4yWTRK9LAdbLf2gNNeLUIjhO
UA+HDqW0nG1YNPOGYdlyZb20lg7mmUpiga4Jrb3FrYQpB5seTl8YEOKDNtt/DxWleRiFsqYcpasq
KBsNJg0adzqSt/bAKjO8HhwyDMvB165L5fCvvShUZkxhKibGFhuTYcxb2Rxb5bVCbdSUSmSVtG3N
O0z34Xbcm9vOXT092MapXfIvmoucuEQJrxO32Of4+jMd1/yHbrpwctmNZGONnSOuvvAiJy1F2yFx
8LmIBT25h6kz0IkvRwlP0DnYk+PzG3R6IU9+TKcjhoZup5nEm7aTnsBCI+YY1+IGCKocX8K3ouZU
nSs7cthj+TvZiqyrkT0OJOMlj3CFobEISgz0vYJARxxFwmDear8elXAj3Z1UFjt7fd+Gvp/UiItB
HnEvXJsbRcRK0du9zYMvOYo+Qt7X3H6P1FcqOTzJh5fZZrt/vyzi5pMKbb+no6hGAhIFgbvuGXhd
WpRW/mi5dljJakwsHegHSACCD/fXsYUfNg39AY4KaNk4rIWAsC+8kIqLl98YbnWVmjtmEaw9V8fC
xpHfoJtKQDuce8hXrPpqY/zLYLiHLMaRdkx9CQLdIzwOf3uQD1FUtOCgsh11qqLaFVabh/WQJwgQ
L4f+kRv5NZ/drLhL87hYiK6br1x3eVwE1WuI4eJXxNItC1gxfKI7VfozUjcBSI+CSHEDc3PsTeYs
QiTScoevLicfDr0d+OEcIRHu7MNupmuylNwWpeJwCxnn5DPZx9oahIgGX+RVfNv/kFtUhlt/Ggw/
n8vuIufcerjhfOmgGLJPxjIrIOvj4zksSnH9n07eVATC0BXI9vrb9ub4gU0H3tqMNMk3LUq8zNVX
YCiCJPrey9eAUmejMsl+hkWGEyZ2vfQewdtWBENbE7iE8pUY07s2cLANTGpQIGfkaoTr6HXhROmh
C6prvluVAk/RFVCE69VjDBOXte6DulDP9f7HAi8g0djjZBDDsb/Zgn8b1YQQnRGQla87Do+5Yo4+
2Zs5lIOgfMjLFOGEF+Zk8fEQA8NJhVHwa84qA95jRTR38YgBDE8D0tFRBH+XZ3m2T8bYMyzwIjHi
cZlpwYttDHmWpmGZUYSEqh9dxtvzKBrq21/SJgNjGytEGhUmobSh5uTdfzUkg7tj6r+6strbdERJ
+QVYAlQqWH4o307g6/7/0CjCGUYMQitEOTn8pIF5LC53l03WgSCYwGXN4lFY1Fot34SrMnL3Q50C
g5H1auX8t5fAv+1cCCyzZ7HKcgntCnXGrZCVl9ilrnCBGdiLe55AHjkgepUx1VdjLEFyWabkqtxK
Lqm3ikciJtMc1gDfNeYB7/F0AIWXgD7WkWRcfBB59MjFZX8CH0gUsUSmkyO2CBx/jzfJNUr48WDv
zTxazifYUJd5biSO2qFFYDSOW+tkPe4CokiV8TS3n9gyM9EuY0MMiicgECErg+SEMrlU4y8Fq4SS
9Abf7kz/Ny+gIdrcLKk5nWTXqYm6YG+7WE7fp3WwAw0JPlIq3J1gSuMmKKlLTmdqpJsD+pxSRd88
VdY/+Q3olWosroF1F8LLzYFB2/0AbMRLggvXyp79OopWiUEraJhU+rXryp5lxYiTjh1fjEorSXjk
Fr1OjyZ4y0QX9m4+bm0xZ2flXpvMMyorZA+NqhUEnO1hOP+naom2cX5/zOX7F64KW7wZY1Kwf/hu
/4FI4drNogXWFR9OS0923dNQAw45ASIhzdBnJzi0OF1w47iza/pjzxiXgwe1MnUJJc5ou6iYgwRU
7kmgHj+BXaV1N7zmryQpLH+51Udppz8zcsKzsQFCRPZpJowaNNocDXZnN06N4VWzC8cMeL22cgci
fEFDsXmasoyG53IkCR42uYIFmbzJtefGE6ZDh5nzoIrko60DIf68kGMhGpwpLAfw0hikXzaTncR0
ve+DT/LnIv34r+J2w0GzNQNnIWaeC3iS3Ii3m5ZpRhHHGDTfLvRyng9XrEnvIr7ITMNUxqf7+3QH
SKonTeFy1KCeYVA5/JcXZapfip5wqvu48znYE1lK3AsJ7qiwANq7s0FmeLaYNQcg3abjc0MVTDEH
43di1IUGxcAqvUVa08zW3o+aINxUG0WXIZce8DbpWKkhLrB7/w3GaryP6Oww5xFywkfk8pOjKLzm
cddhMmgLz/kHMhJFQAdQx1P2zkRTWL4yw6ogB+vsFTHIUGRL8IcQq5E5IYF6Jg8QDWXd9hpyMYmJ
knwWkv1oiUK4Ln383dahOmtOVYtsVjRKPMPht3WKOEnfJHGQ5r3KTDE/IqypoonezYjmSstL++Bq
TTnHIjK2+WSHz2q8YFB/Zhmh0oWPHTO141ZBm3w46BY5xTP+DP+TtaSmq/K9dmLtNLY5JoIpGdF7
x3rhouWWyE/JGt9SzxxnozWsJLEB75oUtkSDSvK13SmA8ZVI+CSIa++USVIEWRJdEw9fmtp+Y9wX
k7t2PtvzUYdDEFoRBDxgIWVbJUJ6KJzejoo8P6oZHHcdMyuVTwMywbQDIUMehy/ye1NwTD+ZXhbY
3Tc33TpCdomT0YJAxvG9V4M2gf3sSwSssE7oa01BCJg39E/5zglJyLymik35M/44/Oi/+PaLtUt1
WEs4YHaUpP5IwQm/j8blAu/O+6jAmvN3K+O63JReXkNHOZSsHayofh0njds1QQ2ZcIBDc6UUEoW/
AXbOqnu9XJuRXdS8SygMP8lQhwcRV0jXORjWbA8Qq4sOdtbWiL2lvFT3nSATUKV3dO+hJCEXGUmP
GxkS78QLePcePnl182/1U8Xp0nSuArz6C2BQkaRkQZBN/J2cHBvfLGehOpzmfFzKV5LVc0X1YrMW
MPWk3gm85vegErTc2Ny49+C0Ig11YpsVD4CG48G1h7JLvfUx6UwMMiT12tzEoZ0Bdl1/ErkL8UyC
PXCUUs72VhSy0jCY3h7VOtzWKsT2TmFWUdXn+Ubk8XxB305eQqChHYfZht/6iEc0IvkFLTmAFuNe
xgdglZIrY5ZnvGFPr6waijcz1G+c7GuJJsTMmgUJwzpgqu4L1e7+rXslUPb0sMxnzLfelcnxDMSH
HzU3CzYi0BeUQK0TKf5yWjUciaXV9Pailwzo9Ch/3ebwL5B/od634gqj1tYzXJsm0bhFU17KO1Z9
X4mDFjcIUapVWF8pYsJ53vP7jsjwYsVCJJpvJRLbgGGNT2Oz4firdzGZhC2tbxHwGZ5McjR95078
mV3VzW6F+17c4TH6Pti9eSETMJoq04AtJlK7lFg14kz/gbI+EpawLIkEuaYi2NWq3fDYjsy1RUGX
Z2u4dV9puO77q4rKB7kaUlVfETxqVTrJYQhvbRqT+JxGAYG/7ZQ/MLQEudmZGXc2YMKgditdYobS
sKtW1IHCEUCU+BX2VIRy9kX0SZfRxGmExwRjgaSQ16XA2scuKGvNXQEnly9w0GWaO7I5l12Cen+g
ZGDICqydy11gsA18NZf6cgPA4ciqgelmgnniJeR3Ct10ix6mN0bgbudLu/TbW0XHWYSqQnWK0biP
FSlmqGY0+KU9TKyWuIks38zrDBp3km17u/ND4Ztb+91gEko6xSKui5/GiQkyCXe1gbQ9sriQGsir
y2Oz+vSxNl5/d+jyQjKZwqoJd0dKiPmSt0KJFcWg9WuhB/BRPMc9kYIcatyL3gxoczaVa016O9HU
JNBjeRk1+RXKQwFLPeQXkzNezw1OudrqXqakM3lKbDRvuzqUp6dArdrXeth73QdPaDqYydryGbRB
NEJ+B38h3qZXKBZrbH0j9/sW4SMcqTG2XO7olO/f1PuzsnhggxQ2ZOj8gOV4JQwWh74Ze9e8N63r
OGgJisofc6xbYGD3wAAcH6QG0lRNlcxnk6YZq5N3IW87FlsqG8t32z6Nzz1Kb+yLdVNJT9XTGK4q
R7w6iF6Pe/BVhgou17mQUFUZjCWZFaR7VIubepETze+ciyvOJ+NkAyTkCWtYPvNazUxUH1y7Br+6
tyCYUcY5nYjxffzWoSMAFiBKxrT5avuvEiDNWhPT9D1LQlKU/pPdLj1+SqfoykbJ+kLfyfK1djbg
Zw8UVc2R/vJb/LOSubnheX53dY6Aq7g16IYivQcgvU5rl29Wdq5OlE5v6QBl7aIISGP+xtpJTBh+
HsPZlXfkyu5hFgd8W1D2lLlfBAFw5yLyHuURoTNshDk27NA5Yy8UvSsEftDolWWdAAW4I5AfJA3x
YmEIn0EmTQlG7tjDwaO45vsxtSvpaZ5oxKmPfXuh9hXOiWr7TeJ1tL6PT7V7ZLcWHZFRos9af6d3
2iCNqeY/ranpLULAsy6DtsOTvE+Yg4eM5L3nefHYE0cURvaQjoYHKtn/JFkUkx1q1tx3Cf5mDSEM
/vLJAIfgavsvfPbBwlMQvT7RT+RzO3cfJTe926N8OMJyqkaZpEhLUrLh7EUvN6QJBV7iGlBspG/Z
IEDoKTmZ2joBjqZCb1jZERb48CM5HyGdxgfY7j7+l+WvcHy2CalEEP1Bt/DfaPbl6mL6DRLawgQz
IPC+F0WSKS3hAH2Pad/jStWd32mrkX8bPBvD5roBdFCOz97zbqSDX/mwYEhgaymSuhzHq7H/UToA
w7r09Z1amQyBHEJYXtYQnzVo4ilofqY4m8LcIGZh9pUTheZreyfyZr/d9+V+FHvhhGhajVl6jsC/
DEf97W12A2BM/JXcrP9QlrAEhWiLlRn41rTUL5SGTUsHYS6MVx2wtBonzyHnl59ldHFdrkYeQCko
yzfHlPYulzlF3t6lxMPrfkAeIO8VrBHPlmyFCxTG8kuo8AY1ZWFGpJZvghmFtD/MdsnGhU+vErr5
MpJTWOmZfWUR5aq1dn+xyLor+su2IUsh6FAcfL3U4lVYmOp6ymhuTxV7A7dfj8m81YuDxvC6r8N6
ll6mpcqOpTZZAI+iz28vLBYwSchYfj5QhLJDfzV841idQaNlm/FGdtvJluogrEfBytvLnYKms8sY
RbIp/kjgVa75Kb1Cy8ZMYTFqfGnpGDOwi7iN6zROvHbuGhPXlpttePO8Aj+QWN+uI+iXjifaGuAr
WHBVqfrJ6Xt8xFZ9Ky0pVPR681XIIQpH5wLUzMjTrxa3Yvz1IZctb1Btvmr9IGyYVLWUQ2TAPtQ7
a/kvYAJgjxyFqX+pTfzbmZdPoCe7DtcTvFceEQbcWD7V49lOyBLKqqb2ADCg+Ae71uay+Fz9KH0K
zuFFuBlkCEQVUNx+kesTqhBXorK7Maw2TRNdFyn8/xOiUVT0lJihAha56BrgGC4e2o36o7BR5OPS
HM3C68piHkvTDCXPnEJH2TYDf3no95sjEaWCvy0dgRIrNjy7BTqo8J1PJn0bQz7MVtCHVpIQTDKz
BjLKl0Ap1OXmyRseY7l11IFPhBdFOl6bnYekq2Q1NMqkjrg6UpiQn7NyKjL824SrlsDKUNLFfPQP
+48sRB76W4Xly1twAMs01YY5CaAMXNQ0Ej53s855n5RLSJ6m6I6JrH7tufTj+ElIlJrTPrHB6Nmk
hdcICJxoKENTXLvwbPlJWM932HTCKRnn2ee7ibVa3U+El2nqx9CY6yIAa5tEGiJkbrAtC4yKbLzY
1CsGg8ppAPJzSohJmLIvzFYXAgxPXCmDtrDpAm5iQ9CFyKYFh8koYTV27eBaZ+cjyJxMoXBwKdW8
4PFlWFALyjewkPlzVSG5YHGrMEPanBrgiyhl2+04TB5x/aEfraleFwK6SX5yYGPtGC2P98Q8JOOL
BvwAe+WO42ssuo8e2rArNKMN9QXI0RYXd6OC1+x8lSX+/byDjKYxwbDr57/r7fboxCpbaYAD51AV
gdX9LyZU1tAsYDWmzKaKgTKzVcCvatM7Y2e254SmJmYlzAXlPktNQm7nDZ4V8EQ4qYNL8EjNNJgR
lcW46t8TJb3ZirdZWxuUkeHU/E5aTXCBEkGiBzPTjLxxml+eudmylnaEbVPBWMdNaZFVlwHLm3DF
RUhyUg/3w4G7LP7wja1MO/I3VRBfgDRu2MxGGAlBiMrxko2rBIy/LAl1FlgK4qeeJhTNg4yDQ4Tf
CpWO1/QxuMYk3PYjKTGvjTwWS85xCSRqzTnPyhw/etcqn+xGtE+3kjxtU1d+18yYovrNcUfGzSVF
5YwO9q925IKBpe132ax94qCy2Sbcl3mJPEt+XnTunW45Tt7jnKkN7vBg5cSjmzUWWxlmhjt7IFpS
LF8H+TaOV/OfJ2Qcg8GbwIOLSXQqXFna92Omn+KC66tBpQFCxPOLNOJEwLvU1XbcRoHGOcOhz+tQ
BD9iD9OoMFlp8bRABCzDM6ECDhYcpkunVauV1hWyNj6WMCYXf1fBPNBCyTRG6jlwfgroWUxNFGFM
N9vLiL1hSBt7Vtl2rOV/7/FIw3vbOdbEXDCcKerznxMfMMXzuWaADfRLJ8mLfBETe3hSjBho8mr3
T90gUCUwSV1lSrK4mAbbJmLrEVKhfRRqkX+fMMLeVQVlnxpTBzCZVbZOrhZ4gzGOHih8uqyFfVXq
gDZqvGwLt8/DSs4aW1eCk79MjbcoSBu38bcfaea2keMFnr70KIE77q6yApIeYmiYIg6J4LY0iX0s
4TUw0VSb7RTr7iHWauou004UPZ/VkkrIKnwQKPMu2kYrOHpa2VAlTItlHdJxSegyZ+a+ZwyE66Ty
3pw44M8owe7zr2GrLvWFjOt95RAsVeZOsE8zPwsFBH6BZ0igGEchWdDLO+4LdQtjEfIzCbmOj8sk
ixgAqHnNZEnJ1nu8VxHNzxF6ZHCJsMwlboU++8vDKzer4YD97lJfhtQzA3pY4fK06hminABqruHR
/S6bSuOcFpcKgDOirFDJeIO/QL1RKgaeB3rN6A96GqTCJZFmIgZaD1Nr9rgztoBRPjF5V+V0PBc6
5ipE36VdubVtiq3e5btdS+N6O9d3vpwN8qiul/XA9GkelxhoSXxv1Kkd5BGLZyevcNA6q1ZrU/23
zvMJeKViNQHBfRrq/J7nHkSj96cmwd3Cmhpfaf8YboEd7ZuPm0dEGtgYTYik3GIxW1uFDEiUZuE/
bS+Enpb0UUucWTHU2trK7gK+pClBgXIrcz9JrRydOQCzzWK26T/hJoXssPi6rqUsjg214odB3MyO
gzQEa5UJgNfI+HPNLIBrgXldUYLHUHCUaFLwECpfYbinNUf7wOug6iLTjSybkHQIIkt9jPlHnlXq
nX/OGoCVeAuA9FHD2Yy7NqBaMYwx54Kzlswl1zDaejsJF5JESDKZm6E+OWjv6wCyvuth4rg4QHbU
NWqCi4u/Vxzq/ralxH4TjfOmrOMROzLAcJmMU6AD2C7bc7fikGp7v2MyNeRnyMD84AQcyzGaNUUY
EsxNV3f/V5eJi60Q9Q/wufkqZhVf5+Z8QgpHyFv6JzAgVpFGXwzAfS5tfMBTgpHN0s3L+Maa0qVq
lUq20x0wyW/NJz+XjxWPf3LAgb59k/dEQ/VlPO6cstjurXSylw2C+fpM9+Nj47+VPA8IorAE1r0e
Expkt7lseWRx754tQCkJ/75LydeDiBioyi1NfTBXaBM2u3tGDq0SLwl6Khb2hqizUotdWRDgoWrv
060bVTbB1OBcMDAPQ8Kbgj8smI/DPBsgNgqjRd6NByGFRump4LDBxFAROw7KIMbKlWtBZI7gT52x
Ts7O+YsKssLMfKmknZF+8dcSAuhi9nlXq32UTJyxksg+YqxG67rF7n25r6GMRNb02LxdDgeVOh4G
ujTrZwNWymU2HetlOOn8djSkzWtTkmfzl/pa6Z2gL/MopJtyd9n4zZeV/xa+NmZlgXAqYYbL0lmV
FnvaWOHgkWlCaiipIzdwzLf++QDm2T2LaiIlvwy9rujPQN68xDdtyxpPRI2APPHmqK11Fe+CxvOf
MIA4OZtGEbMPliN2xSbdjBQDybKBCh5cQn2khJ+TUj7h1XfvGrU1shQ7hdXhO1WvFzEYGBQujSAW
7lsflnHDQxMJX0YXd9SxHHVU1F5RidZp2ms1ZDMRlaBHtQ1//6emr4sh9WoZ7MmHcAdkLlqW9mXE
5JrXFfw71riBjR6+biFil20GYD2MEtXQ0HIIKqVp5ZpnQKfSniaI3ig6/ajzG4wx4X1hHGJRy+UA
MgJ38j6l6/WJyTy+C+YtmUdjFGHB2cVnEkAjiVqkg4XhbzPVSYSlI5OEF8mj3iEr/mXVYqlMRJRL
Y1MjpKQs0mGwKAIJawiU44EXbPbRdakFTIDoGoksgsWHqbzzEiuk1pvDxj3SZYvXLw3KRAoPuXdg
EU+wWZf8AgbBqyJbCJnOt9LacLkJYdqU4fOTPq85kBc61kt5WZ4k1sOIflJkhLc5TBqiVHN2jbAd
WCFrri4oazlvszRMq7tktVD3wIXKNQH9goTCAvpM/3edtqLlYnUUrGeXCqJy51QOye/ssLyfvVr9
mMpa7KK/F9UNDkYZeUjhmhxOk++HISow8OVmO9oHrwC6i25OFYzjrQW8L74sB/i61r0WnU2YjTTW
/pfctv8FPbT9zlK6tn+kjORgh/XfS7r31Xb4gZryeSoSlEFJz+ny0Pf3gWaM8BNfA0oHXrzWCj27
p/gSWxpznBR6v5njwQNtBGfZXq3B+nVSFb+4xl9T1b4H8pLg0NMk79LCqrcLQ7Qtr43olZKhsEwn
8+nMlyUM7IDvCpZupgLxBinSZ/NfQMYZcJNpWmlf3J2aTR1pcRYNLfIKOGjOSB7AJ0Ny5QoqPNgt
OykZjqY67K6j1AgW98usiaJOQRbcvX2kwcj+XQUfKJVKhXlso55FymDVN5YCnJdFKxkR1GtYgPqA
ACfIFFMZBvIlf6pexLHvKaVTyNeo7E9tP6MFLldehgUsmCNHPBFrYEsO4Nc16bOIVyDa9ZTTR6rz
KilXQrW215fRYQR+Em4Ce5oMZwihyu3oozRImM0pbZILd0wiGAUiXDusuiH8cnH4/u/ikuSurX5p
QFbXdTSUJCMo8wV5zeZUhCxWJ5M7Ki6HpqUMGWkPflTtz72pAyK41qCeg4f9A/KxQYjvBejHbviH
tjRqwk2V3DJHT7ng+4QJ6TvXkOxuaLKC993RHNpMbUtRZ6q0XKNePwRSwinofqeG6zsG8zIASjpL
2qdXBQhJjhhDWZiWPoMSjPeGUkPfvkQpyWt+g82lpYbpdq9JmyottVk9deI8XhZFRzhyiRJdSXpU
C41FBVDKGXOf8J+o7dNbrbXtXTDlFMnc65GUsLlqVChnvkdZlrbTNUR0hJhi2Yqrzr9EVY5Yjgx/
UswtvVhy4O27VItPc6EM6oAf8vmJi1UazKEUR5Hghzrq0Xhti+TSWCbiY9yX1+Jy5d8sOw4yLS1X
EoezeOvBqe4BkX/wxs3xVOTyT2V8Hz+Mq4pyXMmA3qwiUs5VtoGAB6XK1uUcZ52NeRQEfaCCLsEZ
TZjZQWK3VdWzNYF7gQpuk4Rm1wkVOEH15rWOx0vhVj43rbNwZNvqsTaOJxc5DQRqrgk5A23Wf5LX
ydbHClXgtnJwrPB2l0BJLr/Sfd4cOeeQ0ES6lNA6scS7eYA8WF+yxBgQLYKICaJ2YoF6F+t1RFgF
Y/KUmkPV9TIv+cTRcDV6uT5L0hsTUWGyBd+Nlsr3KgBRpGGWNoCbNzHyKJYkUpanTceYZQrS9t+n
XyyXpgQ8zeqPUbb5qd6epIT+ShwAm+0QiufAqDDZTO4HWTFOWdGXxSdF6fNw2ZI5bmbNkXaoUoCz
SfPMVuL540gmOpq/u/85rTlheGoB+PrijdCUxyrWALTNl2qUgEh0kaRkIHX+Jlp8YocIyV7fh4Nw
rIRheO7pEYCHFiCSIKmDhMN0KCqMU/bW8SLuYfXi9xRpZ6Sy07q2W7wmCq54IPlzTAz6reFZs+37
AGNlH/xHVt8a4jXVtgWzPwoHHykxaUnFgbjKZWusI4pSK13mFY6CRQToeubiiT40kzmvCqR7zjHI
g+G1O0hpNh3M3NCJ9FQ1zxCrcojNhV0XSer5I2kWUEDGZKnigRlIqiI6YTfHxl2L8tpCrqx7v/c/
R3LSHo8dTIj4aS/EyAYSfOoYAGI8WLXWVWW8yh/lW2yRxo/a37t+585Qu+cx/eMio/wpvx9yNm7U
In4NCIc7zlvXRWT3i8FDFjaXNc9p17AzI6tmdl8RghuKwSay1E+/DAw3xwQnRZksCUbu5+SKoiY5
wEf1IBfulZC5E4qCd77WLpwTW6D8N2HWUNPI4Yzh9na8SiWQic/dKgREekt8mujOtVIbKPDSwojQ
6eKurMUCQslLAKwJ2nHFVvfxfVlK8zzaos6ZAUg1KjQVAclk6KtngeroVjLmW2pEJXmpppz01y19
imdP5xhEiRe4DLXyO0jwlBqIfLLq/qBuMgMhL0wObbGTSUnpB3wCfTacav+DZvQnDqHu+JMpDHRz
E6vT+8Kb9FndIu/BdZ3ZZ55Oc/J4A7HrKzO5+dDlOxF+7KdpD54Y8W/r7/fKdDbpxH/TtOkuxy5f
EhVqQXisdS9NL/SuOinmobA5rbVa2WvcHYCAEmm57SwYzTbV5EFmvw8TZgPNVBi8i5Zi2JjHkgX4
hI7MVPfDT5wvmT5SvuyBtlVVxQJYMvOmVmLHy3CSmukPRY1rso1RdZjS7gFSOzKBS7UVTxOjNvE3
Bvoq1r7gf9FVQexqKcubPLA53arvADJ6f9ueVeSUQmyVO2gXn60yBnwdm+ftiwcHdo13gAdGVFw5
IUbKNYh7g9FzZmStfBSfjYHoYl+SeB8akAu064bOWEzThU2VsTAgUjP/dweHM7LC8IQjmCwYZqrL
hIdjbuV8xo+aPRIWOPo5DEngMoWOOYKiRp1pkS2DxDddWrsoIrcZmEgfv6IBH91GPEXtdcenFE+r
mUMLVmGGc+ibAuz7PsI62RZFcYkEcrMxuT/R8a6kpIIMtTjBGVt9kttfvuj6unWeHkLOP++OZNu+
qpEeHS17CW/+CxbO97tK2S7uQ4yKXb677zuaCY7EhYO/wpai5pUzm6RTXVZCmKQ7GbE9UG7vkCeY
rZxPj/TXYHA+cNacK3QkyN1B6/mKmAQFiULzU1jTuUskRZjgXbDANZLOIpV6iGdD/x8VLmVEuwm2
GKd44Hsi+joiyEH540x8efcgAZPhINZuh97wtJZ4YHOgubu2JSnwkFVZDCDYSW2OoCb49LqwcN55
AcwIpGvt77QCYJspmuYphbQxPIu0bxHpuwXbW4/8QoGIMoF5t1wwpp4E+WUwAyyfNtHRmUjwH2lv
uvDMwY3x8JAIA6fWgaOe/w5/TnFVo0o+4PKl8Fort5Jted3Ev2SCjumTNNwnd2OuxrvoMqA/dUzM
dNxiKwCqbs5HLkfu+vOUSS1mtciTSgjJYNuN7IIc79MeAHIspdNbBXddjkEM3FJixK48/z5Qpds5
FDFAYnJ/FmC3zXzTCnGiz1OrgLW+peu0ubIymEzLZmZCnq0paDttAR70v666kiyS7eigxXiwSoAH
L52zKbVbZ+mEXo2LtHtqZupu2X+bfhsU8dRa4TBTB6LLyhN159zvFhu2xc9WKp8vbL+84g+L+3fl
QKEMJX9Mdo68hSJHFzUZn+2bakJgxju424a9uJclchZbeLUpqDURSSRuQhKatREhsoiz8CRhZGfx
qG7ssMfTfMnm3IJ2LobmBWTnpBj/61pFlIkToQZV1jJ1DD4kCen9fltMLKyejXsrERrZksNVFF5x
e7dI7o+pPsDQBStCuoOkvdDWSi7+jyb2mhQE8HYcbUo6CRlVktaB/VgKYu3IJTJpOYnrM/EGesvR
sD9izwcv+AlHQiiFzxDTPCaGtak88xanoxVPVWK00O7UlSva5OesRRKcUeszI5IGqX/LMzrvrcJq
jpzcsnYWz3WO4XMwokg0dFBVlhRUI03rhP+F2+whs08danNOpHaKVMRVSure0dukCT9BGPp5f5WN
Gh6B08pj0k5B6xYv0YgtPGcTTgA55s/iLCXjIoW5TEUU6t13Y92eGfHRIb5H1ot6AXnj6fBR05Sm
Cmy2QO5W4uzcuZ4mmLm9FAEVoFGw73Jm8rgp58xe093ryfLQktNy3BeHso5uWgqFndj5qgLEEzZ1
EFRA+0KuxBpSZEjOIrr+2Nt4U/JNBTyMQs8CYsAnlIksTYQ5xAgh+ccdeJ8iNKRW86yA5dFHXy2F
wTmK0YBceli5t7xxxrAKRnEiA5DP/oj6BbrvCG88mED1dJ8FlXEDsZ4ajcxv1k1a/zv3o/yuJbhd
g8uuhf6biKk8d8NfrgZrLyad0xXooOlk6cvILLQpYcCrM6yByjtop2kckBSS/ILecUBpweWB/Bng
OQmPrhXxJolz30wRb1dpwiNCj2CkZqp9j4T4svOXZmSs8BXLBdOHcnb1kE2sZT191q4PkWNP5Upj
9x1HuyEGrI6cOJmkBoB2/UxWjrzkZIRd/aHHOYoqnMTQX/eCnGxU2LniDXdIzE763pLYDBTE0oRa
E6XcUHd8BDbE+Deio9I0CSr1m3gclA0ePvMauNxJM/zlnVPKP9/pqmSPM+xHYgXknP5X02yodDoi
TcbcqJpQQP8VZ31scxc1CSEe3G7iQrpHf8zFseGY2dQAuvMT7mdR4uAvatTTWZzmcQvBqh2VRKqX
HQC2Jr4e4PzaEdKDF2jaWojB/Yh+V/oBHkU+yfoSs++isuHs6Ui5tb9V6V02Oc+fQ9zN8Zm+8Qgc
vSq5ImLuN4SD7IKBslkTKwoGwNkpKjDOjOrcsDVI1Zftx8Pr1VbK7tXK8aOp/sC56Bc9N9CqWKJ5
ib8e7VY1YrgccAu3BFGHsgs64W75wIoRPEP+MYYBgtW+vqKia4jh1tUlU6PBS9ZZV8eczHRG8l67
YY3Ph1fcuI5s28+gjqxKEKQFo8XChkXGQtbpXjA2AjfPYVlw4oSxKYM5g375gvJqLGuFtU4yoa/u
KLQWav6kS+cn94En5PyCSHlmicXHbDIHlWjZMsy1TnWtnEX6/UYy3ATaTEQcrkf0yNj0LQpeRQ0H
H0YTZqiMkaBw8Vhkvpm37TjJ5o35bR7CmoIfBiRON2gEWpz6qDyy+67BEJbF29Zvj2aIqlyLiwkZ
Jje5SKFita8nQX+PsZiVK+GK9hHqegt29kvvxa5rEmmECfbRao8bh2xJCjm6IkJ/DynY83dX+9D9
j87D/zTIPywxKPTISUWYDS4clvixGHG2oIkjAtXNn1gvh7VloLYXDkDiCI5kTA4DyxkI3xiWKLw0
JUx4ovz5cv4btcVfg+qk2/9ahSuAlW37ys7nT98CmyciCnJhmlmK734J5tW8CDIGzVru0pQ6jhJ5
g4dDr4tapL6W+bGKLcO/ok51OUY23gPHbB0AN6kJdexcIe6w01OhIwO4Ti0MEEABT2XAEUx3bl8h
fHTRFu6SHmo7czVUFEj55xR197bNpMItHv0rUlU8dUSJqAGa1hXuHBZKxm3oXwYvDUEfGrT1Pnqb
AaPLAH3ktvEC8ZV/q/PmCtkwfYuliaQ+8WZ5RwwgAKWNo48mWh5nOw6Y3YWESUYP/yN7eWAL3VXk
k93tdLtwi7w3RukiTOEa3Bkb5l4aYRJ9de/ViuftGjpUkAeoSTQTD2q2Elfw4VuJIN6PhvPEghI3
Y1flCoEjmIla1b7Ew2U+cEQyC2BJvtzX0xE9RQuD9n68RYE7hkmdHF3/X5rCUFFtuj5e5U/q44D8
UqrQNG1XiGAjML9msnLbU7HyHxjPnhFZPmLLnSGoFXZ7S59bI/8wwW4QiiRGNIYRN6rgoFx6ax7V
ajleYI90uWfLn9NspJg42zm+wRZn8DE8z0xKz4XidpfWNtcRQApS0EV5pVlLrp2k1nacag25J56W
ZCm+eZE62/sLgzJqMuohagadOS/tcoibREpfpE/zVJKWNKzedGN4MTnZxKLwMftoYbrdD5V/PiJ/
yPmaQ0xLp0qZlwrEdZb85ujvy2Xwki5fbPqsommUi0eoH2Ou4ghvzsDRoY9YtAZnLxf4HnIfoJwE
r364nPI1ELpGR265p/0NRkau1esFV4NT4jhg97UpSfsstOSBLH7x/iUHvW70tnEtIBIcbOO46l/5
uA9p28xRf1khi/zwDCnf3oSr3m0C/YikN+tDNQIKoP+iqj/ww9ptpGbC4BRHWDl4lofJ67s/MXJP
r7xpNJoSw+W10LdvcsyVh62dXgCqdpR5aT1p+10+sFVJSxq9CFcDiY+fkp+sDPM2xU8Gdh+rFLr8
s2fkygD3+Wd1Sdj9UonK+WDYzjT0o+2uoBtxEd18JM4J7LKoXtE0DT+VpjdYn7YMs6akbR/wGhv9
D0hIkKAeK6Qiw6VlEU0NTQx55rrIk+3GMYG0ZI9J6rTz75gNkDnI1MP/2uut9sBGZo2VKPn+iOQo
mnWMprGXqjdfO26VP3LQYduEimpzrZO2jW8JOMasXdtCiuHNQq9LIluzWYP2fzLAtvb8aV668CXP
pLCRmQ8J46RhCu4L1Hn/I3+WuVKxg5L6SZprF+CzqX6d1p1jHFYew5q7eTQ//yj8CbAQW28Q9ZZy
AoWo95hMIup3z6QdGNXoIRgAV/jDHM6J8uanqG0ThHV2WjT+pLaG9dRHw/WWRrJDDiSUdl5Jm8VB
UA9VjzIsN3UiY6iOxNlgBaj9NukMeEOj1E5JeTDBkkAK2siNXSAB5dvi8+cqE37KLOvlLXy/IfJ1
1bbdSIr5hGjuCz2wQaB0PY4YJjCkPilX1xxbgeM6ANsf4KUeuspVGEbkMPFmhJ38zpxnB/AROCPm
WiFfBVQYwb+G99178aEHveSlwBFmxyXy8uDsB/Q7YCPnF9M6idRXiEJFpbWmbpXpVZzI3epmzPHH
p9ycP4qCigHNC4pgWuUslaBM6ioUKMN/gjx6bhU/1nUpj2uxL8EqUUeszPz+Vvfd/Qmoecjs88lD
tmPyOFt956DGHgwJYMEQKvbtf7wHruLrT8nusla0dgfD2WNEpOIOSes7VW41nkNfPugqSBkRpye6
FogOBknCwcfqYAhB5F9fEMHiqnQkgVCaKeHc9ERAodWmnvhjx5NsAiK5zsnPPHmelZtjHeDhsH8y
rFaUiPLNKFeRXLFxGasHBZyKe3j1RQLf8NK1i85Ch3GIqIu1O8fE1tYM+RdUKaYzMH6XytZ6QPK9
Mc8OS1cWtVE1TrSOljaOp5dO0+M1GhbxPi9z3ySGLbGM3H71B2mZeM+DGN0AEJIrheSDwd8MJ5bk
2vgpUTKTSWNDcHgvlhWlFWcXp8UPbyMwuzOhjVfCFKupMjgqcoAL5kz1nf2qDOAzyMSINIPc2klv
YN+Mo+/h/mC13dopNkg1WOmoFT8tNUhjtxie6DYAGcT1xLWy0kzsIN12c/d7ts8Ucm6omOI2fLcu
ePP3KCgVCcM7sUBu4yvnzsNNtrOW1Up2GAhEuJmGyNZOolonJntwVFlRDjDNxTUCNEHctyEfcygW
lGjbeJGnEX9qZ7raa+4WDIZ7Viw7jNQsuN8TbNsITdeZEtTNwm1AXZQQNRMa7MyxART5YcxM7Nxb
2YGzMoGaAxN3Rtp6vWC73SpFboTyYQ7kvygITN4nSK8Uxa+Y4epW8OT8NX3GX0Y/ZL77wGggCwEV
1HsIgbNomeUOWvvRhaMMPB49yGbXNPGFQQV3SUNCkA/tmGZ86YwqvVG5/w79ZHDYB01VB5ZOT6zm
EOK751TAkaskpI+tGOH0UNGoV+dbGfBsOqtZHz1E/Xwwtt7uNWkXX4/UqnjeJtiGAoWDxgdT1RKr
B91+wLbgugbFckmsL3+IEZfrm/+LXhNBlhmwUyQqRWN1zQvSp/4hrGP/Eo7t+732v4Z5KAEn9TUd
2PrpDk+1FoOcScPAlcFEvXcgW5EpyKMlecL97AGundWN4HIE2Scn48NdhloLJY3My9EXVdiBjkXi
2sZRFcoSUXCcEOcGlAGeb0/rsdHJ9AGwT9lgZcZD7AaYG+/E4fMYb2+G4871jdEQaafTdkKMpPgS
MP4zgZx/TnD0tl/eN8VNhb36CLk0bDPkVLHU/cWdJs2EO9kmxtm4Mlc7xpcsb31TEIQ5sqreWZ6p
VkN071yz4SObrv7W5bNALfEeCKWjuC0CWJTBayqprbbFP8x38g7KZ4Zg4FUeRMlnErswXYYYykUw
eDmADY8QiI88lU6wjdDZzAGWVDvpGrzmYSIdqyDMQWAvdSf2GbcMyLitKa1kJUmQvUhYYO7vVL2Q
wjX9iVZ6qG4u0tGwNPGzCNY4GP3i1kmr8SPDSODriY5ETq04xu5xE+ChSLe1NISzvWxtUllH7wlx
GB8bcJFdYnCekjA8W99Rx6Wb8y22o/b6zcGHNJ/zWs1wbrAnrSE/vLbVevJo4WXAeJcHz818lh24
qiQFUIuq8WT/V4pthqGq7GR06AgcIkM7S6KxgrfQCWfz6VkoFQ6WMR3l+Vfi+lnVSK8YFl6DOmsA
o9snE1bWvSiYlFDgxTeqAKuiI3eb8yYlUL5vMTe74dZpjt0LYa5ggo3cittR/de2VyvogA+kq5Wu
yUgSxkCOuwtLzG3YVmHuFSu0m/C6/Yp5RAO2JbAwA/D9TRPWpObtGMChxvlN5cqQER7hE52yUAFN
7tAfaK9khB06Qc8lMQDkdsK/LwKLuKIJlopSAn+/R7xc+VJBbo0+tJidzoI7qArfsSB6EPO/kDeJ
4OIz7Sg5aqTsMewjLBg6BBwJIus9PztGUVHR9OpeHplTPfUYxLc+0smUCrHfOi/9/Yo318ln4uEL
cpXrZAs0j64EY0G8jkVv9tvMWbX2a5PWsKFIFltMEM5oEblfFN23lWuQ2F9rYBXXl7DZ7Cv5UwKh
A5kmPwiSzJ6jP/ACtGfhzFlfkwVLhlDEbMibNZfVIX5h4AuwNQOvtiNfgJIn8b8F36OJl4mRIwmX
O2hhF8It3bc69wc3fsg5CjulQMEqh8+0W2rl5jJiBePC8e5/AdDrHZ4NKtsW0y6uGCRdqMRGF601
09F74GLo2+OFSmD/QFYI5tcdLO/RFz7FGjAOCMWSPnmUmQW9RaMbvSTGOqFAVN2/jtotUt5t9cLz
Ory+RrH7HMHYH9GaxaaRM0Ek7qEMG/+xfEfJCLpBInnevxkJt6/jNPDfLH+aKdgaqeb0owo/B0y3
LtDSE9OusEDuC8UFMKg+stuXLsZmomIkAN1L6eMRvll8JRTRQJGgReZ3MqzgruV2t9uzKAWhiw5K
btHQb1moxoDGONdzH6NFyJKHXlrITFKucaggwTHynCVQhomnsHVlbGl48geHtJB/5FmgWwJI79nL
6xY1Bah2IHvxwrXa/j8ccwHGfcwd+KjT+vZmveIkogy3l0g9rbLviTzuyaCpWCW9K3jfa9rno3WA
RU8Im1Xkndd6gtM7BDTE+RUjdgg5xhOfp9KQ0IP6hi+LsKB0mNXAySZsMDr9NGb31hRoJwHvd0PT
B2uJAZ1aU1h4E/2BFb1rSo8arcuWjaidvs6bgM6ePf8J2ykVwpfGbxJzuuRRcTDCyL0vc94SfeeH
QG8rH2T2Ngojki3QwJG23ZBUup84Nxs8Mt99SYlNeL8TACAt2JfKHeOThCIgpmuDIu8fXkvqrtsY
vv5+L0sJQMAOu5DJzdYVHIVWwGP/ETjtjKeJkwFAIB+6iJ00m1kwLa5B5NidQhjFPCGdFowyevQo
Gp3ZZ27bxgSa4sxhqtIcI+tBVG6NHQ83VD4T5XsfCcxqS5xoq4EmVe7rTbAvvz+wfIuMTXT373C3
UjSj7tV7t8XdU58RNjGYC1mafwoL15SUKHUBKqp82ogFrplYiZN8nObFdDiAHKiP6cK9CXYQT8bg
SwDFSbYsMoU3gxg7Chik+kwMW+jngou8EugLSoshY+1eOJVUtWnKZaMcqA2hTN3yxifzlhaqpwFr
pVLGvoHkVlUvQdhOuFuiIZiAXfXI2xDM/fgVHAl2EM+hAcn3vggXgbXcWJPIAQwp7dnFc7sETsvZ
4FGtuFdJE9fRc2kXaHaCDkOrDU6mE5o+Cj5nc77nEMv1zm9pujlgzCsThb/CWpv+Ls/Woq+l35K4
dTsEzjJZUHeVwgkfqIEDkWjvYRDisxfx3T6VaJtrJSB5OHUQtQiIX+ds7Wb9c8bHpZk4ojwUXiIk
4lvLjBIFZaYQmjfb3t5fIlsLO0tpBByleBCddiBbQok1BQC+Qu5B4bNjkBdObzTOqjLCgVEQuY03
gzYrNnWwyRuSh/y9s+69E/1p6hTIKWA+OzeJ0KIQAdbKBfkJPmhYnYW4MtKCywuPeB0E3h7NYOM1
Csr3a1mPkQAwfmT/J7e0CnbJCiQE6CdUn5rRCW2mX5qY3ryWH1CB3R3mXamRYyNhbE8L/m5VtsIS
i0WYwXJ5K/W98jfJoBtqEwrzZ7G13vUTqZavk1M9yOhfYn+M2HOB719+c8icjxgN86T2G1pZ8GsG
RpmX/dnIBVFJKb1icfx7ONwwyKDwmpTiuBCDKE53q8R/jaUnNCWtyGmSKRu7Qhl5NoGDPzCeurln
mB3tJbQcwOUQBXMhfontYLgYlC0rIMgCFAD/zBIO7cz+S7kB9flO5CyLaa1DtbWp0TJz2lVa82zA
ax4eD4LsjZ4VDMF3k/p4fPx8xK1UOJyUuv4t6jnkbpBl5088baZezy6tot5p5g4h+iqIEeDMAbGw
qTsE5gDuwPopkfgNANVwTnlh4cOwtWfaV6MaxDMZJdQIHVOQFNlrlsr7qfhNGmu/OWavc2JsIeEQ
wSvAjnke/5Ji/KOq3qIw7T3KXEHRgN4/Jbzs8IsVXx8cNFaS7P7dt5bt8IlwbqAk5R7JU879hEDY
1jzenjwQe6qIDfKI/c/5ShKSfYCwxNIaZPJyFGmPNvfeMVsQUxxCMNtex6sUMXjbRppwIOgXCZ6Z
IixMOvILqrL/0RGesuFL15qgRpHaBIM3xb3gV9XKn9hc6L5fDCbpBT4ZDaT2irEi8bjAHqwrGD5J
aiPvqn0snJS4qa2eficNBJcYnYHmK7Q8y0y5OPyg1+zqIP8nmfgA8uWPmnekY2XqfuyAzIILyOvi
ewJ240UhLTUA1lZnAKXt/FiHZeXZfl5qqNDUW8AmrkhzSSMKNJvp5uLf79Pr1nmW8UYFQeMSaFRP
xcPASSNN3jDAoXlpvblYHht+UyT0CFxNUyhwjw6JMKGcwz/YYS/IIV2citjSk+GYpqLQmKBqXufz
5GO6BPW21h+EmHh+bak1zikg0CT4Lb8155FZ0zQNiW1Pi7qT2EYN5AM35MN0RsnMQc775CIo/6/d
b49nTgjfRBpgv/WkZG3m+WOY7j++4wvZIjz14X7gngpDO/ivemvu5HOFccGeszhqqjZ4Os22IVlq
+TLq1WmdDQizPPbdMvObNgAUlOMsU3ZG28YMpvf1iC5Vu3nEbjsYL6h3s7R5uTbX6r3h5waSbgEw
h7k2WYIIw8MeM+V3yBCfyHP7mDc++2v1aP60CaXISumvqAJ9ngVfu+Z7ae85qpYx4a5wG50xuYsw
MTOKbIdFAHSCCZ4YekeZi1OOaK3oM19r6YrmumJZ4MpEpm1rXsA/7anhgscIZQ3C68oMG/yZ157+
/l7VP1nVXl+VW3nBBczUD0Mcyrb55fjfcb/R3gfuLt40AoOmDcJ4iSo297/Wohs07lnPLtbvNRor
N+ocIRXbOCBf3eZ8WrR6chX9o0II96RIflkGyG69fPd9mBFWLpPD2j4JxHY24T7oVhIUG2pQDqjw
PbGAmpC1jklXm9jydJ+K1hwnEt3cig2/4KMULJ8q8mCrSFz8o58VUR03LxJ98tEYAWp1UYhsS2sE
Z4d+FmXkAYnL+MvXhOY0dpsHiO0RuYIWrf4SLSMFyl8CunxXkoFX/NGZv6VogiTqmALd2UKUrMb1
fHgEmUafpRk8JkrVRr//hx/bjaWerHdq2L9hZr5bIceiI21+qIJ/SuMSMAUSLbtPH6tuzCKKeIL7
uXx+gdJluE3Nv2C6L9yrhD9+cn8iTGygUXB5D5PGQ7CwF2FkIzlsM3xooS0UufeZvljNh8eT73u3
qgpf4gTqjzige7LJgMVvBXL51CdSOyEZTsuafvbseF18SXe3GmcSVgy/81dJdarBT+ovNTEM4DBG
pp9vYjU1Fnal3mcXxiFsgGlzrkaSrIN+9uc+zfIKmZWk2BDQNXYXcsRf808X88nK96i5l8SUoYfL
sznCdUdukxZkm0Azhg1cUa4GntqxLRRuvlNFi8am0kMlNmqCZ3zAPXJbM/PimzC1YQby/JFm3Lii
HZWJ02IoxDI/xgJBffFgwoyFKMX26hx8u6QMN1540meWVwRiIqcO6X3UlbgpPb/QpeChLf6Rm3DQ
M7SY/vgrLqYYG445FnKKWi5mIEAYtrqFoxmtj0FHAFLyLY8ZqP/jF+kjCNZAYFz6SrC1SGCgzzkE
xgInonwL7igyQrsOYi/JBct/Y27nlhgR1i2tHVIm5007GmserVc1JeSOlrSVW3DVpiBXb6LP051v
NUr/2vgnRCzVN/ajOwZ0dffOd2Dsgvl0yd74Wo1QIsYayW4QjRobtSChaxYBBx94uknQxtIF+dAs
5lMtlMdScwVJI9erdmLbD3ks4Xj6ST2BthUgfHGUNtm6+f75QnPgQpHKu5laVVA1kYRlpH+eKyGo
I8HBEJPS4wNQDvCgjPaB10D0hmx7+yOzE2xQQDILzePE3vsy3w/jxk3YK+atz1Nwz6cdUbRj6T7c
yhYMltbtZP/syywDwBu2ecKWkxSD6SPeWKnd1P7KeY007KG1k5wVBvPLrD+iTb/SLB68V5JE0RPJ
KqQrM9lGD/tsQx52urq9VYLlKkspzTH7ANhsEHbqDH1TWKLqBQIHxSW69u7oRR2C1ya0KVlbw/xS
dxN18F7tnj8zY93I49ZEvUP5iFvuP/WqUE4PGDyZ0Lq8b3r4ZsHbOYif86HGhdxXCpbmWzowfmak
DAFeyRxP/OVBTZp6PH1MeBb7DMas8EO3geggMRAd6pqY5v7BTnhM7ccnjejHrcrNchPlTXTIeCdL
RlGONMlGFFagzk82ulkSXyfoFUdp5yA9FF0ldrgKaEmfHbbQs4z1sC7d2Y9rcEyl0+SdanpZ6APR
Zgp5Smg7ig4aT/++FCMZANO9e3RoQhiB+ebCRih5t+8Z74oLaZLk67A5gE7TB5cshn6hhFxcZSyB
a+Psb2dFMKGF398dKfmIjc7t9xslxcSCsUer0i2nMshzpK0HPDLvQR+eU6+WBBHkrHVvfU0P1BM/
LzsHVWlAoTrTPIPT4bQJnZBKE3IdMnxiYiEu8u8cgaqtujVXFKylvm6Jz5otTqD2XXw99ch5an7P
p4B07gBXuWKKSZXtlZyZIFHE5f4Pmedg5gjQy+Smk3XlGs2IkPJ6HgmKEaUXzWHBJQZALEW8eDP9
viGdvgVFtjJOyP1l+C5utjQklSQixP83uPu9S+OgVrCwcIQGbVYT/KQP0UjiAHyw26tL6Eg7zcWF
UBve07d/znWOAy72v0MG408mABR9cSdvGQSmV18Pv7oDvvngyFptgNFiiVUyN3Tn6CD6nxWuY0lI
/fbK1tc2nlI6s9LNBWV/07LUbj7yU61yEw1iVNheOi6S7P8b1L3fR0FEYoHeY1J2ImiyqC4Zg8z8
kTyoMXIeKGVRwP7NGVWl4AvEYk7pFS/CI1JT5e14xu8acTzfDulsNqRwKq3VAQWfQySreGzQdGsW
vtDMhFzY9LOp7YsoWuoZrgO1CLezoGkQOzpLw1sZmYhSoXovHfI1i75OrlhZNkfj3+cJu8vUr6gL
t2o/MBL/AXzIlBTOkdA1/uBzsgBgNKKwWTrCjP8q4wg/EJ2nRL1CyfKOTfvTKhMr6PV2ByCbI0mx
NymlLIcx17mjTFxU1OtGGduQCHiaZGWTxjfBVVhNlivw8cEfIT+YL7RHYPdAuONAngx07mGbejvC
E/ouwh6Uw+f2fFgJ3fr/KJLY/9d1dn8N1nEh7BjfDyyUb+4PQdiyJ7Md4T1Hz+fAXdGQSplgsyn+
hZtepaaCSJz5b79baIfKsdGBgz3bEfSpWqyD8X5mMJqS+t/BICRPkyXSvQkxGix7B5RqjWmc3nFA
+ECmBZgscqwrsAGxdCW9QWlVFXusz+JSzVnt30Z8W0NL8CSiIbRGgOHc3alm45MDxgENEGfUqX4O
wq/Cx6NT5Nl2Y7oG5cGp9lZcBp56TA4HXFitavakaPZC+LuhlRppToiF9+kFq7y29Tq3rb+rdU3/
5Tbd9a5EqRVBhsoA1d8MHf3ikWautnGLlZPXeLQeGl9d7B7r8I6A4bfbXl8TWYcp1cpF2+toMOfH
s6rGJvLtblrpniyf+/VKa+GEe06/R9OxbOhKQXBZ4wQTzAOWo6edQh0A731GIP1W/IgOOJE8OnJL
YLmsRdMMvBIvvzH0PjIbu6GHUK3t/xO6EYOmHFF7wYThkAVSxQ2zFlpTtXykrrYCYZNvjL0pjcEI
ruuNLGshCn4pH7ZjmbtWKFNT3u5p1MyWziHCAfLlnGfAklnry03ipsNPlwS/csjQM3XxyZJVP2r8
SV2vGA0+w0TpE4twYCD8OFCCS9eoKgjUhBUkV9seL0XA+oNqHSvP8MhFg04cIftJQjt1f/pd1ciA
r9k1wKAWUMT9u3DA0A1zBkgj4aWLSnR+eCboyVw2V9qk7AZe2Y/yqm0byrJzie9JBv16WmJBBC+f
m5aZ8r8pyd6VRU5c0QSaAHq3TZCMtQ8zOmYwbmHmWD4aAtp/x+8shK7l6cAnZNx3lg9LxuCxzCYY
u0CdX+8S1zBa4q4sS7RrPOuOXPVs1IogK5AT2fnWXMJ9beKHC8sGBIBkBgtAas2nsTQyDQraiPMi
u0O4hv9jb4uIX89ruI7lL7rJlsq4/TFK0M7YJnmX2YiH6vygOyipWKZVc4fTGAfkqJ8/s41r6A4j
g2eQtC51ImCRArEN5G1nvzbQE/dMlZPiIIudjj6CSDonVFZXamuZj1f1LK0oqLjraDJnFfY3uZ3h
jNfQTMJWXE3nXkXkc+looswrKq5DdaPwmTh24Nnk7sql9sdc6M1ogt8JicmvF4PXBpkpiBn4sruQ
c8EycAMTQoQng55Aju3kaA4RJ/nzIwp7sHMU5fSX3l8+1zBzW7L4fyA8IUBCTQlVWaYKn5p4DQmN
ARvLiDyajyGRcpmUIpysEErNNv7TbkGxxw8usVfcv+UVmBuHk3EgTeI9zbadnRRHgrjQHB5/cngC
dzpZNYvs0v7lGfStDrnxmW23YHQ7PHD07K+REHBGmtaE6STxg5sjm0M9OioYn0m4tMk9+Y3Mx+z1
+h0pZrn7PEKeE/VdU/pc9UVgRhumg7ihNccNQWfXSQpH/ALO8qZ0zNPBKHg3IwZfF2oSx53wSU9w
8vA+HnV4V6XgeP4U0l7B69RZxx09xEgvwtb1PPCHDE41oL4VCdmBlK1rjMOLsHu41ZJeZD9UCQNQ
/UKfkm86a7jtl5Iy+kZtIP4Dc/LPkJVJi2TsYlZbj9d9f6N0mGbjzfziOH0ZKNom2HC5g6rg372Q
XMdVs9RmMWwUu4nW4z/EnXXqTOZLkZ7+N5bK7JevzvD4NdEKUREy6RbycsJI97vSqUy6WRsfboZD
gTAT6sZUTGx+hA+eGqpJdvL2yMxJByToHtEyxbU/bGinn8FBIJt0aRmbEO0DUTSUq5k2Q5GwmwPi
B80imvpq8MgAYMyeqDhUzdIngsQAQphKst4YUteQEvNez3RrpCBttPPDjCwpaYvwpEwQzaGmYzjJ
TXQez12uRZmYcty0Ot14ZvU7X0V2K1gTwJ2SFtPQd7+seCAQJEY1ljMga1IbXuB7j8U4fFeoTgE7
+2Dxfa42smBbZxI9jJvQBpeNE+KwqOI74VMpcSAAMy9t8jAFX5aC8MydGEia8xVwm41NvaS/T1ZK
XCcpb8dn5sDlUnQXSJiQdRhYEzw/1cER/2TLewOamhq8l+Dhp1qx7UEDeY5E4mo2O14+J+Zy2Cm0
C+uPaE/un9qXTOPCiMR5MVW4i5zwm4xAR3NaCFyMsu3oPgKWJDDCYmqOnzID1qLRiYL0jJJ1eOWJ
YSEvhc+zdXKrYa3kXv8cGWQ4xSf3UttIsyZgEcr+/NVic7gdxDvdESrbhcvGPsAJpWNLbX9rWEwO
HUQcMVrU4i4wi2AeupFFNErNdfarvXsdAWbnBvFqh6gYuKkFp5GMFpQMZULSDrmmOf5TEJXCUjIF
ge0x5c0ufGfEXh0xPpim3oddOzNR5B+9SLQqPsOR0KbrNzKXY6iZIH52w1agG1oQFxBT0qiDBmNf
ihKSyKiUbT3VWUrBdUfLAGEIiq6aIFFzC0A7ckHKmUX8KIDUMcwL81BZDMdFILdeqyCxoAy7jjpP
4gip4tp7Qopiq8epUBI5DUxL65HyR6uOQTxf3rvetF0BfrFMp9KbY4SOXPIFcsgMfrAW6+buEIkP
+1snBofokEFMTH2AErKkcu2LWHI9qTPr2AsIWY9BRfb26FQtF4Jf3LuNCMyEjQEipHG4bYweZLkT
hJPDDYiCNpqPYNkNVYvnANilFtEqG0iiExlTp2kkq6hMOiiu6eRTTZ3xq+HQ/FELYvUK6n2bcMh2
HTrBbOHceA7abcg4hhgb+SAl644oztD0gAbYxhyGGQLfDbg8WtP8ICYIJ4Wcnfgp76bg68Fd7QGS
Y0G8zc6SY7B5wZMQzv9iSdq5mJ85i5JhIsdgzoTYJ3mz3V8M9/Ef/6qXOVWJ6L0DJQoST/usi5zV
1F3nwVWaIvFxnchbD0cau1dhG6aj/ISYE15xsl3GHlKwIFk7BHw84KjbwfyT5+6Bw34zrGgZuMJw
K5dl4iu9LFtzt5gQVZN5jiRY9omxabI6l0FNKgShrUA+plcJ3/Stz9Tm7XMcsDjUTbC5Ib9RM/dX
Q9pV94JPvgvCBkPdUco9rqOk2qACptBF1+CkYrNcmZ0Ng1gTurpDbgbqrDBX6LyB/7hFteUNvHLd
V1EelgM55XKBnQkyLAilZmnVUnChlb2cp/nXdsq5kY4TIfMzP3gAhfQcYGZjQw+A2H6BBiWyZZbw
JhG17M9wrVxtaZCbSvWtguTDN5vDwtMSRGJgouK0mIRHdSj90tV3WQR7/5RXGyW7hhNO+4+HVLmM
ShMH28AO55KFsQu+6dTp5jphY/Welmd0nB2EGg2cAjQVTNChuYsgklOrDS/tAPIJQIfmAlrIPQzE
YRQA6cvKhNQpBvtH6VKlq2pyFjmDpOQX5QDeANtOhpnz5RsdP1fWBBRcdETXLQD0/UYwYS9OxQNo
jktWW0wzaKyCwgI4YKO7UcZUi2xz92QMjHusba4Q4xm9PpUvEQZkpO5IrR3fK00M61EiwQ6PoZN+
QVxPpK0uLEyeOoxIChuQ24KolYYxdZ42dzG5nsaoYV9EjP9V/gBsNS66NN1sWOdJ+5ngqWbVq1ct
BmRBmvPNrql/YpdxHV3EylXWCL/pRhe/x9cYNVNMn6/y4bKKtRKBaf+W8iIcJP/4DsBf2frKBrpt
lz34H2WziJLiESc/KQMNhzI763mmocOSzuz6aoBTq8DeEgg0NfaE0Up2U2JE4n9GmWelicCaSvkJ
BsuN/ReIQyYQ6kz2YmnBtbFqr0/1XFJH2F2Ev5CQLvxu0VJ3vme+qRfJUDA4uwlAv98Q+73kY0xF
v8zOf48kaGWpTorffKoWxpwAOEnbX4I9PyfbIH9t7ltJhrLlMogK7D5QvzhQQwTkl7oQ0meQBE45
4E4mHmQZ6+wzu0GWSIZw8HM+djBmFmcHX6vrZu4hmiEFBUEZYv+nyeUbfBSKQid1bfb9PUbco/Lh
sRJaRNhcolnrfMBFZPQUoHmheu7mWtHQ7t6NbD7GBxYOgiYEhTw3L1A19aS2WnkKp48QzIL8jcbl
pgREruMvTs3jtihYfQbTfyzzVF/3LrDRocLe+a7MOYDt9vYMfL5v8RGg/HPT8iDjOyF6o6GuczQX
6+81Ru+lodbN4et+E4phG61fpz8vRhfszVPKjLjrxOk4d8/WXCsgshv3/mo8RwP2funkfCWTJpP4
9+8JKumlGdWy/MPaj5NBbsW3AHvBIpB0+grfzt4i8ysGKNe7YrP0yffKu0dZDaJeyeAzFUJNjhfG
Qzjczmi2FOT/qu/sR33EWCtKzCSqRWRzS8geU3Lg/3r/bLgtOoWNuf4SNKA6sorZie3DyIp4T84i
xWs5es8w7qQYEABWa0abpggjzvzgF71SuTL3GWE2YNuMsfExrlVmd+8o5qN/FBfcUIgy9PrTmVgU
yMa8iVI9gp3CGq33vuXT9AKLZGeM6SejDzPXQnt4xUTVnYLpgZRaWg/z7Vfsh1AAvGfB351a1n5T
5kRUh6ENH56kXFY36uMus7F6z2je/3nUOiF1zQZlzok8F0OvhUpNzXEB7Msn+ZyXmAulP/yoRLpQ
UbTvf9IXQJ3bQ0Ed2n6BaZz/+gJCIOas/1GCf7p508QUT7344P+4+WWif3R4+GAa03pjCJkqcnOw
5EFDsxOWH99KHUqz7likMAJotYkxVWWgEFRvCbUuMmGVAKpTg7Mes0kbIwfwvkghc3OZ8lKC10fj
aKprbTbIiDbLrlv5J61tqM8TKsTicFeNzm0rK0HIe/bOZtmYnlCzPHi0ipG+Upsy+sY0k5vJpUQw
M/fp3SF8JbG8UqmnSFFlhRscCZFfOZ+GBow6VRV5h2T+Da9JLDmb9BMSgvPfqAlSA9HvRmQbl+LS
n1cn0KWB79AVAiHCbU5khbvGeSXHQ0mYUo6ivVlOfq0UDV7MOcB6uZfe7nXlGO6cyWzHKQwfnUyh
icZ3pdPjv2mx2LJSfR2LjnQajLC+rRWLUERUvl2+W6lxyg3+N5ta8JpzogNcOO5oAZ5dG/NuFAXa
QtGWUvnsCl8XdVko00j8U8hKLpjJl9wmnCGZ+erEX5M3Nn5Y/gDtcIWlhKPNOkOeZUNeH7DTKr0f
JHSmKOO7+T/QbyvojdClqmmyC65q9RbzyisFbvJfZtCK8TXVzItplud6jLlI2BM3LewQmOP8mkMt
CkYqG4gjZMLd1/KCgPF81u0t9dbOdanmHhRMui5iS+nb9lH58mUB26jz5NlLrkVa2lsbsh3x6w4G
eT2n0bq4Tzaf+50lo8x+zIq17FzPUSUVyqPWvSNam703a/wFkPiHLa07UeDStPWDvV0MXaO89gJO
M4lHGhE5k7lgRxfusAnAGsBeQB4sV3n14r6/juUwpb/K8yltVgymuHuOzDc7vheMgclnNtSAUAwE
u3TTod4px7LFm0tqx+ZD8I3JxXyijeuFEyPtBFUcv9EDBXYQZfZT1dcHDzMXYRJfbwGIYbJieBzT
2d/kTCR5hzWggsc2wkOE6TGyvMZA+hdd3XCB6pp8Gqr1X826UwVYXaIvzyrbbULNzEugeh9d67K7
dkCfg+Tk/0u4kQrpJlbTyIVPgmcp6lcjWUXSmcA8q53SnyQ8HJH6QboPWGZQZUPN8UQp7eblklnF
cwMywcqnanesDYxVV5r57YxQ9lyyVEDm9SbjkRN78BB4uHQmGGm62TG+8Nf9QgDOh2s3Fqp+7Tdz
bxWJpWWt+06pQL7F6/oNGl/7GLy3nKVoqgA5qBM1v80n0o7WHbGC56HE1ONDVTI6kUSj8PpZu7eP
6DiFBQNC5WpTCcW1gLYp5S6bzFZWa7Ql7/473MMd9KH3CG/JDiHci0busaelg854WtZ9ChQYVrGP
DVp6pH9iZJDeLpWrObLFDOdKC3QLlfSgCpadsec6i2pinz17ceFzBcdmnoEZ+BNgXWNtslS7otrB
dHOGFU9ilrbJFvv9ybaZfJiNLEXQuO2Pxl+v9Vo+f810e4WFSRRNY4OZBHqSyfl7GZB8y/rYQDSO
SkPbgzEUCm6CnC7qQdiDkwi+Q+JN7ZoRd4CZLZe4jTczyRBEUIAj0U1IZLp9WMkJuu6aWWJYU/KU
JL/Z/Xipwuiptu2VUJS31vYUUtRSCwwd7GjZDbnl81+XIPdk2Rp867EDAALmP5i8ftLwSyL7BEbs
MEAwZ3VfXQVpWj2y0lPsxzgJFfB9WkzPPOVCYtWJE2ZtHPhtr4+b7t5+6doMlEkjycgvfgJT4rBO
Xi9H5LqTf0u9XfjYduWnbOayjIoJiceZ9S6BChwa9uoH2JiYUMa0TLhI0SU08TKnm8eTgxTeWZC8
AmQMVWKbM1fymm8vtYsqXanFW8NApb1yUu+158ib0YzvYAWvJyFqhnQ+sGf6o83QDVv0aIxnXHIu
3QOmJcvVuJJg+aU4NSoGEKLiZK+5fzGf9sKtYQcJYFY6F6VLWklJx+SwosCqKxK4QCiYtzS+Fuim
JhfquoN1XG+e4ShWFQi32cOzgawCLnhwqgjOSlR3KaoWZes3n27kIZ7vRXKBAhop0VFbB0o985Oy
rcTHS3JzW3ppIezwH7ljW5LFslAx+YhotBtF5PgMTpVh8v9alzS7SybfWfdsSyEPcp3DMMhsuy8d
4fUl0BRz7IqcgFfrFHk+UXVXNYH9u+zdqEy+9ob7XOPpscI4u6DZqo8hhPZIm2EfaKnm0lnhnu7E
g4Nm4vABAtVjfKLkg6qiYUUe+UzA/WIoZHByg1VMzBc6mCKhnvLEKVxdGJcoa1oAoJFxT9wp6kTx
op6ZeXIX2t8qGuhz0RMu2USmvClmwyq47SVdrHnB4+Poq8Atq+fyK0pxJdSGaYYBITx9Bj/VZslb
ZPu3KcEWeP252RCN90PJflai/isFyVF4d48IUF0j4n4nKHVNokAitFe8ryodxt0mGqfbM0DrcS6j
BZUg2xsJn3spzUeH8xUoWoenkMwA9vUYUUFEDAGTOKeJY8656vB4+7gZl6MOXKWaNIktGaU3mhl/
f0ZqNN4x+UbmVIJJ2B0E8QxlkwVVmHUhdzVj+JJZyvY2LcEr8K0sb7M5vjsR1OZSN5NRva/mKE+R
FtRWJ8GuOiqWP1Pi6G7owxrEskeMBBIYvmKBJuthO3HLTiZVRX1SEAXJT+/uGlNza08gdVtMzbUl
d4S+2djH/0dOiTGZEFYS73OR4Kz8erZIYcMjsOvivQNZGdf/sS/VLRGPwUVEToVMQ9xUpSPqHAVc
q8jOcxmHJz8XkKVXZvfXdp/DBJGPmQ02mGhLctzozadB7CUBzx1H1YFr/U1S4HP7T8/kx4QcXxl0
9VQdyXcbdsVzK6yOr2XDizmS4Qg0afPn3MVBpQdMsA+AmzTzZPmLAVeykUY0WYRfgJ68MBRZRFpC
xcEGmHeFnCHJuWslrKFGfgYTM/o+0vmejkEtjxjZROwGT/+vo08vKFDgICss+xSdLuWTcqwaKwMr
VU6NlgfrAn+rb0vt5rqvctVKYZ/v3RmYu3UNmHok2alkzpcsBu+duHsaJqlOkTkfHezvogEs24sB
OHGufpXzYzNhnLiA8OaNVvBGPYNUrnuzesBw9ysi/bu1OftQVdnnNmjYpK+yudGTRjJzR1hT1YP9
VJIYWYcDfZVuKqlKUpwidVPsxXZ5stMNd17dw2hr6WSwyaoqzgqE5NcW8f6dEgLVwl0A9KHDTVQp
lAPIrl5vul176CXVGuRxdSoS35ii0v/UjQ6lVnoPehZBbqaPJ30qFAlUIJKig+ePw7tVCHmKaLLV
gboDDZ+1VH3CjmGw8GjgLTctKoscY01FqH2ADZggOUW9cycKAwR01vTmDUufDgs1ZVWeN1aO0nhh
O6v1InuUeet5fplXkj3fVzprpAYcs5C016TzGX7xHPJMBbCAh0029aaFYEH1gMAV2sdhIa0WZNMO
FMOvJR2hNuwS7iPz4UnAQDHu2iJEvNq48ecYnNvLh/CMuzcJvXd49yihhTzDGilL4FwvMubK3ocV
95b3E/DDt27p/Os+KNvNPpfoELZYp8h0BFNde4Rsi9450BGobQ2k2ZNNMZ9sTfcVumTiy95yy6iz
H4mwgoxbX8rtsXESIZDuXIwQZiuuvbvvmJnD885qN3LBN9lUbvSrMoOmwD5APXk9TSudtHQ+5ZQc
HLJWSDRdtQXy6jqdeugDA0R1VJE7WocX89+xrsiaWqBmg+NyDMXjiJpu5tupr0R4F7h5pbdX5Fq0
M8N1BQbdygMYW8kzNxKSp1XRAab2z9r5xx11t0DDTpfoIiSFtK89JhAjkqZ8zeGfwhV1cdDSAsJK
5nljPjNQrAZO3YamhfxhI/iTW90zQzcryIQLBTDKp8dyBtgZO8xg22Kk6xFFYIytYUr3Hcp4FzNg
38GZNFKPOxPIB0dKASCcS27x3G5dzvBlJ27feMAK6q4rHa9/N3ROSZUXjlMlKNyiLdSZNHrIFASA
vd0Tote4i74YxuQKkyJ82NS3/FbOocU8NvaQlqjdAxU2D3Wo2nSDPC6bNfaMzzQoAejMdqxdBIJv
J+y8Ye5YCiuer1yfMv/szz6e9DvOeOHJ9QIAdeInMC/8zKkIPMlv47JNPe3d9yHg9V3d0+kyL2ZP
SoMz1Aa+kCg7C6y6U1NRlywNKYbnIRW4wZ2lIz5g0QA1iJQdUmBl8Ohmc6mi1RCvSxnD0muSRbxF
CZcQ5E8lmJMKF8bb8IMm5C2Biakl/yKuWh49VbWrpEWJYhu36NWW+xUfmFdB6FV+xkZD2ZYGyjU0
LR+utvh6rpQuc6ebffXSY73/b8BsIiQXsHA0FSJ1uc2XCZVT466FaJJREuQfVFiJI1+uZo6pwtCq
zOGI/b7vFqGu29gC/AyYSfpqls8WFAv79OLiUZFggvyypnVAmO5P2L4C3DN129YcVizBldwOdSNZ
IseBvi8pMBUgUQUBGI25ustw3R7T9AquMHH7XHdymgqRIYt/FNQsTx8uMUZckxBGwv/TZSKQ0LOy
MXLOchQmdbyVDvBCpfCx2OOyxcVpkP1bJ6tuSrn2GQ3IZ91xJGr0EjAOHInS3Cup/JAX/nHwJkuP
GCcDuwquJmHNHUxDzsxtAXDLZILE0TXxn/L7//2b0ssmiMajFAdVC/2eDUB6AHenQPOzZq5ZIq/G
gYdpPrWsfErvPTcy0RZwN47xY2lpRI7NEGlDJsJ+RHjezgervB9+0PuAW0HsaYY1VyXQiRAaH8Z/
RSegMM3oYu3ZVzizkAxd+geChKkQB+w+3wg3JDHdA9GeIO3rfaigGK3Rq2rjeb7ROqq2GFjCb6MO
ctdkvk2pkk4fNkZY4VPrxQV5/R3EOcoyU6oSFtwS03I6pSJ5RghY4ekncOXLmY4r2z3EWyfaHXLN
nWH5WO+eBleLMp4rpJCPqUvwyDsb9S2y1HnVmEFsYr5Hs/NrVWYbRSc8ftQZkdnxMUM8Z/WmN56b
krMkzz4gQZZ8FuVj0znBRPVHhHqcFqKD2QP/UA7gxUl5+xihL6mpVh/FlGZhHD7TrE0ev/leDGXd
G1V6EUQ1vShpWQ2mif4cl1fwHNnCiP4vSF3+Y4KIFHOwdhpguCzXj8FYNoHVwC9XMUNb1f+o/AQh
JMFinFiM4578wR2KqXCCcuX19Y5mnbcYiyQk3Ncsw3fa7H1s8UzNgBSVqJJvN0R5n+fgsksQ4+3W
O0rw0q4HqYx80s+X5Yrjzbf+MttonqdzEOABVQr1ZnMMKtghZgAPV9ZnoDsfn6/Kq/RurvZPwTsH
DKILokwzdWkepkoVqOnXRTPcZZCYh0bPs5tGUg4QwSQckPINV5GM+rfl/dSAcDTils5E+K1ynBPl
BstqvRCDKwLPQX7yfDBQPNI/bU+U9r34P29pcQBE1vPdtPcNktm3sewLCSQdmfK1kWSTCBCjlfsc
6cU9Dtzpo84wWJeijD4BkxKTYJqjXmPdZmwUq0ofv6x3W3dSXZ4Ej8/CwqdxIlNs5HXumO+bDTOx
CMKZIt07KJJo9eghaArAcdnUVPrWseMnGJRsKaIxkxVRt30KWFA7dlYXrBzdTw4pDmMcPRPrOCbX
ehifHQkTkuu7bY4Pb9htr4ZLImUjgAz3M42Szfi5b5Kcjp/XDQykWdMEpJ+poJOD+MNIK8D0bq0P
jlqpDYoTrfmNZlW5zb7x9FEF4NaXT74yTyuQXEGLf2rXEMne5LCwcszAD63wN1c/GTQsVqlG9TBO
kS5wM//RkSfGWogrxbwqDYKmM4210YCZg6Phc+gyscKtXGU+2C3ySEVYXGyDik28b7CNEfcDJ2nx
FXSQLVsKJCZVNunOvpeZAiMrssQUftNt236niKrabPoE8r2PLYbIE/a+lBrR04JvIx45f9bXrv5O
ZoDflPYa1Ow0og8nDUdwTWsFlvNr51TMazSd0u0cjRSvaBllRNl2AaTGbjFsmxv0hVDNIigCMhqu
5mS+pvpKhloZWwblXfSSCcX3pJUQRDdoi2zDWhIZ9MdbFKpNnxvhZe9pRX13a0gjiRHw04rXoWV5
XSwEow3UPSuRsFFQXSnM5Yx6BfZEbLmn/zihUh85uzzlZL1rtAxn/ISnLmGjnVDWKnt+6ahW6ve1
kVhfI33SBzGGVxsjqNykRhkvJs4iEZwG/W4e52VbqQWym3eQGn6inajN+JhS5jUtwAebVd+2fs4S
9FuhFsXQBCGEIySTGKhvYlzIf4JmTG2HpulRFkghUmlXu+bEGhf3pG/U0CKySRRP8pPn/8NL6fmV
sBiQzKbEYHHUlO5726TKc/qxF32VZ5nO6VDMpYZQ/F0ph8jcncQhQSEmipCShxpPPAeqX8MVHgAg
O4A8erAz2rT0Dl6nSjtm8g9XvepeaqK0PC8+I6ENOYPM/eIKQp4IVdXwlmsYk7Ct7mpxu4Hv8a1j
AHHaAzyF8s7nbK3sX16F7jHLdQ1tcrdKOO1wqXlKZeCvVNjy3y65MHiqJ91+kQjUndo9ckC+kO3m
OGyORe0om3nB5uQeiMoEpId+lDs+E4Vt8hUQQ861y2b5csjeThu/28xXDCHdb9LjwgtBDfBpO2KS
+57memV7JiJVwx/Fo6uwxje9watJMsEmqt9hPW6FxWNFrLduoe03/Pau22+O0IR9qhTcr7rj+vuP
+iMyPdX8mj66EZa4vAI3OCGXjY6BYhQNdUZwzekr+feKDHL7JLTpNDqiLRS8eoLLwHue9M555b/r
VbjQ3KsmKOKEeieh/bSnCl7qKk/5+7zl54wGNwarsePd0bQEfJZqtt+W1s+1tW0HJQWt+oQXKC/J
kE6JEqG7B1JNXBgIcAk8O3GLFzDX6ImOTxbCqebjs+vdCmCWOWR88OP9mmBh13PCe7DkC9vF1DO3
yoMluh9HMfAV5BmtSLNV33CNN5WcaUFT16JQCKaGK+h8YDT7oyb2iuaJRKapJyAlv3gJwDSV7QmQ
nHiIvOeHCHMa6UDjZMIKTG7X0dQg+i/3v7Y20xuA4DwjjztyYYJF0mpapaOwKBQMKOZyX6APjvsH
nmi+HnMX3nTWITiz1VDXqs1BgH9WgDXIvpg6QwGaSJibX9qCnjOyJtyCZ2mh1sxMpRQt5kt0rNBY
BcLv+4tfUuUvZ/EOXufqAZFFN7aWKn8acORlQhiMdd3IsG2DtTvV/ZZZxB5dWdp/QLg7gIoWuqGz
lsr2TyyjXuEMfFtgiX7GTXd2apZ4z7b+Fgwxvgt01LW9jQ+WNl87C15P5doeYR9erwUAa5i/CzAJ
yX6YKFsYo+DevNke+wDF82x7K2MgyekPBgf7xMB1Ec6NLkXR+4m4B5MfUaRvKwMPhvpIqAqRzT6x
Y67rkTh3V3PgXqrsggGNywrpf6N+sbsgPj/5gj2b2nwtMoz/qUM7u4h3pVFVxXBEcZZ1gULUEjPi
7F0o456k2Fc6hFVWxFg5pVST1uo+tWn4mYghxHxrkVcuMS9mqNxNsh57Pzm4r8UGMXMCTHGS9FKl
U6Y8dl2K/wjlOkybES2lBGZ2uiQTRhf0e0bbKnUtzVwLNvo4FW5SXolCxLlG5daYq5+RXYELj+DU
vq8sblpgF+P5N1/bYU09PvzRLEOXUPDIraKnTWr7hP78ScToJPjraK3xcccZV6SAy7LbwGdiIoFn
5x8q7ubJmPq26Cb6jk9yMsavs8b2mJxtcSIO+cGBQ+17gU6MkViK/5fEDfp0nASRiJBYTxxQeM0m
QHYD8Zxo1Xm7mIBHjqdXO6rijOaIle9jyYlvwh8rrV8akgV2oQoQNqXMhwhqHLJZxSvnCJFgFHbF
MR+K+eI6NtrCC2S7ejYHA/oaFmcwJBnvQgogaL7Z6/BiRORRYKxuu0oksrgcl3SO83qeDSDgAK0v
svZN40YZ2cs3kNko2r0o0tRIRPZUwLOlcKGqI1pD9j/QryldAlGbxWs+z8Ezz95lFpOHpKVmjn+J
PyCee4ijfdZC22sS2MGL2emDHabYAkOa5RQTpMhMoZw+YB7CT3qz474ohJ7APmZDKJ8zN/4TWWNe
EgUwUeNm3olyfFJKhJCXY0gTl1OHE9l3i3muyGpya2gvLauAw/59P7YfgTflHgr8//DTjoxS8wYr
CxWyDhE62HrVjknSKWgr6GglI0GuCk9BUS25NUIJW2XLRfzKiELLGAhk+fdQqGEfpq7xIyCcslAR
PRrk/68zTi9hEuLYntuEEA1S8oGE5yvLgVrpNh2/+iazCjCYJjLelaZbti6lqm5fNcb7uoeCZjdQ
cjHBxqSOnh8S1MxioOI+bbPuXV5JNB+53meDwD54f2xYlaDQpRGVeUN/l9vBmKUHdckNUo+AcyXe
MyqbGz1Jw3Oe1ueHqrsQipK5I1K/zwQY/q13ZG0pbxsmySQyn7yDIgqC/7OTGwruMKHmEuwfUG+W
NTtcBYN1+FU9OGZwaZKJmY90N0LPs3vuAuE9ZOkTFtpgqr88yp4szhk/bQq6Td27CavSRR4CrNLO
RLcwZ2Mek+jXL94Cs4hCSFloqY7ASM7RV2jWII6L0jc6smdLN12qhzToMd4oBd0G43bVu29hVerP
rukEUCGYpeP8wAnTBOsSkg91Rm1v3ZNmuPuSo9DJEmGy+jQOCMv3ahX6wOm6AUWS//LErSbakDxX
v8/JAKICfd/Zb+qxIR1NmHOnEcn2F5RneQBBqP2eax9gRmMlzYLlPhudkNpqalLyR28AnEmVt6ec
+cze6pVb/g9+y138kMG+Rwpb4FdEhqaWakd88wgazJY0xskPRHY5xkpNGmYs24dIFw2bB3Nc24bF
NyAWvykedA+AuRDchgDHeAvDuHG54Xfa7djCGa6tcGF1coVvgl2Q7Q43FaktEMXBc1WI8txiHEDW
v9q98HPNxZCiyAQjE8FXSkG2DhgYzro/CRP+2Bu7e/6Im3jSAG3Y9cnqiPlb1twKwt3cCwYX9LRB
H+o6DIENh9TRCH6++BD7kwLaneJnkE8IJ7tjeC2j9xCnmqR/tIryH8RRQMjXC6I3rVVc85NHENjb
lOVnbtheFQVvoXGCPrcosCXBq8J0aW5Hzl8aGItxIB8lQJ0C1kkSWWwm5LnGSYm11FDPdjbu+tSQ
yhmRQWXdegQWsFyC2o8VledVx8Ulaj/WQqcOMpUbehJhPfnkSQsBDFMQfIxG6Uripk5q5ILDjgl6
51KA45RRdZI1vY17FDooEjnM4O+tkn6Akr0CixmThSv7hAhIryNNCAj6QzUjtr1TXtm4H71U+zPU
WJUT5PvvZdNsPq+7D3ZlvQPTVbXHdNWz+w6ups5yupjEV36hnQb4vI1F6weG/3SmB18T77i2fSma
WgtkTs4H80K1crnA9Q1/h8+w7gm/5/rbcCOV4VG/61UT01eQxYtKQDvKaxkGyShyldwbPOuCpCdE
0kZ5HOTy9dQixqwAfNFWUtObxM2/pFn2rr/raw334DCR8DykN7BKkwXaJKiOQgoX/TpaOakerHUO
+CLRF/vBwCxLWug0FBUsdWi/AyRfRTklkPusom0jyxrP98mfoa5zKhqxn3aR9PcKljgZ3yOuq3I7
BbIINQphDf82wcjf+QtdA9s4epSx2uhcyqQ3RHvrmVNXfNXpH0rVOZaqtseHH2NfwCLFSvOlMUEY
abLmvvLG85LVQyPGjh9YUKw5S09u3g/TzYxhsbOE9Jo9pwh1uWPpzuWNhpoV4hMgH5tBgHJAEzGS
cHMJtw34Q6Mi/7CU3Qa5gfbV2WJ4xOZ4WnKVeuSA+gpchq49OmhFFieFq7UEo1z1AxqCpKQSVzsX
8wJ6dd5z8JIKPc77uc/ABxJjlhNepZ2ixEIJopGrtwBneFgYAJc6tPReocNtPPe0DFP9Ie2avhBc
W6y5SznXIgFySQSDNWQ13tBuQhep3acBxC7/ki3MCArSSfsS8KgJP7eWdwG3h06qVZNIRzicSzvO
A/TTFJ2go7MWnC7sVDKnOA3jUaC266hqMmPT6GxavsyuNbU1hifbkOtA+vwzmvqr8eb9goTWiJ8k
aXHRiF170O3H752+gumpUsnPT3quuSH4VbZPubYjX2zBJ03Zvqbn1Y9KugjTfCILUd66pYKXAj96
GN2tnz4ui1LOCkiGHpQEICkzVaprPP5zYajpV91snG8H1bQJuC/dzq/5FkTg8f6f4d5M0HLL8fkM
Js1Q9ImKHfZDHy2QJUKMh0UNVbL2fapFqUFDiMKz7xybiZa/9BlU3HEdvvf2gM9WpWnikL7WzNyX
Kk49IQM/FyfIdSNwqzaZJs0isYCb8mA09i8SjCSJk3vV8QVRwHNNkTVGCcxyLQjkVa/Vn9oa1qa9
7llbZ70cDIdEozar1xYIeDCwYnfSA/t855lV5s4aNkuE+mogol6hs/RhkScCjuG1RmqkhYzA6RNs
qP49+8q0j2Sdjqzh16lavQq2EYeBm9qsteZpTYYXh010WtP+1UFJSGc2zXgGq5LhZZvW9qwgrifm
TeJXftVpYStmWkFYj/0Djy/3ORHJXrtvFNNNyJ6UzI90ssO/CrWfbMT4GqsY6jf5ivMm200dhKoq
BNSov0mo4F4KCcAVJb+Y9JHxvIxcn0tyYIC4VLQfiquRPNTsOfWrkmgNAv0Q1m6xysunHp3aQFcy
LAP8XvR+DEwYG4VwXJxtRbBp3YnjoB1dEWBubt/WJFMxsEYT1jhLXq2fH7j1Js/I5Wd5OpSoYvjt
ZfKtPSUsZyMcRp3Bg+Mk0EDdeOdKTsFekaZNd3HzYgZ/zNlu+Qg58zeEtcZ/X8z912a4pLc5ExI4
ps1gllhBoIUeVCperCEsOGTq8zbBRh1xNrWuB/9HXoJmmWTbBBz8DUzr5o4xMpZsmpTVVAao6pRK
riv9hh0AdUvfs9BjQMMOd6MoUmUbM+8iEOrDoOT6Wipy1HsN5HmClhncPEz3bIkMBrPaNeRCso1d
8wnew/5FaajW7Gu/Mm6cK3UJOviSJExdcPCXgGz6F8DFLGVaA6uyPjLOCVoMx+KZUpEvmITVIcng
cobaIKoGJRM8s4eGuPjgsCWObzg5omcJFYmDZIunPBgDXlj+BILlzgEmDIhtgISQfzyInqwZRIcJ
zEDz5vL5Yuelf+E+oxlBEb21MWtGJuSB9JSVcLOZLzp3PdjRE2jtGRZ1yrdqKLwxRp3dpnOkfwXi
5K07/x37qHevTvTr+DMRTqu7uE36oeFA8PDDHp2sQSfG8w/ovwj/cE/YgMVekgq1tDqC3Y++AKuW
aGGZCHsaz2647okBrVQWa9L4+Bugzj/MzpOAnhunQprUd9dmr1+pjBf3/ThwaJeUVTzU44hQrHw+
nOvEcOKXPv3sAkIpMYLdoEpjc/kYZf5sovqxxDNP26sZbBiDhEwBk+rlvtedaUZAt5uzWyTrJOqV
PLj3bTWbwdI88YvblSkGAI4MRmtJW88Z9NsOIdauBmYEuJiCnXovTA/p3LR4Q7S9TsKGXtv1RRMb
HEaGGCeo7EOJTdp0uuLZ/bX1yR3yRUrgPuswusTSwdFa4M3dGhfk5lipNXGQsf13AKRQsGH6krmH
QxHcbGjqaA7bZs3LLgfpmHBpkjQulxxbAJ2/Hr9SboloCwPj8OhAYFEcXhpaiCXGwTiKJX2vv5ud
VDR7LInBawDtMt/ne0/0H9cmB0VkH8YyEutWr6hqH+AmCFTTS2e3nlZfw6rOmNBbXGvhHstvlHOu
CgTMzqH/ovG6hmrSuztPU+IYrLtXBr+P8t8txs3p2IUDMGp/GdNjhyxXQo0OCr2TixjCMdJYOdyq
6/HzOAgWgGqXFuXclMRtWDNHuXplXXFvgegVtTeCa2R7lJVU/siY/66SRysNal7jgrSFdD5V8tCC
DSjJyGntOVOCtRejZbapff9sWvuck1ruBWUPgkwtqZA9rTPgByYZ7N7HqrbxP64Qp7dclZ7cgXGZ
knga2DwGMUxa2RL7ZPzljvH/1bar1BaO1YZaSXzdlyXQyNtF5ElI6xaQEK8yHf2WFZ2WybRrDAZr
1tJc1BVivUsHMlNk6/xS7fW8Dt6Q98uoDyRfeZcrRvk5WGbYvZDsykk2lFdmrLrZZKtxDpgyJmi7
gsz572j3e9+90EmsGPOO1iZNCFv0aDzFqY/9c49guko17ylwWK5D+ftOxgl/z4lHBcYWvsycXsMZ
cXVr2RE20Pf0HkdMawASKYR0gx7SR1WtXjkS5Nvwi1AdBCCMSDeSU9b0UJ9mgtqAh9IL6Q1mOUOp
yTCOKe6Yxgnhm30mnPLCdFCWl2Z0/n0HRresxNH4EIaGx56f4v6tyiMWvaz55R+yUJF9bxibXPeJ
6pRUma8kEC3FVuoO+TvwGY1JAphIbVqvquPacBCz8z4qGKPhm3DvtODWDE21w5Rd26bDlUKBOKYC
23jB+W5sSPAur3Pm7cqIv+lQhZO84fmA4/YwIGoXyH4SHzUCpezHilxFCFDlHYvYIly+7Vs2UhhK
kJW+kWzKbm5MnpqsT0Wm+rA3Cmot046Z6YkQkTPb7uo0Tx8H+MOzJdHVXxDI5pqsYf9OiIuE40+B
tPucCpo0gFY93ljtnvGPV3PSYen+iHARYOINMlpi/vzsfufrF2WDPdxVEj4S8yaDhQNsFeafiMbV
GZPYiAq5lMzAT41X3taHqNNUOyOJbGu1Gb0Og6rrmuadckKmvvMPgtyOJQtYpvD0zwnGtyGv8bpj
1sgls8/OgVIMOna+EKTxT+3U6LC2r8hFw2KYrOR967zfrex+tTDqqUn24kZ6G+duFrD/joBEr/wV
vNOV1XVm7IRJXnoZcaeYvaH2A0lmfV1HbZR+OrRvoHn7rxsseU8tCRFDdm+5bu8Q4drM98mthH5N
90nsd+ot9KMvX78OdD41rKPmPssvFLWmNj/KjKSKowAkSCAsu9uMvGPTSNa4KvUQXLAprdL/FTN6
Ka+FHWzcJIBX5h/QZemg0GoGOPQ6Yd2Lsq3vUWpZoSR05oKwwMcQj9dmRrO9fKYbIT6MhOExWl1+
xYyC24dDEYCqVTAk1Sgk4mVjHTqT1NvSISgu5rg8fs5Z4B6MiFLl4ey62tbtoJo5Tc1iuim95JQD
clyjM6ht7P+3b2tQ8QKBPlvamJqQPr1bCUHchLYFObKRMl61fDj6/p9SstrV3LSYtC1DR7eZR7XY
A5819ZtMbFU/UpmLMEj0LCsNMuyv+tk2w6va0moa8PhaWsaM7kgaCR0raiy95kQyuQb5acJdgomk
5Ix+kP3UdSTIHm98nctKdhQWrSMYVJKlOe4WvVpVmSFx3c+3HKCETftswEscS8pgF/WFiUMuJceO
aO7/O3xzR9B1S7jeL/sonQwi4B0zQdw+kWbhCnWr1tvfO50dtYLIuwCrbgpi3CxAvskKwhIMrUVY
JeOR+2A+SLs1WrdBF3+mvKxfzsFS6aVaic0lRlX1WAeZZsyxTqmmYmGMnVkgbSBumpt0+7MUkS7Z
5xuRMz0FhkUf/Y9+0E688SOW1JDeVugDPpXq9X8uZ0czVGzWLnNp33aMvT7ZEJ8jdRhOla9gc/S+
Sa7mPzh2hHQPMheeGDCSEAuH3JRhTlEm6pZD8Vd8dIfOQhuBqB7/XScpbfxxUzy8Pfg92HAJwrfN
5biL1Pfi6/DoIYJ3JYsgR1Vhu4yK5lCwUXcyRagFyRynPjCvDKHdcC3vJKDYc3y1lOuVIT5wpjqO
xz5DteVSLKppCIdo18X6XlXMhFtr8nxlLhww6mawAtv23jZbmYAXgca73RLy4gPOkn8SXT+VNZcA
7N7Gc23nm9ZAdV370zRqT0dmbAbuKLDYtRKkoaXgnZAFfn/ENOjMwVxYjm2EJM1qFiAdlsipcBGv
FMyoaKGV6e4MOAEomMyC32thV53dTDGc8MQeatRQ/PhYPBKQWU3AV2w7g894W/3dgsiEKl5XRxu8
ZfXdvm6k/bA3OBFmT/C11C4TXdRiWPT+uKZ4x5NaHJ7pthAJxMIOWjiWZ0kbnDDjhpMDeiZh2l59
offu56YK8zdRipUge1vqe72tZ67ahNff1ICSRW15FAcxmtoqN2ZATY7Wi0p35P2IZUzhOMWzHPnh
XWQ8u8DUlwLFAqnwNkJn9TROGw4Z3YUP0j5Q1FzSH/WZjOe1NFzJx705/rIXiL4oR+puw41t/4Hi
rt/NA1sgl6at/jI8F8t8673EDLfLzHTmBH6Jbor0DuN2YtMfjY/btsfEB1Pi2YifCEA+N0kN9hrZ
2Jxl7F6edqoNeaAcPXzlN2c69KCsltCT++hrHou5YyfIUebFvqmQBc8q3H5mMh+cBXIc8ZGrlS8d
11nFAjpuLgmMgly8lC3RXZal8LqM1koS6P0ERoJ+a9eYajM7zIYKWiDzywi3z0+y7gY1Vrja6oOL
r2iMHRM72A2WIKkvydzH6E+WLwolZU0/1sxwx3Z6BoX8jvYI0sh9uDfyxeR7rnY61CoMS7fa4uPX
Z8wfjDe6FHTYiSjs1vyhuRKkEL7IkYO01aB33d2uKW0R5i+bTe40Lk7EmxVFKYbp70I0kwST8Wkq
LSXgoKnAydcp6BbObwpS9wDnojBu/20Y12EvtuXE6V3WeVhfy5OAwI5tR0eIgUjt6rifQrBh4CCG
6PC9y+9z6aTYxDpAUby84epEdzkOuAN9QRJR/u+YdCxKyebFVTbMVPTwBGoe13OTQleYmaWZOIrt
sbvODMz4GcQ00vPSt86wdQNjRh9f3ZvXvzqnOY7i4IoeeDPyoaG3x9v0whR/NBE7Xu+gwSJFGHFC
0eZwMKIlbeyrqAfM6DCu71wjspYRImvZqZVAReauBIh1bD8qm4LIyA6hbudRZ3G1rnVtvyl5nNhR
zzyGR5/2Mk1QqUr/ijpv5ruZdbqnDKjZZlhNATQOgCjJl4A8hCWJmEopfr4nNyvgUGpikG2XKX1x
BBZgIFAv85bFLebtjcF7NyRmBgXbZE4C12iGQxbkqyHCJ6HvMNtlKv0r17t3UlJHC+g3uaQgT5Lo
stzUd4ENuTkvozaaDHj4zHXpUv6X3IUuQM7W8F7FTT3ZAg871lu2rVF8I4+WFBZZBpsBhNJ6NjGi
2rSPT8qBEb21Ycdh/mM1i7RlsBbeAzrR4fnPVABmaHxoJyHBjUGubKtUyk6I5+pIqGSNGj0v3tDV
BFlnIyvT9f1HNeDOF/ZKFQ2SUfGYrtoR2bZDOAHvD6//4vGWREdK4k0X8ZwQ/DyzOfcr5mGhVXyq
qFMmI28ymeovToFr8am67XYt9nIxDWA4qPmxYETSdqvdYWmbRodmeA91hcz5c0mZq+7rf6rU5tGp
4I/OUhisomQ3SerOhr/hzKzgcksAxG10QNKZ4aLSXDCiJ9x6kRAoR7aTxFGoH+ZMososxtFyKE/o
0isGhWPylGrgLbHgfXFsz/JWOP6xpZWcmSyozXGmJpHYC2cYUi0FAWBuDz7r4zoMIZcjgs0yTWCD
g0j4YiAkQSBVtFqa79lu8NLVQ2SaQGNWgijqyQ2hQ+hCdRXDtkocQsusK55k9xRVav+HKda+xeJB
79M0BbnrPKVUbqxSVM6m1uEodx3AN9v+zSfDW8FKFC1sSjZkfOhrhbiI3LH7/Sm4BHbzSVHE8YlJ
6pdY4xBZ6cmFG10Ov+WPsUoCwjYb1KngFt996kS7aR6mt81zGG3VzrNs/bRuFi90XcaVkeh/PTvu
qArh/FWgYu8Mv//tTUpbGoZtvE3tiw/4vMDrVnnhCYQv5xnvU/s3RxVSa5MiP8gqRwHNvirkJG7I
uHDHHHgThIjktTvKyvFM4lKLI4xCCHjccdn1ji2sl6/88Q/VVh2W0XHrYONdCSL1iviBBl1RO3i3
6hJW53BB2WLJV1XBA/bB7and3VGnH2s9RExtf7y1LU/Czidu8Xd5se5hGbLAmdcKpSm7mXRkz6O7
vs8toKTY0VG5cYYghPQlrTSzp/O6Qj535sZDiuWqnzde4c3MG6Bb5yBsKpVChHH++IBkIeHlRvkU
qbVlS8O8eUowmstr8aOZoD1qiorNkPGs3bg73NlButXOamSHCBjrnohZD9QuHj4Ps1V483beMln4
DXaWAsh+WLVtUwCrpKqM38Q56X7nGa+kjNPpY1EZu7n7LJFH8AMkjVbmjriPJjmmTSk/dSq0Shp2
e+YwjvV1ObZ+5+e7AFNyNETGbGqoFOzkXmCP4mzvwxDNAMTg8h45zgSE8H6s5dZFGY4ZB5WgR5v/
TKM6f1nmMcf7Pwc3h43B90G/ckF3f9YuGpNSD7nLaAM86W8tUyerDrXePAKHStw2JEAfKzasgn8r
BT8fhbO9zt5ysdD1QEyJpsmY4bx3xB7TP8xKs0v9389wo2n6zM+1ZcqDcyNuz5A5x7R4ZevWmbMg
kcfrkLE2wZWvR57fkmTPKazmfWazGZrcKt6EsG/BnUhvsQqdb5Q7Wy477QHTIbwaJLHXXDREkwH+
4/tg+DWgiEEyebJf5GIBFJaQyg5DWeZ0JWaMH0VkkVFT9RtGizk+7knEeg7rJLCF5/tcNYGMpoIZ
ddiOiOSRLOthH9Ce47b7ZTsiMlcCkEvDVR1jRbxnOVsvRra97FSEPwi1EqsTCPazu4MoeGVMRB6s
WOo61Vf02IbK92BeSqR3YG6p5vHbpCQ0mc/lqIIuoOE26AsfUBUALuo9UwkhJyE6HDcYGV0yeibL
kJ/nmumygqQfnv8y2BOrcupNgE4SVw90nAx79h7dxxEqGD5n+wB0YWuh4FGwz5b7GBbCd0laidPL
b19uLNDPPfpWW1tTEOgY1TzcFClcyu7bHZScBFFLaqV/p98yvgQlhLJmxzq7hZ4bwVbEy/YM/rGZ
DpbGxs3sc80B+OZUFRIUCHDWq3MXSTObOqmk6mWi4P36azviGCO1ZGqU/nzLXa1CGFpqd9/aBcdz
BrPtu5Ef7gWYgtn9ZaIELstxStV9PyWyf+rgVycUI3tGJYusojeHu5kXnRCC7sYEYDVuYdGp3x8Y
qu/o33EWi+RIz68Gc4NXm9hFu5o3pIbpaLcWQ6RneidQpkIVxgUFgW9w7Rlx1xpFgaldirwmSKUm
dS9pZw4Jc3VDfVFSoOXMf8+OqkkBGOm4+fKm+2cndumtQSmzzyPzY1dSTYt1Rq5YerEdboXbisXD
K/sTK8zUdcth63aG03hTvK4w7PZ2yqleDba2TqJy/ZUbU5bmmBZZYpU1zhGeqyEpvdiyloZ86DSx
FNLCR7yXufN3fPawjYPcMiglBKmyrHzcCzjbpEofl2EGun0WXfEnQSa7Zt20IJWGdP8K7hpP9psc
rn7R4WL97mguxcl4Pjh1b+mme+mFwPnqJhaonFs75FQw/OielSRwJW5ylH/IQLRUDOkHJmj3j7m/
MmTWEQWB5LQlMr2k7bbYbYu3ItG1mZjbI8zO7F7T5f2zKoCxvQIVCP4sGx/KVI5Ndm4oRbeD8X/p
P5mfBuSfMVa/uG+KyyxV7M13AHg+8MuP4EwN0sMkR8wPDA1wBjBxM7GKRDd3AgubtMuR+G61yNIQ
gZwzXTzfzPYfzwWxxNa09wZSg5jfw19riH9HnvNT9iPAixuav44AHOu9lPilo6uq0SQjX+2tZFU5
r6MFgocUMk0d+vgV7BSq5A5W9/ltgy4kbnRyKzvO3Wq/PAqGNldOf8B4s5OJg6m5zKwNH0/0/mKb
SqkZbUInz/Obhw4pZ7XKEyVlcL8Guo81AAB1J7tvXnfR5+rleh4jnRqxmjZ0Scu0Fcyi3QyqloTW
9GHDre9MBo414NMfWBab3/oef5XBnsvxurDLm8c4dMJABYrd+nX1Cg53aSSVz8Sk8Xq+IsUca2Jq
DvFkHJA8Rgt+MWVXdAF5rCEtj0C/u3a60LNCzTTacUyiGGooglt6TwTUuGj6psFVWNS136rjzau8
D0gmXQwmjwtQqy8CGIHLcsru2w8cR+AS9dV8BHwVex0ekpiRNz4JHnI8IkdGkeAzhIWmHMhKXm5w
c1915JXi0nOZBcve4XeVX3xcG0aGB4svDQmf/NpVLyffZ28a5qCb8jkoQveojqSdXiYcu3NJKIsk
kQm68k+M4lTTgPJhsoc+9YIPPN8gBxAKdbuoeO2ou+Fjrq8qGobPrPpLMTL7XQyEUgIfJvkumtpw
//Nx9VeYYQSPKkNzXJWWzIr94DxpC6Dn7ZLshEWyFIbulRZ9yAxwzMstH3yv9g6pyPfp/4gaqxIC
J1rRk3A1fK+20zUuBdiLOHY14kTkTnCDOEpp2HGCqm+9voCVwqz6J1mmPe3csKOWpuZ/4CbG71Pd
f5pz03v27WkfN5PEec7AOFhd5i6BYLUO/6ARLf9bvHheErjnSBWQz0n71i0sXSnAYZOuQ6nW8MUb
H5rPCZSkqV7QMbEUe09Ur4gbz4tkFxzwy447A/ibrHeE/UdoePVOp4pEZU0txeYu6FqO7Dj3Z3fy
Xu6+AAD/4vc1L2IGmgEnxepgAd+3U0yjNPOFgItBsLwNyVGUf2peS8YkZaXA8YuAf9LsnycIn/HT
3Ez71D55TCK08Np0160ToXF5wPQ6IoH76JVzdsWSTJZ5Nxnmgw3QCn2MEFoYpR0V2z+/zeK01eVK
xwtQXN/pbHp/kPSWvJ7qh3SpteJAgS2d2IJE3qxeSe4tj7AA3PzbXNUkNDNwe4h4YMfmpA/JbZ4F
OP5Mo5nGvkor8xaEmKsncxycFzTBA/2zxDekxaEOMFootS+7e+nj2MNUyrS3HVuEhab90gGVfsR3
WJsBRDDN5lOwmv7KbljWGGRLpQCkcEw/9sxJmvt2+FVoRq/gH/4aTM1ML0TzBPLrdqsM0jr0jTi0
PZxFpQfp5Hii/W6rOvIzKf9tfcuuS5n1J1vLY+KU7pemx9IomHXIGynMmOEB1XAIuKCD0tRFLEbJ
Qd4v54sFpJHFmZcH1F478La+xroWN1xzWYzoDwdx1yfowpU6oibW+HUGRK9BN9i+PEGWb92jYTQS
r6L1QoPTm5OlYjtBZzC8YSsdF/2wbcCeY1eWO/RpqjjMCGBxSF9ZSVWSRkuigWaDiuAnOFVB25z7
zTXZMHEFSnk8d3zCcLB9RWgI8h1Lp7UncCbIqxLdeSyT9mOVwOdHdK/ajskxHsmtYpkRAqG8v9gw
bMh/0O/KqKgT5AbuIGtwbH2IZp0j8OJTFGJry4CW+BuRvxfsuiNh3E3KJuHMyMofKXIxHJU6EEtV
DwiCtU1Db5mZJGUvOLXkuxEBVj0P8z7RR/LpPIawBMCOVau3Eksc5x5R6WrWK8bXgT8h7AKYmX6K
7NZ/3StdGN8l4qMVF6yJiSP3K9nS9xB53MPXZArPoba9ar16xAkGrZ/BzOjCGxSTanG9eFgIYzN/
kxInBHBEmHbOweamWCgmcARCgvfs3PaPDOPLsxSIbK+JWM2GHmH4Tk/cEXxHzFneU2yj4fII/NmY
ikUiTcH8zLzIEhU/OKzqxnoDIwnaUw3XDRK7fUq9C8orF5yp7OMLvQgD6ociPhFbWyN7C4hbJiS+
/WTFJU7Id/PBhEn5SkD1RwpqhAXuIi5eHsRitDG05dvqPWNaJJv60L3zQqMJx6xwiWhviVtaE615
yNQ5QGOP1wmVIkA2eMuBu659ptvbONl76hOIdcBG6Fja5z7PwDCw3+aIp0VNe2TtKcDAOuU7cnUH
iiPPWihhaq+Usr1ZidMohKOPhkBRz80qEY5ix8FUNYUSZG2M8UPV4k2HFWOX+4QNVe+WK61ICdXe
L5ncRBaISosI0/sVa8Rol7xQL0bzfVgFIL8Xx6ZBxDja+KGtB/W9gjFm6dRMmw2zGghSbZMMbFB9
x6iy28KIH1/6YXxjFsLSrUv45WTK8tZF0MFuWIEPSFWIe6akQMBl76X/gV3N1dES6uIz8YDzx1SH
fRnoBX8AUpp0VJEulHbIv7ZGPchdqCDdqoYA/EPHOiRxdTSmzityo5TJnaPWrkk9y48gWPlBe5LK
0o0Qu7Xtp/dL132gGid87YTcTMZayfGK7f6osKkAi9macykdx+5vtbHdlko9sUjKRmuQr/zcVkWw
AznkeCbJlqfr4XidIBIs5U27+EmtGq5sVh9xGhUjFu8xd4PNC32Oc4kF6Fpx3Z3v+PBCIDrDu9Sw
Df9favpM37ST5DG9L9Igxpz5uwqYMVWTQDmT4au8AaiXvdhhwINio9aE+mgUCtWZhQ6XLgXFB8lk
RVVrYa2UfVIL1nH9wAifpgPVp1sF83/i4PKwLyG1i1Lux3lwPOpNVlQJm/gkwqa3dBYstXqCFkwB
lwmvE8ZCuGQztpxPuUVdR6VA+dGWyENrN692qKfojz5xGeUsaJBCaMJyxTB6iEpQJfSwKT5MrOLN
c3BlKBGB7xftAOSzfm++XTBID2JU7fnfjLk9ehwlM2vZVSCqBkIYlVe1+fnb4krpMufi8PG//RBg
FSzxdVF7WFh4sZD8b8RR4c2oocGr1EPqon5ohWCpy3aEdQBGg4t5qq6FzNpfNlcyNOEXhkDWSxkV
76zwLXeLQ42skPHsQMO1n9On5kjomq3YX/LkqX/SLC5icgUlHICZqG/mKp0zO1eQkgafJ6fgJZ+8
8aHWqrksQpKfID+aRsA9EFaN1Xc1Vh63VpQQ8Pe7B2lX/JphUTNjiITEzTt7nlO+/t4e4PXZ0jJ7
6SdF8v4vl10X/Jg4iqA9eTRJrJjMZc8lXkCvsAPejk1zRt/W781mQNIKbsPf9W5P7KNSJ0fGtR9H
dbvyLKtfy3pVqwFHtRnLsAKTKmQQcvjzUGTCp8e7dB2UHUMh/TFY547uuTDegcd4iFG8UPM53d21
bGiL4bj5LQzP0BnIQAiBCiJmlDn8QhxZgCIC9/7Ss+xZTSmdKpQdyiGEBVD85OxtqYFzXYva4Vzi
mWZfQtwraHAbszKPpOpXDERSkGsk7Mv2R/YSSjE5HpFtMPkoPVMjd6KiiZy8DXrxdZk+zG13wOMI
oIQDWpPmSmIWDlzbJjw98NRh+e8dVDWsL8rtXvwG/1xEhcDIfZeg46fog5kYN+YOSuXR/hpHXoWu
VYcCsHsqb+TKruVpdwkmUNhGbktnVm8O4W3WVj+Rl5m/cHda8h3Onm4UD3TZVlNkrYgugY6cJgWI
8UeNM/nSpnxA4p3RNvnjb/O6z/FqlvK3CCUsLH5GTWjilRXew+YR7cG1iTBydWbFQOw5X6fmRWSy
RR4rq+s1eUbpkVWDg2gy/K/UOIN0GDR8xg2Fc2ai6vxnCF5fQU3yDczHsZrl3emGLDZcvGLO/c/H
K2pEElliYBgl32uhPZR8HhrM44ODcOE841AmoCfES0KfEP18mNScuEByskfpl1nM5P3TZzrTvs2C
iDbgfEV3fODgGInRXyYBXPtinoM/tv6pRhjJNkyn2qOjIm7zYy9Y1HFyLinkLJanT2zGIZYySNOw
SF4Il/eCBaWH3V1OTzde1vmtrNBa5xBQpI3wAgUv6WGG1glYWRS6NhEVwQTyYbW6SjZeHp9MBOCf
zpO+JX8AZ1lwe7pXZ+xTTLe3LAASEHVAdmbcE2D/4bAxnwR2nA1pUKFq62Say2Rt81lluNQApFi8
+lfpRal7Gr1mrSCiR5Gg+GEfy8l3lSxDRZLtdq0QogJQumyLtuoyL8yLfGS6bR4QRNPSs+dnOWUl
fk3tTHJW+eBnBeZIR9u6/qcPODpV+p6ypY2m92aFiLA1IOz6Iy2l3Su9CK63qlVv2h3qcv+YLS7b
n1mPUpQ9VVz2zatf3b0RsPTWWv6MOpzVHRrZdN2HoH2IqBOFh8SYir+CAgNQ6FCSHWyAxmNQ8C01
IUhUR/QY0bfuEWjcgxBCox9ppnhZ6+XLcal1ZV7FFEv/8zoIGoMojVAVSoMSStyjeFeWFSrMmll8
Kth8FYuJbXgKCNJyOorO3oIhp2eqpmLNh6CGM8zFNlWOXs1XreqzffPeGJ9LsWNp4q5evaWn1W86
Q0P56RFGW+sHgI69hzrvqO8ubhJmOaip8agVQPdFc2vp4SUUz0Fn1tr7Dd2dD7Gn0PnwbSPjHmv7
LhGCqsYMjulkiHpAHcSAoG0kPjHPyysr5TGJgbxjpjzwhUiq4ytuw1QMMh59WIdYfKieRvmqOuOx
KRtGx2bo/pGJOcThPazpB4jNcx0CXrxZQ8xw/lYFYseXes6Z4hf6cuBGtpkU1NRbGS7ojEP99xSD
VV/ggyZKw859tWqdrapOFRtdgjEkvBxXzmJm2szFYO0KXjRsxdGiZazHeL74fm962SglP8WSzCIx
+d5otrirGRh8MHZSkDbOq5iXZN2NhmEim5Lb7CukV8W+4yBRN0gyd2qWdGf99ZCWgWlALkaW4CT1
ALHNIRR1FeV+vp+Ob1wRxytD/m7aP9er1SBqiu3qSJDjxy0hpWwgZHZgVQB1Udok4lQwXlo04NdS
6dLXZ/IUQCvRYHvCzjlh840duwSol6dEtc2FdlURqjZ1pOEfosvgqA4XQ7icEy+btcMnnLUKM9vZ
63zD0CYpKNGKk7kaQyqdifTxxjKBf3YsoSCsJigvCypxAAMWEuQEfxfk8zeDWC3I3V24C6amAOkp
L15pF8s5WQnJKJLEn2DdZTcRcgTPyyXemJWW7ipvCYs3eC+8P87goLtZxRttJa+rlhCZ81OPBsul
X8J8+seLfvG8IFr4sptl1IlUOChDmR9YGlkUJstVbN2gC12U4zGOkezxYY9CPFzpCuV6IVOd4q5g
biKTxKUSvHPoNhxCs9cDu94ayzqAwQ6rozzsvLaQm95lnHFd693ldDFqaRnIxBdpMmzfPmTr7y0X
Ls3sAvr60BvWyUCYi0aMZOqzk58e9NbR6/82to26aK148VBZvrXixWUDPWIBUmn2q15fuOjNs9QU
nvxBrdKF1uI5SfSC6MHlQ5AFih81rKw0mrJEsCGtIDGyHY0+2oDBvcEbP4KK3+H/YG6rZV13Qjco
mnOZXfDVCQjELtOFBwQHApMqMoK8IJgZ3IWwCduTiyNnQ5EejEbWvCa4ykFPLGnye7VApeBwpnrd
lrLDKWiPZnEaRVeF4+2Cslc2/w38zdPn4wPYqiO+KlCVaC8R0zXCYEYQdfOVWI+sUj0ivAZJ67wM
bUIIxA5Ggajmxi6voCFzH4OtNb+roKzCBPdENT0wamdYMbuLURv6Ql5aUhOYpUxwcgqWowNONrdg
nUJM5CMjFznY1lL+sZ6I2XS/9xffeUzbMEZytE8d1u6XpF/stycXavMG3ST/adRRennBPhZ2oa/a
R9euqBdUaw5hURIDD3EnRxZbLzzAvEYUyElZmsafGitLWWlltJMLlg04zRDRtSqA5Q+88XHS4mz9
9nFvY/ZPNhVGUtcwM+dhhuDMNoEpr9wUIaWD7bMLYQOliXtc6A573k0JaIXVq0o7rf54JOsi7GPU
p15UMzVHwFqfrVM4Q3J7akd2i5wMwHnhyg05oRAzGxbcVkY/+TXu532fsYhrdpvRoRIR0WXYKcX9
o9//TYwOOIF8SVvovLqbqwh9TPXTd62DiCcbuUxefcl6mxaSiGq4/pFpDlmuotrT05ihicuFJhn+
ti2MtJNkl8dQLl7IEjzIF4WweusiqQfU3zLcYwd9Vd1Q7Zv6RLA3ZeLoIqcKo/6dF7Hc3OeC7bxb
tWhHJ0mXdjS1BGAetbNl+r45C3r4QUyytNmrqF03cSd3Zf1nQr9iFuhQT+UCbYN/IPX3VWMyRm1Y
N1afAt1IL9+ZnsZl89JYcPa+VFNo27dRs0EoscRTopV19isAS0jYUOC7sq5CqCxiRkyvNZNA5ZL1
7OhWgZZqkRoeZlhjMoAjB/sAIHPUOKptAaLX19v1vSbiTZcEbkph+7qY2dcwGrreNW9Jrl0S2CCN
0R294AHHM5KtkZOw1hcGEcxtEoCvmj7ONV62ZtpqYVD85+RLKsOXkHLFwQd9fidqIG8vIMQoLEUk
5sRiJqnOMsPw0jfiTo5rCrHQSobftJakTydBe3QRJUZvvtI/FpnfIVssSmHbkklBXKqBZIaabees
Si7yiPMCxHCwJnVSGtcqoIUWYffkbfkL4X4mn6mDh9Y5fOMgsDaqerlRnF2Ste/qIPC25iOCzcuI
i5SvZJkh6xsErPw0AerbAxIb2CmtH2Fu0UEVumnkJ/M4IAU1ZMMiD8Q0rV7I3gzfLaIAK5TPbO6T
5MgQNqY/mOvBlR/dyl0K4QOztcf1grEMN6WfmOYPvXgfakPJK8fLmZKkJ7iEADdBROS9QuSFmm05
WoQezJ5TS+lLZ3Oxnb4OLuNZkVlCoBqiCZQbgEfhvDZz/x4v8ejRFhHaNzg0oO5UoDoHwdmz07tX
Cq334VFiSVDtcXja7uYFj5aQhjkxo6TwKT+RI/pegPtJw+j6PqtZwJMUKNlwb83bDuxAMz0UXgPg
rdpXvzR/5voTfhncQ6I/nkzTwPGL3owfidK/T/vxB2pQyJakXrG8twOX92ojZto9A6UdVICYLU8v
6BzTVIb6PRkGdWkdJaJWVA4SWlUC2cbJ+MYaYwP6ODAe1QqXtg9pHRuGG0RVgr+JB+z0K6Qc0yMM
osAjllZ1MZlH9OeCevE2YfKfRjRnCMx9RBbYoIX4UnaXyraEM6Ssk+k52HZ2eNzWr/ijC6cSwkRm
wH9mVyd4GQ2ZacZTUDjEVpmgNw0QJdR9bZvNQSbhoZsFp/E/C4feYqoI1ZPt1IYge1bvpAzoIFxG
TaIllzZGuXHJO7Rk6wZ6ewds+Y9NqoI5d/ZU5sZvd9yiou0lr/iGDHge16WZcNfq8wNDi5drtmCg
N/dtVnW09J89Q0MTuIBhNzRsMIzpylvohcQw7ctAudOy65BTgrTK5wJnk3RLjVd8W2VsY4rCRV+3
bcxks+kObVk04fA5p24zSP25G+h9gDSnUsBazFAZeyKFSW3iX1VB3Wx56jsj9i0diyfDV/I78n5a
chvmUO4/ZNmD4NrC5aifY1CofTSEmSlxLaei9e4SGDdoHUyRb/SZpnMHNPSLdMqF1uv0ZkGCWE7a
6SMgKmJPBcFJiLNsu2hp0fVcB/bWNOfAI3ovNpA4pPI61twf7BVLncViJlUnTjPYC2J0lLr4/CEx
O/zFR4L584tnkNGakaGDuqoo4C9KlmqZQz4SzV6IgcFjLMsZ9iGgtOEFGINnUiSb16Lir5g1qaqE
ayE0UfaEu/lVutOBs6TRxTABdeqCmhYcxHKjDq4DdVtTX2OxtymfxkqBtqdu6bPPvWK/4fVmvd1B
B14yAhfpGJAOcYIFuOvHQSg79BrqR+SOzgaLN107qzQ2CQC0NATYTm15x+Xj2PrTSeBj6o0+44cv
cFHgQ/RmnJ84WRe4IcM0L8GU7CIL0Hm6uTOditMLEl9kshBjtyFl2JUcHCf/+lOTItfAS5k74E66
+1t75S9p8p+FIz01bUJ1qXlPWi2EY/ATYX2PEneMxojnbwRld2o0DJUb6r4rGemF5PWlsGEJyPw3
ftmKVTY108NU3oBA1+mD3/MPd+RYhL9jHM5hQZ+VILxIXl1axTwa0YK+pW7h1f4Pl2vXdFRQkyct
leSlXF6Vm7y9DQqdf56xoz1KZXTEOBmgxHCL5uR/Ua6bAWuafSmiKU2wS8/RlmsV/0Whk9qXXgKR
/g0t/guokX6F+jfBEn1xxcVqENXJF9Fq4hgVNXLVc6otKmh+PYfO/PKON8PPNrDZQm3Pckl34x9s
5jubWOiZ5O52rEQtSvo8jzosxyvtk674q0UyA7sKnw7xNcPIZ52JYvXeszxlpqR6Bxpb8syK4xhh
eXiYtQuIXzigq5sNGENKzK9/VpXSysmmARwRKxXk+/JINu4o9qN6BPaJX8G6lQEkCstw8XDObaFi
mxCLT4Dmv3ulynCrAphoz0t+Q20IQUjbRFAk4pWr/fNdMbzzj0Fjlc0a1X8tVFvuD5hRefjTE/4f
v1AY3YJCV4NI//M0wuTpM+q12zbtFD3WSBOx+lRMKVxSna4oUEtJtGOdkZDh3IWBWG82GPY7v7pI
dlFGVRrN36+QnBrwsDmHHb152X0KYmkd5TJNhWv8zdrzFUGvqZFvCPT3/RjPVn+uESNTgJZWA95r
Z4oGTtVX1BUIHuOzbRQR9e65S4wseCYqEeo6Qa71OVfkir9Uz+AUdZ7EYy2kR+RCJyi8hZ8E1BYw
2kZemeknJpJQN2NooByVUuAX6Cb2t1QwGJXFrfQcQbbw2KjWJA6e/P0keOJFGT/eogUsNXHzG3iV
eRfTVMMa0G6hCtEixep0E8NWeEFgx5pZzV/0VDF2WAxuqG2D4Y/XG/u2RweZ3KV3nO1L7uL9ssIL
VqWebLQN00KcrVa5vft8SE/wZV9z/aJIVCDfa2bUtA4R5BNaWVwMouzcmwqwdJYcX2pMqejZ7lUT
9snPFJhU3VNElMIz0DqVcsLHNqYO9Rk6qpaWeGcHHFTOp8n+6F7rFLN4zZMVidOR/MhJ19YUoIZo
j5KiHkZv+m8VCJCqurrwsAFGb2HAR/vtyQKDVvvMZBa1+I1yNk6OfZB6cyManmRszqqwJpe9lxE6
d87dIZ9pQZiOkwD2o3qR30ETjihvhWqtJQ4Pb5zsFQuR7jLS9twQBaWeIhFxfNRhbjjogf6WNmJi
3f68xWKFkmgUdk05ZVemgiDcwJvSwF+etm+c2V4rpKV+lvApYbtlQyb+L0roY8AHfJvshZBnKJTM
PjtXwOKVviuAutd0QKd5uyfsRvn/MKWy0iTrYHlECwdze+PRxMKaJmolJHVCfu05N8NOVBdOQMQH
3LFEoayMj4E28ET5iJ24/GdbAOnQ4lTjdaHtXjmYFykNTIn3W5uI4be6Plvp8YHrZ68bVMbt9gyO
zuidv+qA79RIT5iOuSouFQb+xsLwwfqoRJwVDdolsD6wDeDQO0L8EdTuRmSXOB/LLKYq3pe5cZdY
33TN0HUR5FHNS7SIFoGWYcg1AkgIqw+RHoaewwqmc+hIdDYVLJOmGIjE/G0HQFuiVTTWKhYDsrcX
cj5Ttp/Av9lqB0XN8dzDLxSuwQ1xE+1Q79I2Z5hfftKblnBFdOTyH7EOwSBmzni/DzRg+y7AskKx
ZT7CTfY4mhodYv9ohVNJDtxck19Xv1yjOWgWrDWn5ilGzsD0O6XE29TdP6Kt/DdiMO4NhxK6uQLX
pzbp+bNKCyX9MBzFhKVUVljybnNs2crb6bJREW2yp56+oRKerqpWMle4fuuRk1lBrK6bZUW6+Iii
s66DMb8FfZYM7hhHHOC5NlMxI4mNLNEPBOjHWmdDXKYnlL+J1/rbPSKoK4X+VQe3MWkIWXOxiGPi
++m0S3IonTPiyMdZzgVlqr2mI2FliMkCwBwGOYc9aeYjeztTWB0FpYnj6ZKkHZw+mNqtjUyV2vOZ
IwU4uBJT7j1K4psZVPQk7X6wXkurQ6YAEo6LbY/o1XS8jlmWVFflou2vM9rD1TmQTTkZijQ4FlvX
0x9yr6ZNpl190rjZMm1gIStWD6QdkUEXOneAxM1kwK+ZhKPPWpHKXHNtIstrmqgJIsHfH7r522zi
WpqnUmkckU3KQyfFu/ERgYrp0n/B7BELqLPOUbMA8ZG2kprUtsN6Yt9qvn8ww9v7+cwCJdNLq4Ey
cBkH3W9uchSUyd385eiVQilswXo7sGqXsj9ya/yjz32Alz8GViMSjLavJXZPUs1Rm8p8JXQttxfj
JfXHoO40/TOFy+EIDd20j8vykyvYJa30mf7SaOj0r4x/1kCD/gWYUgCc/hrhQqjWydiQbQ2Tj0/Q
HPB+rpT8tLheW9oVJi540nvqTwybW2THO/WkqpW0Q5onm4jKnsTb72/ucRiAs2gvk4Ah6IyKlkqa
51xjStFglkImTvAa58SarTuFztF03+ALzhv5Mp1rpwCw+JYOA+WhJiO1jwFTtY/JyYVJA1e6GqZb
mQ/6xdCZphMX7Yw2F/tX4JuFOpB/Eq0BbkpIFAeiHY7GjFLS668K3vVoe0UGkwvdOGcs2MXsfr5y
ktI1deWv8V4ufiU7iR2snnCsCZ3ceeg9gll3YHo9iRXtVGX+4gL/Yl2SPgWox1AsYrrmcTA7ggRk
Qjty7pJyQLoa3fKae4g9u/pOy2y8w3PQKlpxT+83RbBohAtnmUjaIzdWc7oeVJU8wF5maqfCdnjV
PeHwqRbQjdo6NGG/D6c3Pn95diRlKjwNWMdcOeGWaDuD7A206yjnCUXcm1Kg/rCosZoCc+V7letq
4B8kDcsjug8mAoRf8pMaZbFhOZPnZjq7VPBQSyUTMX6VvJkJOP5LacgFR+45YnT9wxC8FheHbwkR
KRpnqC1PIq8dLsTPjVDBvNLzoMjpTZQXkAXJqY+XfUxLfdJeZkOjl6ftGQsonPUTELPRBmHgR2KT
KO/OfXq8PEplNWnVVU5b+9aXa7/AOYKa6Jq9pdtYWYYTKLsUIzFXq2VkUM6YWhRehDHstKnVRREG
45w0z0zOf6La1EE8XWPTy6Sxe5g8KhchDelsu5FDU9cVGgvjO0mJIv1n50pSdGPEI53gG4JI53OL
kjZdw7CTYt8ZwGnaMX86gBvqBJQGKe3gk+I1eoHN1bL+fCdzbQ+BEFxAhviA3oqFgA47rBBhvPej
C+t5KuKJ1Fqq2mfGNk9ObX3UTF7J/NzujVPkqAVP33dV2EwJW+SQTwcbOOFf3TnDVigWKrYhASvR
NKFEAAdURNFAhD8gD2Nkms3moDwH+LyyFFDVmH0h4K604bpid/ABriLStvhcoTIEc6E6T3wJqXuR
a0K956yAXOLE7DzFLaAa98H4WHL7dZLrFccmG9vYIUb8ouhGddkIQ8BLqVz869JBEmUfwSLloDgs
wssjUqj7gcPLMfwqRhou0HGiOSHiFwQjo4ywhp8A1K6xwe08cpOqYdiIw9XeT7ilqoJCBUrFWqhE
M2nepV60QyGGPHErZ/Eqt5FbtBRnuz/HYMkLsFU+RIQ58irNMJdzw3qjL1OBZVnfKE1pLYH86QmK
DgGFSBlLGhKKbmYeCjf8rx+r5E+sJgpR6nH7xhAVwvcxBibcfLZ/hQStxLWfxzfc8BeMcjdJMetf
LFNl+D8wIcdD3F9xaBsExF1xixZxKWujyIFj6moPDt7NrtvaR+Mc/2B87/Bjmd7EYskxo+WPaHf9
kD1cnnHuQwDpTyA6oIvnaxsvt79JjVuLSflKetjDluK21cPFM8rulnmOkL+riofGAcgVyavsf3MX
ETakihH1CO2cyimP5VFK2WU9FrXmI402YHAQ1JtcOpfe6MEvFFq7y/HVDUol6gWvOJP9Uddc9MxB
tET7nDu+RHFBf/lGd4JWD+2/exZuLInkyfYVN/lPu/SIGufcDx6TTtuj6VFx3BFskWTtGCnu1Fgg
YqURqFmJQcoOoS1+4s0WRQAXajJXegOHLX8aDP5FpFI5FaIhdIqpwXUNWdGrVlKy5CiwhcMckfcQ
ILVwFAT8zip9zVnfh8Dqf+lJFzu8G4cgSMlcH2vduOyhKAfPLZF0P0GvGTyz3qGVJMSR1zs3K/qg
A/BfKr4ol9Hg7u3xJGqa/nJ6sqj1DW9CeIvnjlHw4iXn1juBR4Q/Sq4yqT5dFirZsHhDHBZ1A5SO
0bT8Cd39Smq3hXPDBoMCOzlMEHtlCbI+lx7Do/YlsRcJdJiogO+LX5hkE8lUYaRNRhOT5liA7M8m
kvsD8W5tLxw4R2IsMuzlJ07Xb9Z3n64ZV8VYyr1fHjwXrt7maIqT7fKPmWO8cWd9uV06KNtDmmYE
LMy0yqmezzvks5Ql481lf/UVrh21fOI1D92/Q3WQbyR3Ony3M/ftHhBEXefqsfLFKG+q6P8Q7Vls
fztYQdMqfvWsz2caloyN36v2I5olkG96QzThaTIVXg34WD0K07qJhkO+IAJB2Q2UI2sCwzivqGTq
MEBiBtH8Gmh8pROQ3GaWAiMC1BHRv9f1aMfDoOYad5wzFjEiLOwnUntcEO4CkdxJz7dPAnea2d5Q
bKUNNODhmc7tNCr7Bra0+i8B2oMTQbBK9aHtb+RkgttrvgaGX23hCLw9FTb2xnZao2crGVpw1P+B
wPgAXQMsMsbHDN5zPkrV9HAE/F36OIwsze6lYDmrWM3QgvZSdGqiQQVr1zF00D80WG18425MFY28
WooJiJvLlCZhWS3qZ9n2zBy/TwPXJcY5I+ka9E777k9G4RZVIKQcOgyqPALhKJpdQAL0KwQM2ZsZ
fsE6Byrrf7nbm5dN2wfNkC3w/QCnW/lsoT6jxwTl4kG4N6cKDBDZXGgu54CXWIgztQvuPdEBTy0y
aJDpzKcR56u+Nm+UyZiSVXP4/+OebQBlPUIUmPqH8V2mW1zwbbNi+Akgn+zzkRfzP9A8RJCcQ5RX
HnZqbGpMmHnyqwKO4mkGRjwB8x/mPHUH/wUF8krL/qHEdXjc/yv86afAJPgAYsQOHXFCL/RURQz0
ITUCh8dLvv50jMBviJfOLpiHWGpybRkabi7zHpcqfBMrFUCECGDT3BdyRbFXrQoerBzUBk5UbF5W
fTvhK/jWt8JxOY5Q6lgS3MSCmu3+b8XxWlBYDbjqJQBx5p7DmLTBxPmDIv6ljcZ7URkyJlyk2OqB
YL7s5MxFbJshjAjW0DdH32N8YKW1PHRRIm3FiZ8Oy9sVw3+deA5Dvsyu7OiPFSNCLpW6j4+4NsEL
ys/tFfv4rKl2xhad5oAvuHvuLuRy8N3AdtX9GxkQhmdUoprUSZEizKRl0/KXs/SykeviAEIuY/XF
s9u5ZSv+2pwOMG/32sWj+938m5IV2vk9G/d6HeEn+MKqBs8bNj/KkTa2BeyliDDtn3uRjsKdtCsW
P19tavCYiL3PELVTYINnpGAXe8Zz6ld/cr7xgbwan2aln/8mG0MQQdD+qXiAQoWlD8aQmFSrZ0Bq
vNDBT7HWotnnVIsAF8eoJn9+Rf0+j+n0D9wVYy1ASBrzcxy1UVSrMCeg4AeaiytqLha3RP3UjSTJ
W/rzlyLwj37AJC2fVIVCByuF8oLEukqOaFTQ4tc+nhl/nMizjOxzjoVJ54UL2y0kJycW9a9mH8BX
fvq0/ee9383C5ExMd1o3uuUQ9jYd01eFf6XOHNzI3DU6xp6ZZrbdH19HEf2Rj8F5B+5QOwRfRLkM
7ksnNGiqEHsiAjNDxGOjY2/Rj2Kqyl0loMcp3+8I1uVoNy5fQaZa9XsXnjd39Z0AFa59kl9IG9da
a7K7C9RhA8t4vTJaoIW5CuVrwDUtDhJIyIcMguUhVP46fvbhDYZ6KJxS1xHbQ0qoh65c8abv05lE
ozEr7rei2OJMbsf75nZqkIvLEM2c1z7phxhM/D9XTmbwGvTXgpNakgk+sVfViAsqfFfBKQscYypL
6XqDju3roTUlRkgJ12FmlPPrK164sPsO2u26MMwLX6Lu3VKrgAN8J2X6gyikCxItzygsjG8a7KsR
I7BUed9ofn+7dSBScdds6789180c5McpCXiYP6vMCJqOv/wnqNIyRNRHeR0dW3pDAudeUaQo3cuA
XOpicRyPzZfYMIfKb2AFOcQuLeU2PL4rg/wVyNkL68Pj6CrKFQCeSalr7l/ZMDcQBvhND1i0Z3yX
xdsGYBYnM1eVELPnxeXJxK85sUB35D59qEh4jD7DUdCE2JRM6zHvmzbjHTm+a+zBrQGcPz/M8sY5
NV8hHwoXX5lp9Idc0MBOFqWrOhNzWi+5HUR2BQXMW5UJCtlLHUdNqdLQBTAyVNf/kJJduoGA//1H
LyqZeg1kh6CWv8E+9WqK4rjL6tEhbo68KSOfLGU5kZwCCD+zVRdQ+mQOQawVYzgR2dnX0tlcY8Xs
2Fgr/cV9reFGDbulltQ6uM2VbWuTgKPI05RRIUoqUJSNBv/gxIrTdK3R8+dTy0uHEooQJeSbIRFj
eBqrFtX2naUXK4eefcxuoirHDEJe9F36t1itfO3YoWmKZEaptfkjV3QYDeFzNXR9T1M+jGSOOeA/
SkoeBXNna/ocLvo2rOuwW/sf0GYbh7KUpprGQ9hgr10x/6kV7G6Gb98fD6HgHsA+BgXKXy3j1SkC
mdV3ljl/QhUboxhwU9uPTuXLzJiK8OIViMrhIE+GZ4BWeX9pYQLRd2hi398W5BRz4eXndvjd8wDB
Kho4mACwrqKRtTl0LrQji5Lt7rEL54zNdXx6bFPEZvU0Pwxa/tnjaBssDmT1mGBQilWqYJnTwgks
CcG4L0pxXvXK25mt/uWza6U8jCciU5WrhF0Xb3I20C2S/mVQCkbfEhR6lInLhj5Ch3tFWV7KSaxb
6xWxQyE1MhHXHgLoJbsXP61s3vpWeoU8x6thjLIdeqb/6UzNBTp7dKdrGUO2TcUo73Z1/YOvBet3
fXfZUE5giXbfDhm18+6avZwbZQmwKv80c+9wVfsWngeQRbYf3Sel6t+PNPxI00ZBszY8s3bODDuG
OKthc5bfVkj419mbAnNt/BhmOKXapCtqBcUTSjAUIJH4XmMhVYZVdyovFJ7VXRumqOu1767KAL/X
UynMSQL+CCCDv2S+ygGSMUkrnJHyz+tzNItxWPWJDb1TRmqMkjpk6UIqB2nx662XdUxBpz47xC8B
emoy4MxJ3J0bnRBAFyZGwuqiuXCq1TQSrUzSJm6YhjezRZ25UqHM5IPC6CU39TOt8exuUO3wUrSH
VFPxa+p7NmGJaC4pAZER+bnld+ue9dZ2pSSFgXlmvmf8sU4vBpZC+SXnINhQFHseKHDpR/Ia9Rvc
6guVdO3DJOy7WssiLvzn833jIXPQdhsRs3QdRqKN9CrftVy5giCH4kYPSiucbWBML19dDJGvfxjs
F0FAEsv3GMS64bNKvOzZDyrE3ymOl1vsejKpJCP8wYiq9BExljwyjhlRx8qbAYrONe1S6YNL5Q8A
8W88QNhJ0I6MWfvxluAwUEWdCvA2fHX/cMy6Dy/uqY2r2O1fWeu7mcKCChZEKQER8wKnCjZZLHxW
NqV9E8vJChhByWRBdNhBsl7T4b0TOYb/IxzQr5PErTLQGQwHS0oGFJ0om/WXaI5q6NI+KmzjnODw
W2cF4KQj+pZ14hlTmPGraJhPk23w1oi0OKadry68abSLOOXpt3ajYV4ZbmcODK/vfsHg1+Ljyyzz
CNP4yIP3bRny9FUBXJ/A+Pm/oaMzuxWRDsTMDFaoidDjvLkeisa8uuXXeCFI+MYVDyJOCVjL5veE
RlA0qYNZDGbQkNZjhG2sj+A2OBEVYvF1VOBTKt8uCmzgOd6cNfofRFJCW/uGHjjl0VGwb/MaxJtF
YWsw2VOl3Dc35rQlKNa91/1Bd23fFxTP5g9zq1OgvqAkt3MUhRIU1bPKQjrXz6zV8z2jes51I6cT
a0zb/X07MkfnBw70WokBgBXfAS3xaSBkpFQvXVnoQXr7Y8emLNvdjy1bwuvpOlex1YtL1LzjPvq+
iOZSPefuLva07sAAnzkan6QhSrFXlA5g2h+uhSN+0amtw4l4EQ3Ckcg41EpVEh1qHVsrmAO1rtT2
uRnQM37aI19sqrHnM6Aj2QCx6lFROvWYAgZ6Pa0GRZem7FMCQh+Rv4f6aBjOchqAi3x7fqvb004i
YQK8eBx/JZa9/yHkobgpTSqHlirIvZ3FS8HVsio6CyoYBIYxC/ehqYuScgKZr4+q6O2ydJuFLfAR
78XqxJKQYFNTXakXeIljhfxmudZH9kS8QSEdDAQXpYuRn9N7pXF7pBbWX7kgCHe5A+d8uX1pfq9C
iki07AgnioU7lZo/BWoUQRM2xLL23/3AH4DbItLZH8PyLwbu5G2pacVFC4/xddubyJel76rVuQOv
Q74EBewr8SpkGmvYa+zpKIKIe7Z1dvw2hmn+I39T3ieyaIrCREjmSdQJi2lLL3JJoHemxzF3XZ/s
GXNCyo30tmMuTIhBZZg8CFgrTuLOtJoqrLjFafzSbHSUkNk/nztriNv6k29BKqtKytkj6uw0McBF
SgPa2R2GSyR6AtbW3c9OTAXdhcZBUlWcL5Il1d/++5QTzc4Gx3Vy35VvWlDPd9MJyCCj41MF77ES
AQ8raVZQjaOiIK6slChTVTvWquJTy8EvXnt78lWbYKoz1GYWadR5MMSH/4IAAdcCAc1qoIzGMzyh
0VMIVAokNKjiWkXMZ89O5zFFCnD9h3YRkvSFV8oDmOaq+fPEuscTDyvIa/Xt4q/tJFEd7vgT2hMa
pInPCm11mwN+BxvWglwr7G+bjfe0j9hZ+DQk1RFB/i+tdKIoZxkbgBHNEYxrWuLZGTKWhyelTDJ7
1j2v7Xo0ysmr6A9DL6KfLWTA4T9RBJdtX8Jkeb2mlS9CDJRPxi4NtYQ5lqA5uMbR/c4dFk8ufomc
6FMQyUhxyZo9B4pFf/6wbVrZSCLlO50unbW82Y37cAEIRkNjao2t14Xv/hnw1seYW5FAesTFiwpU
a9vonZzzuOoKhKq7LYpYsotKvLntmoHaICbQSYb/v6i/j4A8sunsX72bFLjZm1lSi0iG6a/v/nuR
R43qqaxKT7UvkRyTxxInoCULZbr9NPkkhhJBm32937Y+5ktwTzms5pRZaJW/IFHSVSV1JaJfH316
jbvKpqUxR7UXdtwmyObAwekP3GtlTFF1mhC/i85pykS4V7qAm9BO064zanRYo0hy6on70Fx6bXBn
2LfMt2S3Y1FgK3sREBYwsqrrdV66GCO5WjI7lI4aav58mwssh08l6VR9HdixLubOddvEr1usR3PU
VDz6bGARl9wV1SjKwgFXctDoRsI39lviIy+j1c9bFn0ku3IAJWTFIQm1G5Ec5MWlFaifAoUFyg3I
bfNwLvvB6r6Zv7iZijUaEWMOae380X2SYwEnqaZLW9Mb6rv6iQt6CAhczHe6hsEfvpxpwl1uG3SL
9miAUHwK7S0XcZo/VNn7OGjoDzUlAigTNkxhhNIedd/SultzIpTbYNf5kaiG55L6kulye2bFB83B
2BGnOdleYz1dByJUxzqGaTBrhqsHBspzzu+Jks4SH+ILIy9e3kA8oY0NzqOch03wJ1Xt9tQgYapK
X4aQROfOA+a0epe74fYQV8uANdo2Car0ezXf8G4nZu4S2TPSEtsF0TlIU9QTtK9IYYSNx4FOAeSr
fRq0wkz2GUnsX8JITSTUB0UFhDGp9WLrLDjU8rTa5KqxR7rwgPHqvn3mSTPsbXmCmbQsEsK7iXZR
d/Hus9X0g+JxKfXzZoC8wjLMD/QFYTb44ZCjwOgCUGUw0x4J+HxalKfWCNUh6qUfUy20wPMLr8YT
2gwhaJwnfvKpdOTkk367p+r/wNZrSuMIprdZKrDLwkfXgfWkepNHVmywB8VSoHMP+AL45sPzMGyu
oCGo1G01PfJCDh1eIEDdJxJTi/CDl/j9SezFwvhL/Gt5KCjlyriNSmJfz8cpv4zRUEiq5tZh8P6o
2RuKRZ9ASMPbr2H26GU+8WPQmD5MX7NI4A0cZmgSWelNAd+1fugRcjxsVJmvchGFBFQg84UXpTVk
DlnLoX0/GwtcPpxq/r6FGqPIpd5ZKeFlPCgXFLviAWJnPce52nje0XGhXwyAVAUqftU4dkIUwmTY
pDreW5yUWhMlPEcjlUYwHdYCjOl1tg4Aze6tAf574uYTUwxg4Nyv/qAv8qwqn6KAYmnXjaPvbBW/
fnBZ5LdZYvnw77qwAoj3U6HPyw6UMCLTcCRse/v7DsOZiCb6XXeYBU57NQD+pBr6Jg+OGvVANyPk
P2OIsN2Q8tnujmhzRUWnE87xgGzyiM0JG/nFBv6cdYCIOVKrMt490sNskPBrCsuflBKuMkJ88wDU
HbMZVaLzvpxVC4+n5hV45+mVb4f05MUUkHoiIFepPxoB8fBq5RLDykXO9P+hxriWUZfYmGQ3+yFK
vcduf3YqYpl+RMvA7KpGVnZ57G822EUhDubeJ289k1Zibvz+PXnlyEQw6De/dpnN+kC4ImEnqd84
9xKo7z92DtXfofeap2LuNLgso6afKYFcrEhYU3wHz4AoJTqavD6YuHwYWyoAEkFcq5VfKNrqxpri
4xYvQwaBugF59cMXucFpdAc8hkQ7UBYZti7ceHuDM+AgKa/IwlvoV9Tisz/khtQsB56zWfO71HKK
xSgCNl4Uh6vSex1ZFNTqrqCFkKTl9eDFTqXKOIsFFUnZm1wVlEBRh8kzHeE3A5k4FTpHDFPzjFU7
frg2i6M/pNR/m5APAZTcAeaqlizt7uTsMLk0FO4zDVFNhtw/VueoVLDDVhAP41Sj7YsCI2YCC+2N
3HesXlLTQ5I/iLc60ovCdpMOwrb0rn3rMrOVaoIgt1Fgxv/UWD8Ik89GkwpQVRuPzRXrIYg5k3yA
x9bZPRl5tXWNp1Wfkyv7EmOvgIeJ5+BrLMDZspnI8bKHamc+3+6z6stQanaSZq1BHIMhE2dQyRus
NSTQ+P++lIq5f5gLsl0xlLDSMACAhO7/NWJe4BU4KlGT12p2fb01IWDNVry2g3LyvgsVnjWwHNF3
LbfOf23SVdF449jcrQjGfiLJE2xHDOw6/pFgHuRiFrSOa+d6tn4jOjRwct2sEHvWjT6Lil+RipnC
TpsIzOm48dMPIIoKpxfVa9wZDmrCquiGnEUYZor+/b1oBxu0qfLHILXutiFCL6+EyngICSDsWg36
8uN+LCxYmPtbvTB1A0ly7grZU5w9Bymck5ueWu68Crv4bbOOnKfDTBQgjQf5UTigIrr0pZYwhiwG
k5HCw2nYwRuRm6BUCw+kEpGokrfsvWxuc3r+Ece/sLTcQI0AvRRVbahF0Mhan9SXOTLR+Xh3b9oI
m/qUh2KqpQFVZhRN1dQEa9R9n/4C7PbTzpPhxEodw284ih/Wk0I0aTUVwiirckHtolHccML3vUYN
8ZGKKEC8ef+0hprD1VsVvf8M+Zrt2wITC3C1uUEYx4EJYdAcpVF4aDnBDb4cFDCCwVGPWC5R0w0B
QZri9rCh3/3vm4wGywnbrhPczifK4ervA7SbTiAMtZpSzgqs7f72tBZ2M2Vhf/Nszv7ctagEijho
7Ayw9c9abOOoW3O29oowTZLk2ofPt0SKJPvVCofOuIFply2yUZQHYLysONut4S6CnZu9gd7E+l7h
d3CMaH7dieK7b9Ezu97ceSVK6F6idbdegDG+k0ls/v94AAH6eunm8fiOadYHQFEsBz3p82rqqpSl
MSiY9KUm1634v3/62SJo6MytMBGNiNd01O649UKeM7Xl8sO8I8OnYfcSh/8QcHmXUkOUY2XC0MCl
M6TZplPrwN4fq7oaAB71l9lc9hjiuTdH3qfbLSFz0ta0MBrJERZ1mUN/ocWqJ74i5GH9ZbTk6emf
mXQF0iz+RrI5dsOlI/EmwyzTpTLu/rVXkjq0lG6QlbcstxcoDrTwOJ6Zaahb5WCRxVYnF02TKHpB
wJesaoUcwEXFVSimIV8pZ0miG1GoB6f5SnqLqnMCZHxAr3XQ+/Q/LGnGE7hCwZQX3xqyPyl5IWfc
+9EAQUyWj3+DEXUlpqaT6cI6y8vX3h31SZbMkxBn5NYXNrPhQbkj0Nm6dpm489C0j/SLTbjjiGdp
R9C9rnOnR+hJ215LpHEjTJwAHYNbEBOdJSnYxu/hfqO3kqXcCTUD+DwX84Y9hZvkNokx4UF66Fzu
SqoPfquU11rt8TNwQ97TLfCoG8lsp2bmDtWS5QI4X2Sg/xcRL38OIKDo7JlTOf7lgQLI3u53fpPx
dKUAV1m9uV8C9PcWo2CvbtTIvyYmk6/dKAaMAY34+ZjVhOPpesiEg5HptQYkVOtajvV34nuaVg8q
vXCr1luEf6+vOWJNogMSnxnZGRr6bAuklrzZQUNWz9j+wmhpNcCsBLeAjuTd+nps8f2oDU5ejaYW
twOb0bw1ZJD1h43wgxE9iTEh51DxR8t6yrbuLAgBN96aaDwaqOTAlRArO+EiSjAcQDG4Z0MJcFl6
hHaOmlmHKaZ7DhJIhnp1m5Dsu5YePiTpjnkcd0nENf7tN2neMws+0hiUrU9pZmAVZICe7VpVNzpX
R0f2uC4pgQey2y0OiCCaXFaD1bU+uHQqSxVsMQ87+WtQ+UEUyCDHpkjaWi8FKIxRi+999XBIIPkT
rPYhV2dPjoyaIzTwOoXQrhAzLbNjnYLmR0zErzE1NuYHKWF/5s10EdMqG6Uadp7RTEgs6WhosFvA
KTHhx3aGLHqsXqXt0vHIUBDHlcDB6GzRNWpzxNoLogC+zKwMc1pScacS2pMuw7DFQ1aS9x+KVYwR
pMbceq/xHyGZgUmqsdAgGyqf3pZNd/AUSUWHpU83c3I4E7ngVUmhT1iNmxeCWrGMOioVD7bSbZpR
4c6ZWHnA2ozwqrF3TfRswhRh5jNvaUkbepjpMUzhyG1S3pLKSRjuaGlAwo44pcQSWW/vptPNVnBV
UnXBwRCSdki915E7YKJuKOxJg3CUiTu0kb+0coXBTdnNuvkbygpQYabcqdOPPJqW01ht2RKErNEx
tVSQGGYdwBVOeoICl0ZFVnQ6mnAWB2MF1rnNfDLLdsHxwqEMito6Uxy1Ydp+Tbf8LAP4Z2x3Lf9D
203FuGEwv05RTG4AlUT1nEThzuhuBqbhDm3/ctbgbpWVpm7EgyDhklRlv07bKYjz7QE3grAjFtqQ
KVCwMJzlAawoauZl7TXSdZxiz7aceXhC05jAM46AdezbpdAo6d5wsyalZe8WQexf88KcFSNEtX1F
APoRTQIQSlX6VI1crYDqwOndV8Nw0F/LXaDUtcP3EeN4JdmYPZsuy5fmI+ZZmz0Wil4EdRbp+CTc
EFLs8MSGX736/ptqmbs+ObN0XlV5V1onwqi3qo0LMY855J37OI+8YsDGcf4BzmH7ltTSX20W2Jlk
FFhWcvspvizuQygsc/5JdcIQE2ncECOdG/cS7j56xqTZeFuJP0r41ZkJ4FlLT888wHw54FLJt8BM
7AjA2r5J3iYJ/f4hQIwKWuWX9gSoJHyrs/Bv9NiE3QetyixqPGpNFCqsxVrobm7pMMy6mWsMZBbw
sEEUX7zZxoWQBTUbe8Vug/nxb6rvLOLdky6RbCYwY1JG8ZPCf8hJ0rh20j1JVBGcndev9TWoFNfB
rxlAgObIsiLghwu4hr4pyK1nKVKAWtJfvrqeOCGcCNTjfG3YpcIMQdvvCv7kwYvwwnzePyTNkhLm
QY9bAxb/qUf6PFGLOEXFOwh3A4LiIJzygzjjAvdK4LDHo5Wbobe0vxHN/p4VQYqZy3soHmGVlsg6
mZTG9QG9L80DcZ9EQfi2RHJsg+veql3DutQtBKVVKhBaRTd2iwcAZYjCcs4e3IRFHlrDYuGQGI1F
Eqs/F18554qVxtXLj2mH8ybOofNlr4+0HrO//aqghfAcw5QNMyoczWktEOCGPk4dOokHMiZ8ukru
Z+w6aWUmNFHqczi6ejeGy3aF8HFtymMHYasEUFqKvnpstGpMNf8SPZKbHKn5r5HOkKq0fKeZrPwK
AAlx4Lmxto+IVThOyFdImRQpwNrSabPo8Snk4ZOSoH3pR7DGLkwGaSvDOduTsUQVpIBP4r0Ax5h2
byWYC7nAZO0/WNiaJqo3QBb/Omazr05CxF/BIwCOPWuBlPApg8r8cyUkqUTBDxEm6OiZYuIWyMbl
z8IThcOR4uKlmALgkQ527lCJqjmb1kVhE4O6Z2FXJxXjlEd0fsREyv7iUGl9C5H2AI43RB3hHhvx
QoV9bdCgiTvQns5Yxp8Nf/LnyuoMAu1bXJr/4JtmteUBfDJc4JIKyIbq9w6+JaKCiZw8BS9CeVq0
H9GooVBF8QkpiusJfKSmTbhJOZSu/vG/2Qqi0XxY+ZMlN7vgkNKW9G/gnOrcHoBIUZDFHa2r9g62
qT+B9XIRr6Cvfuwg2khtrPZx01z88NHJUp4MYAI3R2Z94k+b7E9Mt85T0Yt7a+XRbix5l5Ero/1P
RBYxyBMLPkBpDeTpE634XIvtXnk6yOibJ/YJEIQ1mupOC292BD4AfKzb0EL1BZNttXC2xtUkrfwO
NxXXbxla4FzeBsx8DQFvBOJb2sQaO2vQ9Nyri4bdyH7ntzQOCOR0QIBQeLI/Ys0lrCTEukzcdWW6
fRmkNXvvDW0ZcB8hSVy5wMP3K9hV3A9BZKg/gaSFDFk5QVbrqdB4lzl+fYJ7rwuhLT4GAo3SGFHv
ZA5Ee42z+A8vjxRelea78rocBR5mTsRK9WdzLgi7AVHF6E6gZnnm1pVxu+TaO9/bl/ievcxZrxty
DCikM+WYWOucG+1H8s18Hz+RlwgnkxrYDXEVbjxLemRkWGAWCGhUPwTJgZV+ihqE3Fn9ljj5cZfn
6FdAwzLy9rlsPboccuAma33jrIy8iuURjql40+LCnGZRd2jDr1NaBj2t6/lC8v9ey7kal8lZoqKA
EerZPloMLY2890b3mG1jgoNQQFMn4+Hh/eR25nyLnsBEX0/UTaFCNTIeebfu19NFQyRt26kzeJAY
+hcKAxuvUfV/TmJQw+sP+sTFV9MRK7h6VeQngmc+xjpJhbEyJd6feeGm1drySJnW+jBUhi53A1PR
Wzr91bHTMLZ4nr35dVtRgyJ8osez5Bbwx+qdnwcU9LsAvbCjNZDcu+nYOJ/KRFf5TRXqdHbcPkdk
cCTudKOIEtyOKh4QUB7RdsPvB2KiYoF5oUCYkx/ex1ZXMMyNdTljN0XYGs/LGNKXzKphrZ70wHuZ
WPR+shICVODTe1h94RD5IrxE0ocY5e6Sd2JzPmpENPKD8bR1msCk4c8gSH//Es3tXZ+XGTQvWsAO
slHH7Mvb2T5J3i4finMT2LMPNEsJ+5Pcp++CIEQEDF/Cdh740p8h8Nmk7LmHzmlLZpvmDiH+Qf6f
DtrdB6fuWxOUwAs3jrfQjTVJ+5qMHjEu5C8ei9FImXlFvlew8APDzjPViV9jm1kk1DT3cjPGE9j5
lbQa8uPRrq0qGEsn2Nsn6kNbFSb8bUMLifTogr988YTNnzc1kv++r8JSdMMUJfsFNGvpEggcpLfy
5OBf5HPvSC7BTxnqPm1Km9grWo4zQlPmAhfsN/SMyC4WUtE4ijB42PuAWXQbUeX41tWb5RZUAQ2E
yR+1qSUM9OLiYB6Cn9ohTj2KKY8aI2EaxGjuXDSy4/VoUXuswq0/Siab6J+ui741DMqPoOvjN6hN
9zm2jz7MbqA4qMhrf+o2LWrAzvdjwDbqxjoCbLD3/colIIE8sTB23ouZP+KzVh+aiCeqO7nOqQm0
2IBCeBOPqICyUUVVniYL+p7/hiyWIgvKIZ3XDY5278P6ClZlf7kPJQWxSlB9k/7r8E83Xi4yTnmB
RRHQRWW1itWqqtziVnUgTHRRDazfb5i/IQJdPNAmizPRAuNgoxTNHXpAK55G0g+jEnCihIHX2Eby
fU2WG4B6WA9jQUatjdOtPvLVQyRbx8RoUVEYJXLs2KDKQIEAf9hbwhdV8YS+OX0twYpzhSNWnN5z
4kW/WBxNHuIyROM4QGLNoobFm08wq9XZfyHuaSx06Mz3CDY48lV3p9XY38zFLtZ4u6U2b+YSYmdt
z8xtJp2tFEFrwNGQfqFUksf9qE5sQiOli0U0rHajSuHbMaLxLnmH2YxcmUmCLO1h/pOOc0CJhrQ9
5REG+w+WjU72j4xx2XfV6/w1K/XVoFiz7wDV32J9ktio/bvjyykSzAclUIqWLUiSGZrMQTEvfcCP
Y/O/FgRmN1SHynKp6OkfUa64vHPHmsxF8Z2IOlNkY9gQQs5hfwFd7H0CDwCLGbRxF3d/HSBaeFGu
z7BZJ9aA/l15il6DxvIj3Jh4UiIuoGuiC9oU2lSbZbXvME8KqCeqtSEusAHaaBuyVaVDHlR0HnNk
h9DdxZEiDTJqPqVZzkw55MhqIclXgxky2h7SFEsEe1fxzpgxsLg6/3m9M7aAGX6+BowebxEbxnV4
lXdErraEruxICVgmyw50YrV+5DgaQ+nuZg6ADySFdsFA4Z3qCV9pPJkHErssXOdEsWB/+ATgJ++m
hhS5kcHbu5ij1rlNoGfLKuiteNsyZEvbt2eRma1ldYi1V2xjQy1wocUKc7h8JE+qcXXxO1s5vGaH
51TIGfndpS9bBgbi3erKSMUJRHWtRQtzhHveqcEuolsFKKj9Vt2ApSTQ+qF4al5qcGqW8f9PH9bD
DZC+vtRo/oKQYQmfjGqTmlLY7ifcQzNbxZS8JdPZ14pYimxI5hMvdlBBoZ4oa33oDEKw2/sQVJyo
BplUihyJtct1d+l9ACiIoXQFQm1D80VtVOUuE+acOJxfPJoTESs9JfSz3kvmyksCAWhDSaU30MyD
wtPuHOoUhcCSZxqlNjO+qfGindqhlAIZ5iFHmqp5u4aHTqi9k9PDcUO8hR14LJQ16D8M+g7Q7Spd
wgOrsMaqM8O4rLEPvvjhrH1yjUDYhhXzm1+YPTEgp7a/42jxBW1D0g9iui+GptH/bzQvh0qsEroW
jHfy3BVNZY4Sb8QVFl8qrkY/2B+Sm/k0lyH9Pnvj36TTIsgNXhiJw1v7gPAGbyZINE7pTsF003TW
iqdF0DZexu0IK2U2zuUGxaKmZZAWVCYnvaeffciP4NqzpHdir+B2kyzek7JbfAdrPh6DUzUzg+kq
FBlVqD2f5GIoDCUaomor+fwUQlaSazGKrsCGTJCIKugWrCllyyBmXkhQ/dsbHTeHV02NZayP08X9
Ynw262vWcj1AO8iNIF3CMcP7v/qAxa8WzhsaQePLcLkOp5DBlJSf9woB+w+oz7vJH5MVgPkEmxQU
/HVhyVU90hucu7qqdSDMRgAZMF6i28e7qG5A/yg1LJvrO3+ODzg2I/pRAQoFdO8XQQKs7jYq/5Qh
G09pehUn7u7WLH7QF/AHRPn3ar8tRRdEePISFBLcaguwY6MRM7fbRYlxthbR2gsNqRHcItkzQukc
iyw8OyQaC8R92G475PoRupA3IH9vTMjn3lJzErLcIRslPc9XZeJ8zDbqOBf5mGXFwIaLog041KN4
b9Oengu1AkqcoYVd2BhAUx8TpVO5qDozbrqk3oxtbwZiJfTHncdP59GvX+et6WbTFS7f/Ysdh75a
EgyWcwPY5rBKuXi7noITni2cLp2jBVDze6wpdHnd46Tg9IMrubIjuDw9hjC7YfInlFWl0ixcT0/F
mVb6JK3UTH7055myZPkg1Qbtac0VPE31HI8/xOgag4Rc4iXibqnz/5Ulmw8P509ZzzNHvxSEVCta
ULKsho+6Zn4wLnUnsxwjTUdckZvO8TQ8wD1wuFwgwqjrYXKXO7eoAwROSeriV1mgNGD+UbP4vXLc
LQY6Lk7xXaaCfnCxa/MlpLcroaDl32d+7jrzYRVlAQDP1V7WE1sAdfVAZq8YH7D85KTwa2m+pzQv
DOrBeWMlN9yWptSdjrYzReNkS9fx0sLKk407EZDg/DeK0Eiqijj7E0YNrMndBI5Mm/pimu6x8s9Y
fgEPXl5q3MfxEgmkrBxXR97KG7loGRjeEspeJVn4QPHf0sduKGiA/U0KRwpcN9UdxX7YEdbZVl3I
Hkcx+ymdvWOJzqbhVXjjLVUuwwmruZLJDXcOXHyfLcm/ssICygmeScaiFfbb0aM6nuyM6JLYf+6G
6Op03JX1E4c9AWtL6ApnIhvtzhnelrIqhf1umA/wlhk4hQ3MzgK5ZjA5FYruwPCorr3f1ZHZ1PMb
l9Mq3JNtrrfaljbH3vjrqNrrDp37pYqdWNLoyiRWAf88NlkFPNqYJi8G7qDL3A2f0APSX5J7cMSG
zgEl2ZXUFwZ0stgT8zRd/tKV1X3Z7UEj27ChBITKNHr0ZZbZKVIIF6sVIvlq9iT+zNUD3YpUB1sm
vzT5bv1j8mjmsXY11VuQ1/Q+VdeEGA+OQzVjrNrUYfbLyd0SKvn0KxfiiSVgPNWxBoaDJSafJpsk
dDCwzlDesfbZfxaenCLiOQWVQkH3IVxiKRwMsxtUv7sCHjg507mmFo22EtSzsif83upgbBF9r6i1
Ot/IA+5JiHwvcLQugu0TN2RtYwNV1j5VG4MfQKKSopz+rW05Ug3VTGBIF823UoYzQoGzodTSsqMZ
oq8Nmm7bXzhlTKMRvDZQiqZhEX7ntOUUhLOQt/GjJKuipYNHaW5ngnTPnKoygYicsaEQiQBz7BYY
hldjl+pX9DGYxQw7hBDSu8M1j8lL9gLRsm0PhKO5OSXhUo3zMv9WZy5leqix7daEsMKLZhyqTwiQ
5p5M5u1FU4v3y4r0XWtXNmIAKY+s2vDjYBD7wUa51oP8TpKpldDLsQQNhP6Pt41HrZ5PWkx3pWy9
k1ApckfwkYFHG+CGdPbLEEwzNDYxwHE09pgQOoLIxduhjQoVhPb00QAKaUKLHnfDCjgwrEEWcp5a
WNlhX2DwHx/hNisfk5+SJ5kUqvtA1EmF+/ZH+WaCwIY57okbTisEADCGI/0N3VjC/b2fr1rKmd7D
DZ3aryhaiNTZ64yNNaODR7SUyHDAhV9184u5Bj6s4xZBAzSmOglrNfn7sksz7qDfQAVlKERU1Nry
kiNha8dOSXLfVhZquCeF5ybfSgYbQskIaGi/F7kr3i39aiF2iCRZ5hl7vHNcdy/nnGMFFyw0XAn9
KWdT2L/XXYXFyylt6+MgqOyyxrQRa2DOa9YV3WEcPgOEW1nZMyyAHem0RLeDEGdhVXW3Sbqynmv4
mesyaoz5gf8+Sm+6gGmqodUXYhQdFUz7l6pZ62IKtJFYsQe3L8KLd6qtEntPyX4syMgvs4XWoitV
BTeIP4bn5texZEORaEsaOOhQd7ALr7h77jI51TtlYqR9UfR+68tYAt0qnpsJNBiYr1Hrn3+pTTpr
ND0g4AUPiRKOgeDnb6CyY0xhtgpST+WhpS6zBDC0P5pbwPDSV6HPxrJ1HYvmYBRhQ/M4wZOTeChM
CuDskJXB3g1JFqkLUu1VkKa1pDne7sJGQNkRmMjtx8A0/5i3z1iXcsH6MHPD3orW6ZJfgh3xlko4
J1nIpTjWEewbLBCXh3THZie7F98irPkyBN9bLeNTOjDR4ZwSyTtqOi+JvahZ/mFrv0ergOpu5o10
uYG2UYVOFTQ2KLOvX/vVuEqy1a25PRo87V5/iclqKkFMQuZkJgNqzmIGc1oaFen+ZqABIiLKdNuf
0Kq7L/dmSU1+/2XJv5uKSBpVhlwXSHrdyOX/R6NeWddXFhGFr+//k/WucdpzqDMyyIxSpmFgpIJq
Kk1DtEEQQ19+V3PTrjLY6SWcGh8o/kbsj3MYpuoYLBXp2OroFUgkVLKoEUpJTiByYqnwdjGYdWuT
bWgr1F/B6RzTffXKjMPa3ddGA3X2oJ1LtCTtEMWcsMnCyXQyPEPS9HjihRGEza+Sjz5ayymRczsW
BuCcnEhScny27FC5rY8hDxrwSs3nmFtF16utHUO4oXigcNTk8gatvnFxdp2rCh88Msvp4aWLILaI
1lBaxXvsECz58E2DoZd+eDyyHhxP8PxIczjoocQnIUHugVdP6/tfumshGHoVvzYyUL6q78pLfMRw
JSZCQF3KNuEBa6GnMkvMPuMn9Kak46wEb/jEBycLWsENlOmJKyUjuumH9SNLG/sYldtZ00307I+T
ppYnlLjDbTEPBLxukKKwmR1R7d6x4sNMb+uaB1U+j0pfKWLQiX5Yz5iGvHdfgaV6BWz2Qgr6Ngrg
Oa1AAp0W48N/6nQXXZWfkyfHjWgTpbC7YWhFLFZFwH0sHU7Kow14o0k+PzSWC9O0Qld/NLW1jToC
spSeIOjq8RHhb9HQ2+kb/cKS4QGl/V6z9iuqZ4T7Lpbq9Ub/8ZO8741bz+EjiHeHxwqBqScqdFmX
5jZ6IIL3q5OZq8PLg/xo++6VUTb+7slbgAYPWJrFlqO7Atw7i/t59BnVfMoFd1ZaQxRHDK078Pjw
10bxbVMpDd/RMO5zuS0p7kkjntPJkHK+hHviYesfSSfhh6qGcDy/nE6nSgvfvUm337B4lPCtId3B
yrVjiZMWtZxyFdosDrZVjFnCQkoavwBiQf2Si1ESR+Duvr/NuNpfV+Ztb4gwk498EHmoRlWpViSM
gOhWLzo7hMRHlMA1Kpj4FXdwfixduvN72SmsxQe48uOW43Uh5Rx5KqghkgH3K5Uh+Db4JJIkF5Jo
GELwdXOsHlbr2s/zTJ25Ml36cmeHPA2qrEfsl/67ApPV8n8enU4XeltrRVvmht/jo7UZwsgF609Y
7G0zMOZAChsjgGLh3RgVSl1EsbMae+KerY3PKgCXByWXplqoQ+kC5NhmQVtVyC/vUtss8E9vPa10
Fys0fEP+bzuPHzl0v5bmfAHl5oE675htqcmU+ZAw5kR6s+iSjsXiRv3hLuipWEVqg/OYO1CaqVSq
8mzxAMdJNZ00om1+RM/NH/iTkuEzdpSCilHeQfWw83Nn/oZBGRyNplpK0PoNOUOJr+6GHVJExgeB
/561m9dwvmKnvYZ7D40M9HeMJ9/I/EhYxP8eVXFnYv/gz9q/ZdS5QJM3PgdCAlkdMbrd7X6W52dQ
Q3PCyXQoYDwAG7CDJ7UMQoiGZl3jK8wf6IG4o4KJie0NkGluIF4uY0xyeyG+WgRJYD0tWCxh1fnO
NmAUFUjRSrfVKhGvvnLtPCo0AJk1YlqwYIMceieUPwuRhG3sdtSQqkLYbaNPa6Pxgmw2GJFRVNPp
1VT+VCX5IUDmTf4ioMbCFXTqN48Xza9DB8Ak6OPm2BEnGpeD3OpfcxnkhVFMpUW0l0Vwt3/VBIGz
lEhTAnQjBS/Zv2lhFUltN2XD7ZQ2FhkNnuIiTt6ua5GV3TY/uoXy3qCLx9gHLWAu4anBDY5TXArr
hCDe5g61b0SC53cf6/pgPN9hAyvQsNjqEi3/4po6zA3z9DS3Ewh/gu2Y5NjdottR4iaGkFo6RLmO
5csQgUhOzzrMwf0uaNwSk90KEwbtkEyWh/GlqBStlOmVhCxTYvbViqwBf1/Itcv9Jd3AMxYx1QDx
KiT1vmWjsBcqsKn2Xq2IutER6ff1O/b/DyigLXnoWUwLGokY8/EeluXSaLd3P6oD4R4CpsGkkt8b
BFHZL4z/Nk3HmljDqnIY7DuEM1QnaBM4kBEZPTfHNZtASZMlNmY8ag7ittsUHMhNqHdSM4YnvPyK
yjh7rXadElG2Z+A4sTCUh9485/qto+769lrQ4YY++xKe9bqegiLnW2Xii/EC79ugB9R7CtoYS1jS
lvIsNQMbMgQ6x5pHNViQ99KgG/b8MXUQKAeAODKVZPEQktKD2u6VeRiH/uDALgLDsmSphAVNTQmj
SaKwTr2qSdnZ5t6i4f4nlgTBxavQRsPi7jNKd0MasUhTPOPJoVsNWJy9LIXYUcHpAqrsA4v5hvEp
r6odgVbA7SA8QiQor929Tsu7OidB8d7f/HKGkSe9+QNof7lYoo/Hwb7kGML0x2W3dkBADNtUqO5Y
Kr83iVzsrbbol3pCouznFsD+HJxN9+mMPyhszagYNAxEYhE9jF8Ezf/Mrysnqg9BdHNECYAs3gFC
6wFmtmvn9ZU2Tl4MWpO4zAqTrcD0Flt9TtgxIOOIcoDFaVLy6LqpbiQA0vuP/Evrb0n0HkAz/YzO
beGw/JH1fqbdYl/Mo6pZHytrucOfYkMMsiiXyjdO9iDr3d8Z3StENFFhQFhlxE6sVm1AcDsRuRr7
M9HGo8aFVS/P8Vb3LDPLXPU4f8fItLut2MyFfma5cpnI8XrtsUBcRdq5A4NgS2qHei2fMeVB1sIf
lusHKhE6fKx531iMiUBiubDexUorCg3Q34ZKcJU6mTjt/8v4dPHU3XdXgKdKmWgfiSd38SjdWezX
8+KllqeBkXGr9qCeDbaGCbaBw3m+3GjS7ouacR2X1urRrauxqeoW9mZ35vouRufqhEtSNL2e0Ft6
2zQkk4kwqMgLhWUA7ls7M3jwWuLYshOtrWHBJNp/wONsUKZaeqqZKIs2ooXfPvUALzWuwGFAHV7K
azsQaygtmCKoKz2s00qoVIuEgPJ1BJxZaIkJRibiXaIpY8snro8Ksp7x6gXBplA1Z10ekHFvEo95
at4W5soij8UcnEMFMLutw6yyxnHhziYjBjtTfFD0NbdJ6SdZF8CQhhtVB+e6MYzemAm0IuwL0tO2
5v3CupxfsOXUtkUvjzxIeo5E3TKs7xtMwWo3oSRObKy+vj24jUK1gjui0fCVbIlb55N6nGlbvlKR
/Vl5Hpa8HY3OPT6pvzaK8mG/kBrnWBzhTLwrICjpYSE1bPIxf5UVk7QT+MTR1JLlgfNVboEq7gwg
ZrNG78BJ0Cqvli2M4nH0msDCY3L7f6Gxugnc+kNsarqqEfmgvZqgqjbCbAHCABhP3o/FaGw2dDzH
w1qfC5vUtQCygWCUbeyDgo0A7jn6NIS6MJ5dcW28yyIp7lNsQk+8T3SpRJomhC9xspZ9Mqm4alVm
dfcjplGKV+MVZrOlmiiP8IWimVOLkWzHk6hVjfAvjJCL40WURoRi54EVR4OY0rLlDG16d+m3jV7T
4+dxSGt2s0cNkXU+4siBYMUFUcfNThwNYPLz2gY7wMQnZXO8DMgYOcTfdZ6wPLlWdSmG3ypOAIE3
EYUhiWOvAXUBQlI/2fGGOcfdOtESEwrxm6YuJfa1FO4bBqy/QR+q4G6xm2JFA0KCM0Q/UHJrrqWz
l/4s8xtZENdS8SRgzG9uAiyUrW7Eb4yASqCmsG2ewNv04tZBGsj+GUwjYPIPlXfAJg+k8q7djrLC
tmHOfiIafuAGW/WFLVl4CNU9mnfXtwl9jOIQX4l1EOGBDteu0Ly3bMyZTWIF4DJ5XKRcAMj/SqAK
Dwb9TSFKd/aF8Zoxd6efVSgCinuLLW9H5SmwxCQAoh7NlGsmZTyKvxYu4g2/CWuPeQb078WJR9R3
3Ji3kK/2ArqH0DSx7TR6p7vxXdJZvzWuAZqxkQvgWOQFY2eu/sVY7oOmgCX27VSS+v32tBIe03T+
+KHMCknnMPsGQTRa7jhjkeVcilr6AZV4qNAsUP114NyrcMecT3ZMoOsfNzlrOMKKguRl0m1HLuQP
k/PU6leDA1PVreL/73s1uKHFSddAp5c++DGG2OTncczhi5WPhKTjdbuhY5dlfBNdF5mb1VKk52sB
mb9NTWuRsx34GwiG0jCD56IMg+WeBsoGNCLZJOfPUTX7/DTHvq8nMeqiHRuY2V5/nKWWcSARNebx
4K3gCuvhsyPcLQTZdDEquEnDZWnariyHME5m27L45cmDVi4cLswUQj8EibwOdQZYU1P+k3gfovxC
/y0ViFTEkZn41S9kglRHbQMV2bILb9lmEnkShVuf++uxRqfZExo/HGmzv6MDgrBZG8wr5HpWZL3e
gDZtFcT7aYm56TbsHNsSGDQU9RXflnR8wWZ04L8FLmQKLJwOAlR/W0AUhbBU0s5x2mX/i7ABPtzx
zaLLeNqXgb0p4U4W5aQM2F53v60HZoYjs2DP+dKAk+NPmsQloghH8WoDCx19fuCKf04puhAod5ea
aRs0E5TKfQfyvMDN5ljfAcj2eJuUZFhAj/B8iET6sWjcR9lrOktwOO+q/kph/fv3w+vXP/y6+ZaV
tQV2t2e3sGD3571rn0QxW8AO7AahB2ZR/79p1pV3aIX4+7jpwu+sFxHCjQxXqvKASa7jtaAGKUHA
1X2U2n3vGLBdK/FCaJIsF2/YrWiRkjr/p59MM6H6lk5slnL8aFfM8j+waYOMrAjIu89f1iM5ZQUW
oxKJqNW/JnT1ytm+0S3t74/CG06cSyiszxkKpZBdXwP2GZyn2LxttnY6sP7ZLj2ItCZaFWlWIe5o
GauzrbHZJsPsgdPlCm3tG2RzlkPwOXlriUlxJpULa1Z+l3u2UpWnMJuGLpT/lD/MxoWL5YE/gsVa
6sttMfZscQfel9dCXByxKmz2djKKZJ3yO7EIhfB5k98zXRGUCOIZRARJybM1IBoZ7gqJcQfIfXdx
Xz/XPRoJs3hqQHUmqkR9cQowKtqjwbW2wnsUapgA0ggJOC2Lk9v3Y5exTzLf8pVO/Kx5793NDpXH
KpJ5spfgx2zAA9d8SWzrdQ7DeDV77CmkvQuhW8mtX/R5wl67Q3UVDSnfYSi3rMU5SW3+IY4ICnLj
4D/kcW7zDZlLKXVNNFIprG7BirTdS2hRzMhld2LfwdWxR/ZfJSrd4PgCcY3B2rvQVTWYPExVhKo5
mZw3U1m+9TDls8NJwyBPnk6irvZzuFH1IAEcEl26E6C2X9/CiWPzaq8VS+iYuwS3Ar17q1YpZi8p
ou2tj4jyoeZAi91+GnOb4a0z+l9nKoo7psKcDYluCUtbuNgr8X6f1PjNkWbDWFpJ5avbJWQylxKN
yR5rrSUfrtSZTrafMhC0SmAfkwHVAQ88femt8KS4x0Xkkl5/QA/SWP/flrVO3TlT13DCSIhJnfra
WSysQlcCj/Sas296/DP0gDwlYkaLbDzZr5oEC/3Fbr58jOzvQcnprc96MGbZO9YH1RJD8esk+kxw
uQtg0r4aoWwWh1EZ38/k0JRZinjWofZxC+20ExiTYoKGhM59ZiyTAEJ8/6td6i7lQzJ7mnBKLkRn
r+CNm/B1tUjqiGkwdAeTUcAoYDix9ED8PQ9IVzNaI6uCPE37HouQpL+kbkS/Wtyri9mgh8I/NQy0
KLv0ivbBoWgwTK8+5HZG7WvyC2rfY1syuWiXhUP964oZFT+w6ivQL15Kf4Qwt+uD6n0JFq8RBZX9
vLsifrTsFQdvp4Pl6yo7KlG17cNz6LVqHU6HiXpFl+BGF3G5W0Y9M1MT33oRP6Vsvdn5B+M2eoBS
PrSn4lLCHGaEuljvUcRm7hWfu8WtAt2Janx2XPBCNyKS479IIG7SK129YIEfl2s8Z1+ru3PIS57b
0x5oCvgRFrcz8zkURRKjZw+M/hBGZRLqxN6Q9mO+ZfDbAcekM2MIPIE3NyJZjyIyHLtgaA2+LY3o
xTdjs67MYs7+W6XwL5ypQKaFc4pe8jjczZpIl3nYpFNXZRyB4H2a0QfIQ2+GqVC4N96g5XcT5pEu
YEYQzuh9uGZ5tkRgNGBR0CTEUVsopqmNb0W7I/vXinbmWk3NmKr4o1QdD3l1SkUEkaQbooZB9t+d
/qT0l7hESQrVXhEaiGzHQ53Mp4Sf9ujPJ7qrmwcs9zWBX/3l+JRQFo7UqeFXfAHRUhCg6LYAjtRi
fDzyUpy8kX4DS6UlgAtY4pfg/T2IEVkXXbe/csweakfsI/6kHkJdHXB+elk1pb49AHwnaP4NO76a
1kDLy+NPVRblUtpWLERwgeVpb1f69vVWYGfGKV/uVXUnaJFXFu6UhDpNNUvw002HzJ4layXoDztI
PWeDWXOC8ChrqTbjYCyEUd3zIGDQY/jcQQjqJTnlIkSfAZ6v7kt3+ptiWNdPA74+HRpfTYhRA3kr
leeNDcG8j57Mn2/C3FVNRd9FhjixJko005WvMVnsv4OkXsqW+xsTXtRjDIgZlQ5vU6TgAieKd03h
/WER8C+aYQhTvay6CEHD2d0nTsQsPJXS7cL9wENg4AMrYV5Bn+vLGNlVt15n8KKzu6D/2keACfYV
7Gk8pxQgEcS1tBmFSZFcZPquvzqDdWdPKAmbcwpMCaKW0JJfeKRXZgrqeHNpr/HqpZK0znpQklgD
8xPYPBlwf+vdML5g7JOwytcyMtj4ozI1p18ZLbwcjC9g0XDTIX2boOCC1PNdmCKxlWFGaUyXq1PS
gokpGLeNacZ8E7RlwtLEdMgxzmX1iAnFvwPqj4P5B62isTrI3q2M8NVYA3sLW9hEP5lvBKpbYdnl
cvm7zwB04KbAp1D/zX/JijWiGOpweXX3ftzIowm50NXucJTtwHgB2nxe0tZqt3srlyJdzGiXGURr
9g1jMevrr2BtBb5X8qEqUSyssj8BYQaVeV5bjKBiDYjd66shZo9mV7OeEN8GJ6S8E79l7gF0IHUe
6uBB/9FV+hXlId02CE5+heBKG9rSmzIMPoAGP5h169Ubzex/BiQsx4rjrv/vn4jOvxIuyMaSPo43
WcqTItRa3keeNuCKuWIKCtFEB1JL2mAlYJW3/mq+CJ5r3YVsYvFjnQ2PREZ2lCbL/JLgFLvrYPiI
2INvjOPOq5GYVY9fFqMrHg6c5gTpdE8RvxSg59VVdH2Z6TyrS9607TsmxK03dru6xc+IfImAhyzw
+r2pUXH9OACVKG9wrpzk6XSL9ap0Cz3dNkyl/0fLvl+ntpQAdMTMEyM3GLSPClQSKrYtV/Uq9CUO
8lziaOLLGY7UX3BHW73oTOiQVjR0zuoQVQ/NuBx42dGA/Bh3W9A2CivmwNb1Y+JZTFFLfN4Xojlf
JLDfrzu51YcLMkaDsUw2R+ROoYncVIyCjiczBXIQ5TrqsyCiRrBKFnMJyL+C11RjswlhiwR/ierB
wr6vESnRNgcojKApMUK8NCEhDyKNud94g5halOlDnU5swDoLJ17IYzfZvL44Xu0RwcaqwHXBa76j
COTbnVxV8N8JcdLBvvpoxCLuIFnQnkfoQEEycNd2xnERgGs1G7VN1hg8tAuxM+MGGzzbJnB3SxUp
BjT1j3bBA06F5yr1K5pCuB4pcfDTKbpqLXcIH41PPRk2GJhD5AgJQC2x5su8KuRG/Atn052SrO4b
dEijnlevSW4jqRbX9V+CNWyGKTQzSNsZmSQ0ILwKOaoEY+gCFH9mS7Bau75YOnUuEN2KFS275gr9
2k6Gtk2IOF5S0DE/ZZVGVbRPdrJwTEdEyiA/ydIqbKZKfqpK14T+SKWVcgPs/4LrEnKeeBhBiA36
TYnS+zXch1/BU2deG2x3VL8ORpQYq0CUOl/MixNw6GP5qJfNOrnuwifZ4qwiHFclwGs+MHkNsPWZ
oaNDjLmsGR0gVD9MDBl079sd2DzfKYL9orTbRU/vSedVRbyAjpUj0fdQmQ1t1K19+9JVhFz86/1Q
m593reP+ZosjBrjmOzMEM8HdfTLcP5L8/jqBCD5Ew8LMuMCPzcI1uPf93eHpVrM/UevQ2fpfMVPp
LNL6s5juxfORgeEQe4yyIZR5ABqdlolxMp3xbghln74TiBkSBxGFSPvtPZcfQG1oFn4ueFBM0L3O
IHewNZFmEccg0q8veHHJvsi9m2Unx2hcr0lca7h/isUeI6mL2btRW3BP3bBxQpFua5uVy6/p3Bw4
5k26XxRLblpt0r7wb1kx4wjdm3FZT45Zwu3WQiF/aW7uTWLZWArUXPIVWoT329F4yOdSKPrVlh0W
CaT+OvgLgdpO7+xIGXhwkOkhRIMpTnjkYg7DANbX/edQmnByi/md9muK814YC79TP8zawukaxP2K
HKfvJEYUhbJb3mg9wOvv3xvvIINk89V/AfTgpXmsROeYQiCbZmQVKFFtiNcFVeLjbbvSrfSchayl
2UKBPu7GGmrxzK1H+96SkIgHWLiOiqGrJeA5KdwGZiD9ryTTDZFbe0fwBRWQsroR5McF5Id/11Jn
YNl2XsvWN4DBHWwe6bZ5mWIN+OuBOEOUuM3CbTrNx+y63p/itdoGDHipti8zwN0POKQbZWAA2u5k
cmKfY+ab/7qa9k69D6eKqBKpA+A/CosIFLKJREzQ2XVsN+tpMID2oatJDg5Zmif7IRCR4qgMiDLE
RIQ/J0vCy6deeMF+W+lUXpRTuTAxZmYYb/QqyNRuHdstn9PK9nEpiyFncTkVwg+DCPtyXJMYf5x8
kR0zf2sJXqZ40/A5yX4VBKVQ37RiwU90AC/yyU0bzWEApirHXE3ntGZ447vX0+nekAbH/eFMIz9N
jNTOUv7+YEItJmzggJBr/PiOz3z5jg91OasaW+j9Y7+tGS+OpEqR3w1CU/f+0Onku+UWIR7LoQhf
Tw4/oDy83jvIgCkmhy64m6dMCzrPBakJXT2i+ZXKB1UhiHI1ct4Q2IYeSmtw8vcKUZ0VXBbgBH6u
j4r7JofNGTjlPxToAJfr4wg6QNDZqUCLkptl2nue/NmA69VoG4bLgWElcRX7DuupS2IE5cSj7Yge
Dkk3X8ky6brkek8r+5bK+pL6Oi9gQeryuyR07In+Utkt//Xu6MCBAOSKbLxzr6PGP2pVOhCRq1an
B116SNt00Z4/aDBX1kvHiXQQa9J16uaZwJ2en3KzBSGf7kWSb4qnypk4CQmZaewObbnjAEbCRV31
hxDCD01jSG+VIB0zT1WbuFZRGfkFrZb9KWdI/7wh7DJaU8U8UV1KlsuQCQeMH+db1sgJF8c8NFz8
u0XUecxn6Yej8899Wd6gzusyUclLVDzLJ8Lb4OVIOX1jyT/GVmX3T6tCHmlJJ2551VEGnGRiQu/r
7hjGhKZSt9EBRGEd3y6O007QNmwOOwB9AK5M3dJ+KccU+U58ggL0ZsjgMQBevoDkpdDQATNkQHaA
tjcB8dpAWQsxr0RpBP5HJvtjzNASRgrm73UZ6U2Udhswge7phkqL23z3VmfUBMVK40rpksAsYB0a
mPj3IpIdWpekg+sJmjLgNvM/SoPiQQne2QOI/+M9nc4maBg9emHpvlhZnK1Lzlls1YMPlBxVNo6I
wtjzHkNg77f2Vf+OZKsTPEl+p7Feqprx74nXVKnCmw+DBcV3US/r8TGhsLXal1An9O3GcpyAH0Z3
+HXIei7D5ObEiW0M0Z7pu06sqYoWaiCCEe7ORKEmUhqnGgDQRHkroScsRJ+OxlkBFTWX/G+YQ3vE
2c/iEYvw8M+7VAbivCvPTg/IhRv41G0bqZb+VUoEUWN4lFWcTYPJCBA/e8h8xnCxN4dUkEDNGCbK
C2Xkke8nx+GmeBM+TKEngI296mTc0eQGdYBRfYj5rX+BEt4VI2q0NGr0YJ1PjSfUKw3s7/E9PANw
p+Tmmjzo2G7Vp5X5liCTKnPmpIjmCOwqh3MH1+zCqOHDFqM9BWgR94MybM7yUJGqw0e8U58n27NP
W/KIGjpqfi21aCW4/GOz3qtv5qej9TEHXPXMy7x7Vfpf5vYhnIPh8qujVdjA9d0uMkW8pIfRxKRc
yBoFpfMpqb9s1MLJF19uAYlMAWoICmii0pGFedGz6//d6Rt7SZMWmHEXURQZS60TshUV4FNy0X9w
f0733ne0ydCo+rCHenEXsTkdVVsJRmFkiux8h70PiJ2kzUJXMr/ScnZoz1rFVWMw4Fpf3N7QXp5B
C7yfhbzakp96jDJjXguOxKiPiU0YaneDDK9aftOAxAj1IG6VZjIPJHavRCGqipJ0VfnUQrfBDQJX
8ppqdi8o+JVNj5XdC6PmP3auPYIzstulqoG3kqOZw/7q3+la5rg85gxtZ3uE4G9yCrKy8dWETBCH
gVwIlZ2uN7ESWIEb4PaIuiBO95wIv+LdrenWnuUQjKlLuNY093sOZJXOjeRcCsT//qr1cn82uDhq
Uxr+lRjo8OdcsB9TmY6CdLujDwJx4X/giRQCmg26UNkpKO+TZoc5C9WKTtXJ0/66+kW2aPP1cPXc
5EkscwpLuQ6Wcq6tTYQZHN7RC95vagIkan32ESwTmZrfoYIdUmOkBUR/liK99lDdN+4tiO5HDTy0
1YYab1s9CEwZT8EDnHVZr8SkdO2s9b0W4rFUvLO6o7f97WDEkIR9CPvXJbfuIgcydXutxatezfnX
NcN7iGZIrgk33VJ8nj5Ht7vCP2LcwnD6Ax07gKIJt9imlCWqF8lHHKVV1uOCtQhu6Kh/sWoTsdcw
TkfMZaYI1X1obcOCpudV8e4IekID5Ys5urCBZ8Z3mB4PyAEnSHWMJIvdEk3s6xkzDF2/0Nycm8jh
t2Vby3oNWo4s/jT2HEzdeUGwdmYJ3Zfre8Y3ONCXAYHt4hmP5lGg0Sx9Pbsw6G9pQEio6jvKwcn+
zWvvSQyC/fJJBJVAjMrgliLhZkXHb1jmk6XLcuI68sofKRkrkIuPxcmGG773pIW3RswCkwnocsXP
5PlcdOODJybPCwdFF2OHiYxifqI28fd7Q+sEJaRYk8DbIyITWvWxIB6r6bt1mfsz56Q89vDi10Nj
lpVAC0ghCmenGtFD2RqG3F6bUo267qpH8RiAkmhtIniXdfuPalejLnt9AnzM9Ifl1vCbczxws+CS
aEKWx6coiQDmal9UVsR2Qyh/5W1wAbA8xSzsxO+DC7unRUs+QfIUSKCox1tfGCwyXMFFHpHY93UG
xWuuP9kNfp71q8zMA1mw6xyoLHvC1O9WL+ZcmjyGRwuL2os5Giki5m14quUjh21ddT2+TTzvwqpW
tv+6+WVdxIMz6tXW1QFSWivWrv2qnoUAlnWr4jVYwB89zzQ2FvafgoMX4RlT42bdYaT14vIKI2SM
PlaxCr8PN8CEH2Ubyr+73ce011zxDMzBS26FPLfO/16NrScckS2iRIwDsd0/S7qt9N9jS8ZvFP0Z
/GBQJDZMdAFkmn67gs2jy9S2m0bngldrf+5Pg5z0VjBWmkxf8pDwOg+moghKvuVSyiPaETYYdHP1
Nqa3toTS8JOInSeRIFjWRlrpd58fBAYunZq//vEhqHcfZZwjBdB0jG2Ysh7ZgfjQ9snDW/aahN2T
EmIF/1pno9USkvWnHTW2Kw0ZDDo1vdPHdjHSW3uV6vjeVAGfZsbaGOZ5U9PIVORhFsYgbnlTOIPV
VxPhAO+zR22YnKDKBCRLSdVnUj3LEl3c47U6k6nmK0rjSx6mGKMMEcaaTkkUGJDhSK5SU8EMgV5F
2LjSvUsve7LXdUuzqszK4+rSgKedPKFDcWNbHGTNbt5T+HZpTNSc+qaawMK3epCaMmBxPesFoVFE
Fc4UdO4XgajvOgIordOnCPMp/GqaaLBYIh6Uxp1r7boFCVZxxTLbEGQ43AEIXWkIW2MFB1doefsZ
CcEbRiEe3euozAaVr1YiIY8WgFd8H4x4FeEAJ+WJ8flt01fLYQfFjwzs9+duUa1w+44KMnwan7KS
6DSRCwUr85Aed+RIUGc/X9q6zIekjdd1S4S3SAIeUfh+0aHeB3ub1P3f5Kdvp234gOEnz2eQ8gYs
LypsIascX+cnC24Ihk7jq50vRXasr7nubKHIbD4jQmUFTgqCYIxR5E+rUBsI1fQ5W/f0RbJjIq71
AiYrWCzsGxmqlVHm3p8qfiGMf1Gm3ZjBTOrlwALzdVQVQFEvGpVAkorxSQi8Fi8EWRD5myzEnE6N
hFzR7kGi+SIyP72T8A72UmCSRQebb0SHGLjeEaS2V3HB9OfmhLDuiHdzAaMdj79SeQeDLft7Sveq
51ss/8g6cY7jh76zYMboU+IHfYj2fGjidRZBsB5LqGYeVjxwTN+lEBw5Q7EPP8YNhDrtZIx7CwE4
qpjSEw6u8S8X/216Mqm7d792s+YlRIin3tubdOsWHu9PB4tZw3dMddDa65oNqA11tCvuv9uAOoIx
sbFfnfXUTk8jKaE9v1Gejc5iphKhMhvJyS/iOAyYTY3ITeB0qQLESl6L0srzO9Wgqvh1+XPn0+pJ
HtVQmt6Tt02xglBUvgNy4f2ptsIDiibjNrsd1otnSIuu4sGmeQv/Fp8aYzAVwXe/jeaa2uKVSENq
0rS0OtDuy5L2D9WVQTWufmcb9R/niUcrbs0VziOsbcvZNI8SfTCJTN1dyzR6+cB2JRIhrp1UkU6z
p/eqf1F+6pSGi7zYpi+PvgUydJyXFuivoWIQCEIXs1oRa6cKI2cH+pzgiBhiUUwmd2Y1LH14Zc/R
ZUha8vtNNYEPcoDvVptun3/nkDHM1KDYyxt8cVhZhiWUG/HO9LU+UVm3M9PlBUVhjjx3cJP+rH6X
SByEvjW6WDhWGfeI0faC8pvkiUzK5kjyngKGWtAqU65cOOPSqsfLQ6l1LWAFmcfSW9w7UaGOTgAd
0KCcvEiDzGX9yZLIsQvEIcL5gCB9XbSPuynNMFL159mhrdyo0lRhydp3lEpzuxjtB5FFdq98gDso
UMH4goXdvuP0R6RbkDNTxr/peLih0kTY+D/N0CMwoxBPL57XaWWGrHhA2HmSJDMhO3bgbr7W0OzR
D2gqGu6Jcn14PjGcZiobJ6BYBpyEw0rzuzKaYyhokHGzRzlgrV6AvNbVcrpCQ6l81SAwTLayAy7O
kFvSsKm8xzoH2NIjIbCi5jQcK0LfPHPmlBtrnVIXTYk8nDXBtEmRS7exbPTOePD1fX+CdIIxUMs/
Wrd34bd5Ym3gNU6Q2epC6OPIuaCWqxiUduZnFXkDJkrg/mjBNIWOvD8zDEERZ4bhWTH9JLHb6FGZ
tJnOX2L62Fhgj++dRMaIQ7SdiTNCLFkH9PQuendPCb0yqpny8GuTp19LfbbZHPxjBlvqAZ5WNiUN
pQQg+Tpn3v2bsUHUQVBJ6ZWM1j2y8zg8MfowxJabIztyO9Lc6RpGuhAoKpOndk1K+4ThpQc5CHNy
eGVP/5auMM/C3m/sYl1ZyTqF3mYAo6VytJH9IwyVnwwKykFP12ON6QsFzgA++gZ0Z5Vu8oLTJDdq
02ToYYqBL3T5o7JiK1Eop39BeKESzDb73RrpnC7II7uqBnJm8pf4Q00ZJaFAQptq2Q3QBiNQPSLd
0EuRr14lbOInZsqQAOuN6LBvnbw35QTDZkBYaqx+pVwXql9t+JY/GOBeb6Zj9rELLy1H5Ny6eykL
mnHzhzTUS70q6u8u/z8R41UzuiL7ZiE+KvqJIlWXH8oOGB+6zZQkBvwBXmGuIwkHf1x4XwDCFeC+
Anc19ekXEpMqE6rKU+XRiboBhrTz9OFw9ChMM+oKyH3NyggOGYWO5C6WNDGYrMx6iETSVYEbeO5G
Ld8+UOXE/sEf/q8eXEhqYwCIuZb6r8lqIxwbLkMsxE1vktPnDnbDBmMl0AzCynwjhVJ6Q0GWxyq5
uhK148c8afMH23w3ibTyye8CvVbqkygbi5sQdpSXAb7zqzUkX2r4hxea1b3Yy4TXsVONOD3HMHoY
sRrWxxmi+WVMbYJ9HuYDz722sAt6X1794J9aoT/Cje5oOLfWrjX59SChgrIq1Fyb145+WFfcSURM
G2V/0rNuEPn9nfWfONFjG9tUdvVvQ8E/xJHMXA5PknGMrl6FTMc0Z+LSXfOSnmBjKpdqpHBYNf1+
isG5WSXdUpjO1JI34r1EIf9UFFc4V63yvSnK9Td8UOyE+bOYitycCzddli9qiU1B004K6qasbcO4
iuf90CNWnRVezCG32TD0deSlF2W1dJ/t2VRMZ9bL+25U9zoKx8kY78TOEYvuq06f+70Yz8b4/wmN
okNE2bfuymgiUjvYJOe7rs14NpJclRYotAx9C1uEeWW7n+Bu7avznB90PGn7A54X6d5y/lLU0lBR
LzdfS/PXfBKp3nryTbKIzxf5VJPKN1WOu6HK1O72PWh0YZwyVgdVIgJLSLePnpt2hXq0GEGxe0zD
zK/6f8tZ2xpWk+8KrBMqCqDej3E96Z/s70XA2WgK4Xcistiyw+SnHtH9bcyxi4cbSLwB6XdCNILB
wXhppiDdPTn2JtrXG9Mb5l8bfixullZ8IS5YrEgyIvGCXuLsR5J40o99GG5MUMC544odkzO4+sdF
II7va58LAMf/Il0aBTsbp1agaMlh4R8rf+40yvOYwCRU4EV+1mTTRJlHLuHD93NahG8DY0nIzWGr
xF495k8hw5d3P4sC3XUMeEuugmG4doX9Gk+yJFW0SK6/2WiZ7Q/QaEGnaleIIKlr1lFLezQwb9y0
++2R2bbDHhDEyMToFG32jboW/8GSqBGiRur7HTP+r5b0mJXCk1ANVqySwF2LcZG10BrZGLzJE+ci
ShpA08RTjGkAMr24OD2yNwvWayyB3/NeyZB+4UY6ksi62F5nRb+KhImvWKEBQIgr/0bWu1V2fNiK
xE9+1EIl50Ylk4yt+aSQ4zo1Wcp2wX/4yPy3RNyhOf5Gp4dBZY+SXiicsgEDubq3R6N5THButHaO
wNqZf4qWnldJGVGobIC36wVHWlWJGHLVKCqsUaaP+89vXqP4JN+Q6s6xQIHoMJsDKlUcUA09x2d0
WAVPEh0nr7NGPp20mUR95YzcU5AftgZJSicWBosFYqJB08xFmiSsOcyPJueBuMVl5MH+N9wXvDrx
UKlid/+yJ9CVWX7ZKRP9cYAFfatgeKyqIS8KzwHUWLcqiFV4BloVBq/ZGOfJ63HMe/yRohBZu2Hm
ppW8j02x5YsBl3d2c+Lqdw+03OL1SJn5d4kHvbW11wOH3cVj3Bj3F1iyS73djxpd7aLvJUa9czYt
2qmlVkMIDjvwsvrjmPaJF95NGG9R1ASgOG9kUc1lCQ5TaGDcAIdbXKHiRscwS/Q8TcoOlNc7elRn
bXcwW1ktmNmPoPTc+1sSwxLUmt2zalbnxODJNUOqKd2alUYhc27nbQcGcGz8YB+rLGKZq5BqdXaA
jwhZPNem3lVVQTYNT67u/M7OKvh211uf2wh/R/A1IawlHrf5w0HVloTcF3w7+OL8sPfiv40NSiDh
kY1IsMKq1cLqD3nbvNauiudmoMdTtaWqX5KFVmcmqlb+ySNBRWYYKQQE3hbQgDavfaNFq2ulyooa
nyNBefrJ1ngPZ23I/+Tpq3WgDBPF1+9rE12gsENEPyOlORhBkUREUzb5/OLPcuvl+0oDw5TmpTbG
lsMUbB+c+TB/L32ZsxAWJFiY7t0ijaoplvCZ9FPOGf52MMvYblBZYTlSXSMV9iAaUByJamq311/z
7aLqp+PMZfr2TQ6XG/Y+DqavkKwsmEafDr0TticrS8ZWnkdqYo5xcSvE6TS3OlAlnJlftRsNdJv8
ZRBBnmDVyiuHzpDlj2qU0E8W3vYkQRTcVq6dNQ/SWcbOqDxzNuZfhhA/1OaJBLndgXujoas1gOke
KB4kUOr1ga9Eb8031odBiLrqtgiCYB3vMcC4/uSNa17Y+9DPTx1wYKG6lz9CZ+VOHIF106QEwvQq
Mt5qX+Svy2Wk0GDQNUfJ00s62nh83GZx+7apLLxV0lRHE5XNaTE1kl9Y9jeDhwhm9KUWpNvOQJEG
MBWTGot38D9UwAiKpah7+XEVSM1ODjaVTsGoLJQ7UQWtsB5XDB06JHTQ+gm+s5qTcA0xgdpWCg9G
kF6bOJNiT9jq2H/4wpuj+CTYluKB2Wh151gmW9+1MqvfjEHONL+D3w3AXTz9SH1F3+9mco9282jT
NRSYTQVOPM1FfCM+AwCCYC0VMyaPyKI1EdPEah+PZWe8W7WJ0jNYks59SzjqqmoCM8io1DqnOVk2
ZfRsEjJ6crc0avTStvOYnzkcaY1xF3Q2VnK3j9UHtPXO50AZfEzuxPihHCwg/CvscTq0XGsjO8LQ
xseaMk+77L1PPhESHqkz2cOhOzSDV6jXOYj97BXHNYUxpz8zYyNPCNqd8WL/ef6oS/icWRjTJiLL
0VN+04QpATWwjgLeKn52wzlRVNnag+RDYjZ6hJWiQUk/ZSEe1mO22l+nFeNkbPWYndx9gSRKzeOL
QuaV58qcvr9GlldrdlaRcILYHdOFJTR1Z2EWxbQ7dfkUhG+oMN1zoDsI//xmS4bIi3hRl+W1TtCk
q48JGdbLLANedCmiGhCwHQ+yjaZK3HRyLcAtdANIUsj8549/AX1Q4BtC+0Y79NJ3LeIY2fAxNdPW
kHYJvKqAJptxTP5f+BqhTL9hDdyY/q+mtqtBdQks7M5GnGW6q8kmIOSSxQDla6brRr1jV67fekPs
KzL/+/8bDOeYRpeaOwlcyxvG8S32imZC4O4BgLFnkj8ZHTzhE+C9AxGLrMUFS2NBLvDT5sApz4SQ
VW9OIb9xr+MK9tVTaxKMglCufTj5wPYKqyfFN0VFDqAam0a62Eg0AM4pU/VQmTLkMvejixd9mByT
E2xph7V1u5n7u4rG7btrxK/iZgwkNmX3gBrxlEm17OJ/K/Ut4h1lG8VadeBHnETsg2InHFEpZ8Ne
nA7LdIybGwMozB8sas6jA86MrAqnpV4RcltOK4MA0wF6ZA7cp9x138fJX+zHYKXKouuSH4q81pdq
n4qW27b35pzad88qpfxnKZlyNlV8tWnvZ/0cDsg4OfvqOxQc8byFLtDj95yCJPH9otkSMcv0WDzI
YrJVjMXK61EXpn9WATGdbMyKGPQG+ftzHdWYvjQRlbMLpefTXrZ0NOPhWVcZE3DtEEfCK2GzEHCE
mjZlZRSSEfZPIuUr1HxrPV1jD2So2mSy2Eo0A8FjLnD95+/U1WOpnSDQfSK/GSwo+x53zNVDJBH1
68wxflzb74ob/MCcnDKzZSVKVOPK/jYOGPUcdPn10obv++AnQ7T4Eo2tGX5tqlEhrw5KM+JnU9+I
p24pDPvAWlf6Gkq/FijpU+Eat4Hk81I7fpBB/UNspavy6k2ER0Azlxw6IKRaokaR4llwNTCbLhc1
khrMcOME1GTpHeKUVkbtPkfdqmHXFc5a381/OQoeBdDg2LrboA5QtscBFfhirTdaDkPUT7jczAqY
x1tIxsyZRZ2wD9cWhnmqAB+UWBtRpwGh1xR7H5HmNG3EYALeThnl0Je9n7XCyyRQNmnP7IKCIgff
tmqdc84GHC4rhQ7UKkT4I/9vXmCiW4SkmVMdMe0dnRrWPZ75pv2L66PPGcbgyWujw0OGYGpNjVEq
MfwAnT2HYLWoeDUIRMHXc1PHeRUnxWNqmhNtu0sygo2fIFkpPC8b0KbDg+d+lDpgJwnj4p2tfGfX
cPrkuraHfu2Vw6/Wu6/t20OwHdyml4KHr4VSznkXNan/dveXs9GVT8UPVw76EdJusks4mJ4nJ9F1
rEkvFwphhk22xfm42t71a7BsDoy5a5otrRlZu3Wet8WN0Fn3aU6meXACralVXFRSK26UnR7QiIJ8
wVisde2fOuZRrufNe3XrF0Bllgb4JsrmxYa0zYB3DkRf2DTO7SCCRMZbVqhpo2iJZeFb1OLSsfC4
iQvNaArvn7GIvtL0ozGzRQrVyl7t6W86SoXyWhPPlzmL/NZn6+I1A1a9Q/wnnPV5pto+qGSKlU48
bVBBbVRYFb6T9S8SRXwewJeGQzl3GR7QkflETHWG2ytRfxIBch+qABlkkZIln353v+54fMfaxkPs
UrOvTpeqkTJi4ILJgeLn/QyKX86cmZQLIxfqezVoP+U0ogAZG/fEY0celEjesFDFST7RQf91hThi
BY5F+aZMsVEEI5UYwWCDIFDSslM/9sj7a+BFXwE5J09nmozbpN4QDlhVBlYRDaFGkN0mID3C/HGk
pQ0YngM3Y1GBTzzzenMkicK6/Z2A2LJB7uVOR+NbdiuWPMLjh5bnYZVhEu2A9xyXSm7oLMSz2+Lv
VnbT3eJkkjSIPLcHM6TfOiDWvaa0cuwZLXIKPjFqE5MAWYNjFQGGSIUcHfS6gBCUaqD0wltf0N8d
LeGxu3PTTP2cw5OLh3CD8BfMPj+K49F/XZktNuEG1A4kJcJa5bPs2w0ZZ3M13+OvLFuo0M/1dnQz
728PVRFqwPo7x6ksYcvC70/TjCx/jbtWTvww5E6S/WY95bBB9GSerAxES9g+glT/2gtzo2MOjRcd
uNfaAnO+RDvMprRMKH8xpveILGHTvRp20LzzTorAIJi86t1ikKkbNTlxQ3aXX1L5FHyIlXthJKw5
DqLxGHDg+q+xwzt2Pf8Kj8RFUzWpwmVWFRSj5ssa6GVvcvVzBRMffH1l9X0dKg7/06Q+ZVp7l3Dh
dQ3pI/NPWT5qH2csrF2YnhbD0dklguoJGxTCr9/SPLIrpgaHFSkJgbzeDnBajiS5RS1Br7YRZBTm
01Lf5nJaKBFoh31UkESe6yzNz944oe5bFlOThsaq98iakKMPpAQPx9mrPp3zYX6exe7QOt+ClGnF
CC6MVZIYqqdMmZKtJKPAzB9CXnwKwR5XYw61lsiFZyCKRR4BnSgCoxusjx9CkYkJEFdanTI98wzx
0/V+ytaGkCfDoQRoiyeyARsnDeP9vD2TZCpiB40XxfUsREw7M8qQlUPy2aXllM3UYtkwOuZIlePT
EusliFUCUfjZWyB90O9TR//aSh+N+IvaTKR0b5+f4AATDO5Ur9YBmIeiGd11P3BA42SQ7hAyKANY
Hvuq+oG+Nsb5HQZcw465MEfHfx+eMmBZk8wgwckYPPpu0eE8LmiHhSOxqa+BWw+g2RzlhqO4Hk2B
xPoPdf/OWsPFK5JsQ95ISvFPkTP+iG3MKDmwdY7EhDjXOxhSJ2af/mi7d4ahSChetCLQTPXHfL+2
FulEVCVwIRjNbTBoqfyOe3X31ILWA2z9NV2vjYPKAr+7sWIRyDSww+G5d94ZQaZL8Dzd2tJSd14p
8y0031P1HQlMx9sJsT3ISUOb07KAZD8zsHLhPTuStvsdTftW3bgQ++t891TnuO5NPW7eMs5oI+Zv
EVC2Ot92E9K0tsw/1Wo8EZvKDpoMh/3X4aU5Adz1zoOn1LDQcBMUJAM4G0BcNogDX3oUZIfhPT3W
2vikG9Ju+1hvtO/4xSVsk0/2XxCopdUa6M0gqXO98o5WoCKb+Ae36BEgxrvxLJKo/35Lka5Ih//J
zQsbS+UqihAbIM6TkCN18qXfTDty8mnXgY8+ttXieEXaMk7teF0kRaBAAmBV6YKJUbDRx3TGVyBD
p7QX84j8gD6uX6zIn3pD3rzLfyWDlJs76EcN08CC6Eua+s2KdEKkP9Wa9nbfJqtLww+ShO/s30z9
H2jnn+6KARMc1CLl8VpJT2u1HJg53O7g9TiAoPYr4Rp0fvqpwQx/NJROe6TEJwe4Fx9FfvXO5/pd
MdAQj3EQNzosWPYvf1C6BaYprqL+Dixc5jw+VQ+tFb6i5iixLvQdj5u4GgW4GHEaA56nfIR5hg9G
sDtzrhjfRkFgqTySffMLRxgF9S9YMeMRx8cpDZITgG0o5JBCPorYs9nSvKNJpadtf3U4b8dbSLcT
tNhTiP3rWwV6UiWNOqkLtlHU1i+g8FP/Z5vogoIBGOG6MziGRoHEnBHPlF3gRR4p/DvYF1nAZDIi
V8s0cuTYtoZx8LDiP4uz0xt+lijOsLNZQncdf5XEsTfhZSrXRfiAfHpfa+D5f0/jyT0cBJBmFNNM
U5x2iFbyyUcTcrIAzpc4Uw4mQViFYA8v3ZJidlim7kA7whzta5tHUfpCoH0yH/5S74QdQv4S8Uh9
oEtrDWSCx/9NnMyUXRl6GIAGKFKP8DCttX5Unu9MZ62sBz/h7hFOO9QWNL5sRx821EDLg2GELWGI
QdNhpEvcssLvkxbO877cug3LgdrDUYiLXkDaH5bbxiZxaX2s0KcK5O7Ou5gxMhvK3xsssycIUOBP
/0hmcBvAmcKJP+Z0AqsP4Y2dGnc3K5cnUqNSLHvDLWFe1v0Zxo2DeFgyP3ZRDE168EBo0lCj7NIF
Wir5UJMx8q6JV/zPbjlMHoDVd+zjHxniSaHoMfXUHerbrJ7UIbzVmr+SFPl4DSNJCuj9uwHT1Ni7
/ZhAhyYQoDEYeZlZ1HnU1Msg579cGC5kiU4HFLma2eaGhrMWViVdekTdHmb0Tte5wtOUiYgobhwv
rFjBBZ2hDYTSWHbcfFmb08yesabnZh5RPzoNDwWFyGU8paJuoK6HuVFPjSoAXrjHFQfune2hqkSN
vsZnFfFJcr9GVvRx6omXSZOLLxEw+34WoHjvzDhsXTAVsfpsngZgmxVtJcYEVnGaadc1YdnTESkX
/mix0cbYeNvBC3wnKWZr+9RHk7JkDene/9h7K/1hSSY4WIyBUE214QFiOnfPZPzL73B9ZdL0EqaF
lgAABCg31cp4h8VARU5bJdwsDv/DjkZSvuPRwWLBTb02aa+B9xt/RD4FwGWvMdcx2n7m0xyitDN3
S1jTaAyjx7IwtxAUuo83ObnQM6bj8OreGuitlFS0///yyDpLVC12FKYlSvckPxTLBQ9ZLRaZvWJ4
+plr/TEUIqyU56M+fdlmt6vPbproVdDTz2SYZZWQABDY+nwKvE7qsqU+qh7Vh0klDQ463YWrN1WI
7nIYd9X49i5QOIPV88b9szsYIohtdQ1mAx0zGdopw7+2ZCXa3f1w1TPX4L4dt41lxicQ5WR3u19m
nvJuOxM/ntRWJjvuNwKtKTFLf5vNVPcVEvkCtaISWh0JzCfmTPruTx+QTc8tPrPN6VMJDxAZpH8C
IBPHouL0RYZ6wyqZUwYs/oFMf9KrI3NRuOLPeUr/G3C9p1vUgTD922fpVs9ZDMcVTUlLIaJjtfbr
6ifLB+qdZGdVcvl7p/W9I6mjuvvZn/0n7SPOCRCfyxUtQ1Ui1S1vvVZyYDw1X5cA8iLBXTkKZp35
EKixf4xAUzAFXzBn4srfGhWQOITXStu1ISVnH82/gCnR7jZaLKGD5Ne0bo7IloBv/y5qnSLAWDaa
2DM/FEA5jomsWqduBA4qvXbGVT+JQQanitCgxINZYb2SCYRQ4Yaar/QdrzUOVrqZzgLpVDK6CoIw
aNjiYsSkbzKMDVOvy/L4x/766+/cSU8Dam+vNvhQJynrsMntMxO+2Qp2/oo2LWlIshN4GxsdvDKl
sfJl5FiKN9mazeqFofZT0yRFs+nY3/93HdofPv4EdN3xYU1jhO+vdgFEpsq6nHfi+PfISfnjCTuA
Bf5+rxoaWdZsQuBE64m+zysro2/a7DvMwTT6hYkgo34VAbx9csvPtKUm18IG/qOAYE46FHqQ0r8a
Ackz94OShpuMAB7ccXxP6zRu1OHTEkSqYNLmZMhVRkZxHX8k6JCCblSu90HbW+WhaoSm0Rl/CKu3
K1dqDLikuwZGbb0zhPKTES0oo+j5MG3XU+NZm6O7T3aLjhiZ78I5FrtYMeAieje4iREVE8m0an3G
YvsY56UezJtSKjCvU2JqNh+lq1/FFhqGlMhuSsPxgqecasycEFYApRH1gPj7jliLwDkhKz2CWE8J
mZ8fQaHtxBb5LL0NFSBOD0xLUskr4C4L3gxrJzvHltOYhUNV3PjJsE0Y6uKfqwZtAy4vhkL2r14r
CNxOKv4NDs+2pR/GCPcz6n3SuJq9cncKvBD1VdoACMu9UBABL8bD3ouhFrxUONHtg97RIm9D9oIr
60ycuiDLuWP9tpEkVzKfcj8mVJ0rY6NJ0G5g6nRKa5u3Tz0q92FgZESdLlgr9JNjW4Zn9H4N06zY
Km7R5ap5VBU/1HXNOfMzkr+5x1bfNKrtGEQn6rN2vIxR3gG6s1U2xcD0QseRSwmhd09HR/FoGSDT
fcKSU7ZJkgW6peILg5UP+qRcBwdrQgdw4nE2Lysz3LHoDtHOCFxxRYq9qVb86ERFyO7DZfJob/Bh
6YoxIZ2upDz2t9lA9enp2UtcKIjoV15v9SAsRRyLtqSaWqnl4+OxhpT8qf8hyEjRIRU/+h7D8+wG
vv7nxZL1cuNkSXLefMuteGP6zQSlGbNNyCKYAyufHpfoz+2NAjFoXb43rrZG/BQFUG3dTlAZTQ8e
WtS7V+jc57Xf69irKAgDBzWz/kOxi0ihdGdJCblIPWRGFVMnjTPQ8sFJxab3JJPjSEbXET40p6iA
JffGN+hbGnp8rgnXRbBIu/HhqN8JKgn4NW53fYLAmtev+/1aQF2gwm+U8+X8s/rHevFjL0Thz6Zg
KMvAg5a+ljPn5uOpuywBMSd8LQuLZlYtmXnf8ndLgnhQJo2/+rHfUCz+4biQRrJSUl0exy315C+D
7StJ9rAgBXxF7AbgeN3/rX70FAYvxsw5d/56zw0jv1EjZVYgH8qBnHbrtmO/TpzMgxe19QOKY3Sq
xLVZBidv7Y1edfuagf3zNbBm1I/DWJZh8DZeE9btpoxgFL6D+CM8gV7kjVVqu9KZex/iQ7dzISha
MKFGj3+G9DpgXMnElwoDGGZ9PpaPehej0ZPGxQWDtGwodcmN/eykb7iyTB90islqOrrsrUKuGdim
PT8s1Ar5iz+jVqv2wNfwN3tGW1SC06ykjbwQXZpi4JPczt2AN2q65ajz6k+x/gWJhhfbxkB6ZFN+
DfX3t31ScqHy2kcxb5rDNEOzF7md3rJuJkRjZSSQ6mry+3VojEqR7rfGRkWnWjUd4r0L5YTmEjYn
Nn5wQweiA92VQvm7+YYdXj9SarlvGVGU/MpsGDLOM3RLD9spo+aNj3OxC2MK7nj0VQevJSpXPpvi
JH2wo17+hBfCDRNG1z7H1lETFfwPRP7+fAKyv9LpVhYz/AiIpkohsz/Rm2haEcM95uscYfsvOKto
YL9NvCes+d87C7i37WxK+O3w9Xe8QBYjUOkzs+Dg5WL1W5m3PU0AKpaSVaKsI6DLsrCJ4+VlmKl3
4pmPwjsh/3sLkz3YN/JhuSkZZBPwcCUJ8Zvoi3AIQI9fjh3tiLKhzMNTkxKfSIv0/jWHuz5AAhG2
i8iWn3iYhMLAph5e0cZTdVgOv6BWKSdwXQ5lHIzUfskrgkevW39T1m5Mf4VQgLQsf24+aElRmNsi
l5l5zWLXpMEl6OLA32PFRlBbGRwNVWFye7sO0B/ol86vLPC4mAaTXbs7rSzGeXArJtk0Ch6DBBG7
VDZauRr0xUHn5kopJwf1TU472aWCK3ZydzsqoGmdies8iwvanS4F/EddAqIAIGPFfRsCcX5GhwR3
44dED7WtY7NcnpiZmnDvdKR9MaHYGV3LcHQVGRiPx7nwmrOnblyP85hqF/iqojf+qCCWOjB6m8gu
x5fq4ElOkObiQ1gNR29sq4XCiYaWIGMDc57TmK3YQJcrc89Tp9XqQwAWTzdnnX1IAVvy0I/JpOLe
npQ/4NEuAtdHu7vHO37/8ocFd/YKSPJZQcMx54wSnRae7F+z/QsMh1HZTG3+IEP9RYIRt0JMuH46
+0A4uGxryHPdSLspTK01KAz2u8hHXWVn8MC8IZwiLJXfcQS0F+Yg8KtfsWmV+jKkPOWFSMZREX9c
sufqM3RyojwJvjblOghdTPeu8WxrhwENqWlVut1eynObHTkJtiyULLRVnsa+gvbSZPrLXx2Jjau6
8wpjwffPTrygB3LF6WhvoXJgUaguKhwNpiRMKk9SRnkXBt/iZIrg6m4by0Ovj3rsa3k8F4pMKazi
BFPFCIxEiU/umsnvGvCL1vDDQlHrDX64SEky/ZvDXOfKlhAqOzsxOAO0gBC6agQPo0JktqH7wcTd
lNMzs0xpHvuS+6vl+K88EUYTePF9P2Cq3fgO+Tj+jwaczGLkb3WXmY9fCpApfxkhFFZpB0MHPx7Q
M9xY4/083u53HNM6Wd3ZhLPMerbsW/zq54bW2zOJcO02oMDIUXv/cOc/KwLc6IqtZY3hFp9ZAX4o
gIGTT3polwiOMbMh2sGKzkSGNE0nvdP2KuIgpEKlEq69G6TObAzOyMzFHQASg8LRdVUYcZVh04XJ
ijHsE59J1MxnzZpDq/1/GCKrWVE56pwkkQHJJ1eRdWsCLwAdW6QfoO43N9zRujn+ezRN5V+jN/G9
TkYEwNdXAlvcagrLv1OLT5UYNNeLqn3U6ERtj9YJPn/uCFDsnz7rQK+RL2s/3osewxdc7DT2Dvb2
VBsrKKblHokxczo4OqRN9fI/fqmx0l4zepe3TL/6BoBqXJlCUtXJ1she3YxHROen0nOk/+sauC4L
ihqFZAKEJfDwC0WF3JBSCgjaf7xEYDzzbRKqCXzjgVuvpYQTP0YsDrZ9HDv7LDxbHfhHliu0snD8
sjWGf0NTDnvaszPvzXSEFFZZSxaRORhOuslHqdmI5PoHlNnpXZsI0ndPMj4WTwHM/KQUYh+cj8zq
hj7GtjVjYRbvhDFk2eWQ/z1ydOBAHIL28/7vUSPMBrZs7gXfYB5Nx54+Eoh9rCpTBU3KJfJ7hzp4
V21Qy/CK0XMTHvX0/8s5nMadv+M3ZKGZl7e1vLW2Rg2He+QBeSa6UfSbWcaYqWUtVO7+yJkrTlm0
Oc/bh5d9rbcBjXjwtjD40h9uQ7hOBvs/wfUd/h389e43th/Z9RZO6cDjEA14bkVwPGQPcBoOIeae
n8UwP+1g+8rqQNNabsOORioB4LYbIv7oTHyh1/FD5mmFx5RB2LbLawIgOzXaDINS8G18ELhbZwCo
HXZEb5BqrSVkQVXW12GGykr+MDy8d03Ml3D+XTcWv4CFJbQKsoLw/zYXJW//+/68qnH5av+bkfva
WGmKWlnRdZ+sXnRSJM9LKN4aCOPTMN55noCZp2PGL3ux26Nfqb6sLulvWPIukNpS1rXyWWxnUmP4
d7Pf/GFJJ6ZdlE+/nAmbJfbvEiu8nnbfVoq4UFL6LEIvpMFv7ItbWtjrQTbTUORKH3Z8ZQRpwEkK
kaeYcoK3FskbM0Qxy4tTWgLhhjZeHWa/xw1Q9TesBxbuocUia0ai44s08mrMurXYqIMf41+IyD2B
Xe2P11IxyeKtVz/mVE+GJbnofiRCjkHrJOskV1xpGCBJHAdHOyucVyVipCPWbK8yxvvs+Yj4wSwR
ZJxjFOv0yTJM0E6Cwj5Ca9Sbc/oDkWCNnR40KKpUd5+JnTRc4kG/ysy9vaaU+DE3Uk9JzewIEVDi
RWKcBnTiRuFCD3SVVsuN4s0dygh/XCyjXJYPie/uRsfNM05w3XhGOS2iymu9VGLc0k+VO2EZNAlV
iAdp5qWH9cWUrvEW9LaIrWkMS5SnZAqxw3JlJEefEs4FjpoCirBv7/og+9r0K4TeQP4U8Jl/E39f
9Rlo6dp8dnEDzqG+UKaUyqPKrWtPsawPE5hGHsiSOeVmXch15tlgkTfyZAfSLWVc74+Ly1sO+G2e
trp8aJntHxVhCNDmY+KtWJhHs5fbJdmdQPCOieRrPSjSr8UFgsvSKe232BbXYH3abqp/TF0jo3jD
Q9g32G2pMQvSRNRGRhianeHa46f9lRw5A+sVus9RcecflibcKKk+MFRsIkud+i0Lljz1Kw23Fg4J
p8HjX55PLbB8fnPJ0RhW2NJWM/KfSAeFil15hd1mEf3uL+3vTt5k/FgJJau96VYnz6IgN+S9L2r+
2K4JGn9HuZfSuYz1pjImfz28FJUg3zriWIvYYHuuGscb608lfKukEXiM6OlvY6Zzc7M4GLCCooGi
HKKc8AnrxN+FHHrQyTHka+xpor7F2mPt1BYCI8/BtFAVMM1iew5DYZOhC/GElxpk+Kef0wiBtms4
m4CLZy3xalPFEGbKy2JyL8XMh9zMu0E5meNiifbw0H6+LW+muIDenF9M5wzuoDYG7rZDHjeArmXK
e+31OVgDzok9ipDREUkXtJRUWqbT0qAKceFc8bRtEAXkfmdBNhyvHvSabDS4m0a2CVQPdPG8ZWkz
eKE5i0r+4E9e3/Cttooz6rR42kp3mB9l15J0fzxo50fV7n8Ngo59su4ziebyP5D7hpAIuupeEzA+
d9oBcsFbpBlQzsdpGkhXTlZcWka+bnrp0+syJP38931Xw74CA17ntq0VwfkQDbb6ZBPgyNOAYVmT
PAlgr4p1SvRtn9qzRgZc7ZUE8Do0rIPctU3mwN6tX3uJabemn1mGOVp4arJsGXve3PWE7IczmsKs
yR3cZvRTQFrgTBQ4YEZcA6fjAsxOAQBzKZq5TpBol05oaqGbchN7PQkejVqr3zUiWwDRjXVr243H
410jRhIIBd0VJg5aCTGtV7OdoPJ89EX24IgsJeToJPDQ5eTRzZdvhohmAAlAqqqS6H75XiaqnXVU
hJ83wkFUBGYjYNoKC0KM7sC2MNa6O28IGNpDEXRTK//72qxFsYN5A29LkM+ReErxm65iBSzN49a2
GZy7xt96j8Wr8n8PS6skKuEHF46SWdl2My9eZniels1iFnlK6a3U3cjBol7XJ9cBjDvxE12TD53y
pSuj4Qi5JsH8QXGneDg35t52eCrC5tmZogf7oMRohmxcJ9/9fA7hyVdzeeM+P6I03nLunjp1Q1vQ
4uVquVd0FECJNTvMNu3mmV0rUMWJcoOqBvNd0oWUD3R0VpSM+AvG/wbouzUDBh1vdWgqxZdbKME5
JdJBj7beneAfDOeDLRqf6ZWfb6FqvedvPPrkKv4CPmxE2Q2hYdhFK80qAnTHzLUgK5COlSsqkp5W
QAjQkSMpLeNBHKg+yLOUwJamdSjBTcwkcdeyKIDq5pfGkAJQx2K6zGYy4G+6zBhF3QfHVVx0mQQB
nujfBB0B7YTd2mvC0CSKRtCRN7fGj2T3TtPJlknfn2O977k4on88Zne9SKAWS1iq6SoxmkeVwBFl
r1pjDps+u/7Cefx7e8mCPyi07TuSMB8fa31teCdfu6HV/22cTA/yLbsAqPg0pIcvJ3JbU2RoQJEA
BkgvkCYVYwUHTGUBPI504MWZbp3d+kFwcSE6IUgwn5REig6/LUPeixrGEGFTnVZl58e+Kp0fLFsd
sGNEVvXxfJFW2H6JWPjW9/8s27g/dRbVCuZggyTfD0DuweaIJfNAz0vAiM228JNIavGd07LNNJy0
u8q4qOg1cX8rdjTW1mvMcBY0ArfkEfgQPAYObVDJdPBohzBxqKS+4a/Xlzi9rwH4ZtQo4kpkNjmJ
PkbmLaaffo3n0JTO2Ero8HIhotvpQNeqf3cEPrxpkBL9eguZAwLtS/I/bs3w/5iPqAPLynZ9FhxF
5/kuvCl/LvIfWFgDb+qeu8Ao59hc06iu03FgpFe4KYd8OqWqVhRZhugau5alLZu8g87kLogDtAqr
U14mkmC0Pp7GBMPmzQNxYKNqQ7Bmji1+ZYa6RhMFI0RUn+Kmp8MWPIZIoPcS1FfIjgt5dK8TxJiT
96ZesWt4JdAFhhcIwY0mjQH7GDlVhEP9R/jx3DZEONFZ1hbwnQvpV3r5WZuGQpyq+D3zT+7kw4yQ
n0eqVeVUkLK5AdofrmqTlqG8OznCetvZ0Ma6Yzl4zWowGDcX7EF3cTMRjyYMPc0kuqosX/PCnBxG
uJr0PDji2bVsdAesbSAvy50Ab0KKyVLnhI8mV/jpHVfuKZnIRyZ2loI9XkIkgIIwswyx9Mzf9Gm0
3VetRA1pEG+mnslE4XgVp5sfhijEuMGt3WVoFR6tkcJi8lcetEK2FBB3LUw08y+PxpKXOcJZj5kg
NsrvubxkuIGczus7UUuJcPI89sM9LUhPZLLH+FvhVrggFaEyUNDYoHNycBdLRsd+tm4xghE0tzLt
rX7JQIXnZFC1eAWmp1Nn0O+emQNrGUuI7Ngr7OKAdgcOwXUPm7L0dIQX5qHg0q8EsDSlr7CmLGiy
sKdYgQJCY4Ek09i06rlj8Jim1iMMn0m6v8/CTAQj6xaiZIi5CCEM5T2PB3HN2o2dJ+MZFu+k3mro
jT7oTTKnOlvivRXxyge9oOVsmCQ8gORPi9dy6JXhv1UE9E6XyQUz5Et63lpjyGne1wtIii3L2xsO
XoEcL8vX8olZU+/btrMZZE6uyjBRMpoqz9EUJB8j1D8++OEy8+sNnKmObELVNg+Cmz2VEq8nhnI3
4CXVBlOTqWXFDv+lmc1rlHaKBLXvMwmt3+mxcqNpDh24oJjFCvKaTtT0vcboQOfjA6mp4s+/IKnV
6Sn29X9cKTJby1m/IDQ4psEdBT2+AaOu8LWJJw3QTRisY/Y1Z0hMX9suvTPEWEQVWSdj65f5A50s
dnHa9iC4gYs0ApHTEX3l169gXNprsfEwqOck3Ew8Qlf+pDuuFAZSubUXwEDIabfHaOz2P5gLC83F
FG9yuIssJH8T0xMvP1zU8sP80CgVQudgH7oepIwgwSKcmSP06yMyZFz4TJ9W16/Nwwq0SVTUSRRe
9ertbti4OxgegSi1xUEyFXuVweP4QZBbsibrFlrdO2KpX2Mg4+DsOOzHGz8yYcW2XYJv2cmUZbvG
KRMk70p6FnevKY1Xe2v2fYJl9Tov/QlfNnnjMafvm73bk8Qpo2WBFn6uSc6tg5A5upFv6XX+nlUn
m/wwyeak3KlhSQnlBvvBZuD1txSzAH5XjoNEpD6bDSamjeMYZXHTB7leLK9rOs7OwVJ8S7l4yXzc
LeDZb58ui7O6rZXWFha7P6c/jjzWO1Kum0XZaDugfsIhOypI/8hW/UlebB95NCzPFTL2OfuF1gEI
DpRAwaNPMqIePhXRIcHqhpli0PG+iHQ870Uv6RMYTTwYR8DhCexYU/JXcltkG7sfHronCkvwri6K
Jl8T/5tRloE0Pfa0B9MRUUsJTyHsM4hP5qyXS/dOvyoI2hKkN1BCmaaPFmik8hC+LXBpiT4VbAxV
kwzXjHGNyDBJYm9DX/V6HNHc7rPHnhTzvcILbA6z1ynLyeHbFojlvaGDdzZC6RFSD+7j0gWoZR8X
tQHgvXyAb+E9BOcgHFp/UOj3gvAtRJo2lDgTjTzHwyzWJ5pNeB1Ow5d1S2jwNuqozBv11ib7vKxk
EJYzsHMMjeMwzAFHwDNhW1OW6ssDQcHm2BTnET6/27ngRWWplnm01+YyqggEdyVBIrHcb+i2iNR0
hfLgpwDk6eqvECokJWRHWRGRaWorlLexlzFwbBN7lOF7caxCrmci7pN69qKoyZR1lVWphrE30+lp
QxUCQmrDDjPG2qqcvUKI4ZUf9RNiF/nQGZfbtxInXogXb/Q/TkEErV8Vf4THstI476r3G5L7A1k6
tT8FCS0WPCzzBd4WRXA6tq2JBBdv1LB1xi/FocQdyeZk4Y1b/LweMuOasRL7m/ilYy8qoJp4u1P0
ldawDGzfviHPEYsA/oRTstgNif61zZ+Hs2nSirxLtrwja5vUGug2CeRcBXQ95scxpA+Vh9YHQJno
QxGM3T/cWtuobKrCAfe/uAk+5zpmgOky5stJT5wNRHGNc4VB+rqOIlyjH2y09mN0HnATUqH371FA
CgkrNKJAKrwAXrzn2ondYV4xdRSEUhc3tj1Fr06MBEPK6JZv7BFjab9DxfKW5DL9cFaXZjFiOkkk
GIWN8C+gfhU2MgetyOc3frmCsxhFbq34U863Kn6Rli8hshQvSA+BQ2pixsWva1QLpdlZWCORFuL1
RWoHV3tt37grFtcDfoLurv976vsOUAFRQvGc/ylDrzoreaq9/m9KycVRCyWugXFjb4yR8Pz6qrl7
2Tu/eB/VZuqbT9RzQCB1DuQOETBgJfS2J3xCPtBUQWgaZYFM4zWhCUECMQEnLaeBCbygZAcLWF0I
5I0bee8FI2v+KQ0R2NPCxgpz/CdipVwcza9tdHYRnlluFCHq3ft7eON3POgbFAzcouO5kicDpWlU
SXDbDjI/Le1AmnTHb37jAR72q4xwPe8KKAU+3hPvhwb/+VgzKgcL4cpWdJGYNI4GWi11hAtp+X0T
tPhaGWfk1o4inB9jlFOzCNWwHYrKwQKV+Xtw0splWpg9zzLFsYrhLjgTlf+rOf5vr3lyAVbzqOjv
3aEQfhXq1ynpiIo/e0JKHcjsHhnhciXSbDC/WSbILScsRs4V/L4nZ1JiCXGzwdg7xj5e47FWTj7T
PnXVVAlH5YESdzSBfiTrutmMAs+oOubEeW8xN8pq1+vZV1RM96uKCpWIfr8vUEgtfJIG38d/cNco
VIASGheObNqizb5/oOT4w40aWGGbr4W6faMU34dXh6GfcJbPFkTVMcAJcJOf3VSnEVHqlX7pqXOe
O+NKYQgrL5HLJz3mqbaEp6A/G8QnQAJl6kYgHfTZ9A3OIJJxOMTuGdXNf5P2MJp8TtCCwAJA9vpE
oJow5YIS6n2eJC93BnVjxNzuXiWYAVAD4z9P1csSAhdp+viXZ8twEjYQCYJbjxlGFDgdTUdKhGBL
uA61k+i52GNMoZIgKhmW/uBXF5kBbA7rM8bFNmEALEi0zcoDxvBBFJmjN2nx5reE/xO4thaoBi08
xvCAnsSmgv6HzMosnczVVJYTCrP/ZOGKtcv+uDNBtW16K5wW1rzLfwVSXrlVK8Y6w/J4NAo2kVYP
a7AJ56/JfDxcZLceIwws3l6OfuV23dlY2sTbzjzPcJAHmiLdtE0oXecfS8SMktGAP8E6PZDXLo/s
SHyrXb/uElemA+owwrLLGyx7aiSdMqVAceetjUYd+H09cgdRdWviMCzInBjQHysaUW1Qa5Cp4wnI
ImuWnhUsCO2whVVpdvW7hn5TWK1NZAPJA3zhc5wVyhcWp88PxY0CfgiVmtpKZ7c2FMrc6xVpbLIG
BpJXgoiJ6lDm9cpLFrhmpP0puD2AgJdI75BieagrUSxMNQkABg1ISnOEHopdns+epNCrDjIhEd/n
DH3zLHzcCi0xqTv+xUAGtmnCz+1p9aQcM9HZl9rtGj5ePTx3fZJ234zI8OeVKHv7s9OxQKjU5COR
oW+wimq3/ALqDervwrqWHGpxqlBQN/CpapT2ccQ5xjuBkrMTH/Ysu2bqHlcT5q6FdlrfFZe0VdSw
lkSdhSOqcTEQxIAwIsd+TQTU0aSgfwDg4X5j+5RsMlkqZQwJ8GvCkkAoxPJZAoap5P23KeXWAzAA
sRqKRmUhO1jQsGoQsCINIkTVlNMa+eiwgR+z/S+HlYIV0T9YmT1Ts5rQwvrZ0p0vyZukNXd19/8F
HvjsBV9Dm4EIVj3TC+QljEF2M9Rt2PVPZNCaTIZCygAJGAc/3/qeY58mSWIi+sO9f+4HQYAGf1zD
txV2gQRagliu8ehiMzxY0RPYW3dQWJMbw/5LoIbzec8oWFmDFOMk8eK9OAXcbx34xEXyHuuLJ3vi
n4nMnihPayzzopRW+sYv6mdC89LduI1gBgPaOoTIdoAQL/xCk9L8uzMeCJS4T2f9fJyZ0wDHg8CA
Ws3KWu199tO3GkOa7q4pqL35GaLB9t5BRKk1G+LQY3eofLNDQrv3waIilQgcQz/3zg2TWI03PQUH
XlICU1KE5mEMZlLHVqtImIF8523xwOvjRcCYE0XvgbvO0z03Gz/nocq66scojTzF4aj/HC20L5B3
1uKvqV2TxznUkGrbq47b+317ys9mkQyA0Ria+K4MKIkrym6jSEnnQ8fajqYnJFpS+mTW1/EqfEwA
sZKLxYx3tcNpw7T6nBdllyQb++6nkSzl7xWmW25FGKskGQfmG1V9jGaXo1Jgtf6eDUaF51+3/p/O
3rp9AmImyEX59xGLUrLg5D/2/7Z/UchvOzt8A3bcCjljRbMEAF7+8K9f7iyMT5jY3npuHCZEiR72
97ORK9J1hmZN5K/Qg9TRBQUFj/YiRs9ysUWjN0at8RlqxoWNYZniiKnER+lKgc87U3M+IM0hlJuH
lOOasJaldU6HC6D23BxMEuXnYwvsjq3VgEoCKF9twDPNTgN21GgwPtxzQNCpfTRkuO3YcQ1eXcvz
Rc/IIIMIJufItKZcjTwfWPSMaXFCTd2jzzW3OE0hPidspNgmEwZrAIQav0IWYSbMUH5IL9+2wxq3
7dOQ/kQpbdQaALB7CbOOofZiOLikc7ycl0x7sWFr+jj9Lrl3kdPbfzVmNmIQ/gS8ZG9qHOAd7EIl
CHkCAnEAJ3KM9Hx83VP/7skCR6+I+f8fRnFF3H8FA2iNBEClpK5WPpDBbjBLl/q/r7kPfTDaMfAn
a0MRDgDKpVq3WdmK4r2bFQp0NdA6Nkb90rJw9MpVt1hB6Vvj25rRD7tqmTRL3gP7oSwT3Rm7ORGH
5IhFfHNTAVHK2GcMsj2mLcusZ8aRIsmyzDwDzwVq0v+RREmuDAyY2on/RKNwSjjnWnBMyCpYwwZH
gvZz94zTtoaTmzRpAP9B/1lOx6gTCtGWouIBmjOXPwAY94GEeC+KK4KeA7PWY3pZrz7g86kkLJbV
vR45QieG1HdnKrP4TqkZX8HLz87DAgSck1/FtSFkum7pNQfgTXM2kdn4zc4+GmeMJ/16wtCA6LTF
8R/kUwH96C3EwD/kzciL8PRuKx9vVg+cQmhtEC+vzCeN9k2mQ8xapm5oHUcU33Z/yCOMHg6PbFjC
d4eXYodSluWUDMVIjWMKxf7ue1uax6IpiNxROEnsxze7cRv7c4GPBhqk72aaDqCryLqdyJuBwC0y
xG1wPqbLSuFG+VxQmtB+UdJ+JYYtcy0QQg9yFL2MArdRorKt18xQ+u82MiK3Q1CSySS/tc8kk/zv
8GpMeCqXPhzWW+SgD9TU3hjcf9o5Y+EAQugGQv6LTBOPQo30b88vcGytmLYFOdWe6vgen2KRA6Wm
98jKYtjd2ZBFPp2m/3Z+SiHrOjG+sl1d6O7vInPEZkAvCgx3muRcR5v2nJ3gDZyHO0cqWJG3venW
Sn87wRNvRzwM0rKEscapqurpCxYrBqJ2to8Ni/LI6H8uXg6tMpJzK2hN3ez9c/SMh+HntWdShSKV
/nXYsIU9Co2qE0hP7olUvvg/Vnw7nJ3UWhmvCoRCZDR4+DSwRNUJDQoNdnyJfS0vzcXAgmacMRHa
6C1uMBDvhI12Kyv7EoEiPEouWCcF1f6TTHM4NcLU3Ort97zbiv/TA7mHjOxKLUesq9n7JgEntdrg
cV54UiYhOqJKoXS8zJcE6eao32XId3sM6ZF9VoTq6WuKqRnYEebFGLvz3gAnxZwh4ve48F1ySLCm
9iAeFAMNBZp1qOrqvW+ezcIb1Gz9LURB02Fv3dSvx4UEyVDeRkKsJyDJo9+QtujF1hYK/6hTYope
gV5t0TLhAB0LE0d42xRx4mI5B1kYToquJS3LTzqJuamjkeLK5B1c/AemdZnHy/AkYDFa9jWQg4Ul
Mjx0XlZX6WrI94DdkIvE/KX+M1RARAev8uNy7eoC4OPcEzxmEV7APSqGPIf1VDBvkAo9c5XTWp+Z
0r4evhl8x/jkzmsE3Z7JdQBdIfzZ6wLsy9LG7nP82ffsyiO3RBRQ/MsNpvf5LLDtIy6t9hRZsnEH
nPqehqIxI4JN5UgoL/RJQofxZ2PT///s6X6MBSMZL8bsRlzv53OzOWJG/p3/vLWoqJ54mnAa3Atf
8AwuJhRuUE2Eog+fsYhheV6bFjHI3Rl/kXvjMtTZYjeCUT7aN+i3lacDms+tYHppHZLvOGwSAyHh
PqxB01ccoeg3fXld/A6Fd4LDis9cUmxOmZZxkwe0fzQW2BkVZ1lup9h4Bh06mNdFLYgjTCmz7gff
uFSyf4n8QWZ5nexMtKaR6kEDdrvK2ZBVXmP43BfsWbQ8p2LEiXWMymm5eplHHxPSVOUbDc7ghndl
9Eyd3+b9eFyVU9pdPPYJ/OtrAJKcHGPvhhRoPsyASdfZl+WQDktFx22EXABj29hmVVvUX/BuVUYw
4fryqvQaI6g1OvMRfyfq/YR9DzpjDwmSTmHo4lHBD7ZfnsZ0HS6085/SdpV6n8wMQ1NOYJv3F4EF
+pqttnISMVqZvevEF6A2O78O1PjUh/9PdcnDUTWZA92bJWmnTIfEXA4fcpuMenTMgQ1kies8enDU
ej4BWYY4Fi9u3rGLIf2r0hbKH86DFFxqqV5d4zwS2SayNqRgfBzPXjjNHTjtGtYs9s6T49RFAevO
jZoVeYYmkh9kHw3pLYw8Ax0uF3a3V2LugjXiCtbZM9vWN1rN7h0H3pyH5fb8Z1Q1Yf7k0D9sODfn
nCvXrVhQQ3WnkwcPiNgANwcX+0LRBrqmLWYEkvxq6uPjB+BVxfaLhV9JWsXagLIwyNJYzXHs8Wkx
G5vy2qW39p1jGHkJfo0+nSnvi/C6n2S04xraf2jf1w4a2/EQbYkv2ejVKnUay/Vv8hhj+dUzB6fz
4pAvMHYEzu3flG5wpJSF49x87td+kOM6gTJau9rBk/KOgEU8+ZRi5iC/TJtF9KQbBl49QeTiHx5a
zLItz0AvMLPwrECJ6qgyJtpe0vOYDd1hmmjlomUTvZUiMh7nQk0rBzh0Ru16p12MokH96/uGcTz2
xQVnXk/rbsd5hFUp30++KMvZoPHvy+kiR217J9CiJppcPMjwzLS0hzE4fY3xQaEpGvJJ3VWmZzY7
JmYfC728SBn4LUxd6zgelNK7+w2hXZG4JfvNHbQwDUtD/nlRUpMEmDZsGzWZWr8iCfjpWng6Rfum
r+MgSDmhdXq51TxepWMeKepdij0Qd6hKEy6FQVS0yFcRPY3AnI7Is+zxff9a4Pf7w9kiUJLzy6tJ
ufgwj/etWq4TJnuEU28XC7Ms01l+eZ6BtJSoA7ObUup4E/TM7LMftVTBjy4zH51yj9p8uoPTdoLu
viTPpSUNIETXIqL02TAU4/EyvexOr1/Y4EcqPohvPx38AOyihQ79rbfwwucb3asHUO6DO7gnJVI6
MsCkfM6XF8lfWzEz9PB/Q/ECzY44LpoGPFrnzya7SSv00bAdKNrrtCU/cpQ5XtmlV+O6/W5E3PUK
1GoM1xUXxc+KbPc1kzPLYezUQ1Zq2W5bDGI0SpX3hxTwGI6F3tQjnZd7CL/j8jgFLqTCtRLOFfZr
+eJ4YsxcWvfKIH8Za8p1GSET9Yr98DkoLD6BCp9bX30bkpONZ+NAWmdXr6Pdh7GJ9w6jIeKxdxhg
yFSg2yeY8epWJnz6uY8cBFrNSUg1iiA1D6pTSbE2aYeDGHKk/SN8bSC7VqwaKZ4KcaoBarHtyi9g
JC64CSOKGDRIMPmi+yZ+hrSC8ceMiUAlmmwDMRYOTB7kDkbDqzhNkf9EyFE9V/zhNnd3EoNg9mxN
vBPhGjhnN620/jiu0qUETS7oR+wlIvPKPyQqRePRg2Fy6+IkbwxYmNEQu6eBVaqVFfZBz+98L1tg
Uyk4a3R7nENAheqS7iJOgkD46/r62pSGOk+bsFYj7AU3hqjww6SimTBCRxR9GPj13t0E4zU8XNMA
VnKJd17fwD8k5j6otYaodNFZdx84k0cekrditePpF/Y6YuVVv9Xv5KZNX/pwxI6gKXPdJ1zDdPIs
q7kt2DVEzPgdbSdGjA20XHyRXEF5fRUNvnIsbfbcWZI/JpmP/HbZWKjAmli2M98gP8GcHMzAzoKj
pPEeFSetXu/Zl36htyBOgwmRG5kz4DrZtkZQDHRKn4K2iCWMhIwDWY8Gc0Uau4+fAN6LD1wFwn1p
kM6njgvOpkE6kRGBXy3l1iyThF+Hq8mJvsXlLCJu069078BGDfnRdM4zDBFAZR/aRp814NKsQiA3
gNtiljJ2QyCym6SoThvyjaG6T2LxCXxSDUYJ15DXwPOMbw6h/28N3/DsJjqw7Lq3V70Moh0oiiEo
ohqu3xWXQKU9zZ+YbqzD2m6mxGFYidnJiyQZodMFfDJz84DDxIxYbNqIiGSEelNoK3bYn7zyW7no
qOfhfxvJ2PcQTx2fQJ3mJJ+eXAtlH4i/zMNFhxk+3PkvEP2EK7bZbKnXOdSjASo547fkTHpcPVU6
oEL3OX+wN6ZOij3fWNsa5cgM6KpIYtlwhzvkOTkJCLa/cGehxMKo3pP8ibcxe+HJTpR5PM1dDa6A
BfhFgA2zAmnZtYSSJ33bssSwOTnhNCbfx0ZkYcz7cQn4Q1r9NzFEU0gRXndHg73E99Sv+wp7wmis
yorKg/5jUq8KWmIyx7OyDQntzaoIkSVNLPj4dIG3sVhiPO9drvc5rhgkh7ShhuZik5cOuEjsnQjW
WbkLQcRABQtdJZXPWx3euTdCKG+0m4BdgDxCI5X9mLc9OdB8UcxhLSWRB6FGL2Bnp1/UBi5rSo6i
rfAKmZDBE1J5A5ka7gSgblsILnsYVpbRoLsCJaGEeyNIlIslF6tunTnI2labBp8S2sU2A6WgnVQk
8bw1KX6mxdgrAEwuMPDHBUsSiBccZcQ9nOfMg8j64aBf7xoRVtkgQ/xymvbrlPRaV6A2IXq4CKoy
Wo2wu+pjCYUysV4R2ghIE1pm0vWv0Nv/oFRFdqA5EOUplWaQsD9gDJ2qKJG5X9Uba8Y7B63fZVsp
4UqaPfe5c8j3Rr1BU0MnTHAOHeyHP3UzWqPcgHmE3hGRmByya+U8Rmce0uz4UQgTjkikpbIAx1Is
AcTZr3fvt3PPMV8ei1QsVzK5kdHwa+9xI4KOT662Rty4lCDJyk6D5xT0XGqS/id+l/JHBCIxC6EL
MCJUTbDBQTTI6NpvW/S5bLh7sGpV9riLTpbx3kHnFC71sOAWFVrxP5pEGyF2XQws2+jSyfXj+m1Y
u7E3iloW9JY6sYCuOpXxPTjM0BaGOtD/rOmk6D+dG2nRuZ8igXDyzmL6OKMepC4IeBXFXYfQ5KAo
QVkIEmcKljelizIBDGM2Xvl+syWD2NYrNFSXmcnCWEZIYG/4t5MivTvScT4XtzawYhaQ2IUtXeFc
ov9zHR3wazuSkJ3YlbqPxN8nWTbpeKRjX4vangoLd/DUqFJBMwToSua8yylBHBqPXlcyTXx12W/I
YnfXcZghojE8IVVFHZZMjEwAo+HOjbGpNfNw/RaY3sZ55Rx1YFr34bcSA7rXxZI3jqTr6RoEcDNh
8QOuF2jB6LNmOuHgHxTwmmEI9kIn2CuXxiUJJzHiy+e49sKj4qCkb1f8peSOVodGQwhS3KXsxDS9
TNXu+VoIKfJrlqaV6l432CxrEj1eBnftDcL+bs9wiIF0w2vt4YDPYQyYvfUhDu+/hZTu3mexeh9p
ZGscYcEjERiDo/IkH+yJ6vtI0YjckuJg/fXSB3aXwGF9d59kCELq0RrXNXwBTPWfvk47n1/+7I2F
k8vh6kkccLdjXm470EXS/xxb+9FOUjG9q24n6fA5yXDIx/lVcsvSxzvc++auo92inPZMUjkBGGQ9
NZM5SrA+cIR89eP+HX7Mq9GjQqXffejllwpsveT4e0VFxoh3V1Vup+zZNhJFWkEvJxr5Ti8OOPFq
yIgJYmHHekz5vzT5qgiDVDbQ1KJqjHZdbPkP0HeDqJAnqZApFKyx/l5zgNw7xQ1/26yWDREYq6z/
saHW3QzzxKRRLorkFNIr/mEbjIbwRsfQCi0gNY41QqMpELPyi2GDKoS8N34ZIic+yDJNjF7vxlGT
n/ugv8t/+VWnbfV+T68WMsjGflR/tDilVZRKSlyfLSBYzRUG7Mr1FRkHAjxQ7/54FUviKMd+OI31
IYFFAre9JYpEDzwILRyBcnm4mx6eWs8u8LEW+82h2Fco72roOy/RseKjSKjhEWUxZq1k83tQctym
/5rHpzOTYLISNv3GvkNemnxxmRH2fhYfTGGd8bgSg/Vt9HBYQ+Ci7RlOg8mmhNtHU1pHRwRPZVPQ
vjL7ZYbY/R2AZvHW8c7eXlHvoQvOEKfJzTeukOaCcFO4XLbbbGdSY8z5a+EdGcwXNJm4rMIJI5cP
15kqzIugpM1HwJGwN4FxUbTp7Ym46S/h0tSwLL5wA4tAzeqWyFzDR6xoM0fmGq43V54qx8+TfpbB
rrrECJwwAzF9CvQhmJksJXg/UyIxddUIiBVNTKsMtWH8DZc8cG6jmOojOj79u4n0ymnaDRfe5hPk
g0N9f742SD3lS/FbdMe90tXDMtLKs8a0rkLJRgZAOT6q0EgANjQtsiF5UlRtdnmxe3F6F3WzplFt
XkRjClf5go78ikVqqjithXLINaWEe+rv0/AY/fbBeAWDnM9JxQ3aRZ4MH/Ld2Rw0gGnh6OnyYYUW
CAaz8qTEeonhczqbVjD4MEzdfJ2IKtdZ5BB6UDyYwh+nf8M0ztc6wwil4zJSbPP5Tg5R8KVrrxmm
zB3WmZh9jvcORXuiPq8nBtwv31ukKneC1VkAEOn1trx7yqgYA49MzKCDgfh/CmkQwKk89YYm5Qrp
zCZET43iyh7kLgPJe88/wi4eCljJIg+wIhBwSd68ZBm/ySov+uxSB+IFGVtamCD3BWsR5LBgIbrK
pukveWOXnwhG5hO6XRXR1Voo5ymv8eSCLOAnTKl84LDk2hLPGa9BS/pv39wj+g48+0kn0zFIhpyQ
EjvrCq+i/GKRQhQfQulWOO/rVtfM0zOAPW02DCk/MpYNClm/5/txjNFdoSzztpRZVpzx8bPf6Pm+
hnvfuOpER3lfmf9VYQEpojQ6T22Dx5J4o9eFqeGYOJ0IshBdAniV7ynbzcdRyC60EBZl54F8lFO7
ZHz80KG+TQMy94xins2CVi5YLJuI8i0S1KrvLjH0+xNJO/ZFx0vwZKuiJVjxQJytBkqmAL2EgPv+
a3krpNqijB50GTVqMlPY+OvXBRVoqq4X3gkLw5JfON89h/P/jda2bEcIkU7fSgQ8eah88UUqRNTX
ylLAStdkWnHa/yU5ZmCCsl7DBnwmZxhh5M0xg28mGRwJxnfy26KOk94WXfdP+Ygjo/ItmOCYp6DO
fcLKgoOKSHq/6R1Pn/lTBl8ZlQ+Xla9OgFzjkWOOFEIewOpcZuShF/POtpU3eZ/OAcnfMIQ8C6cO
CAAgYmqEygPkVphgc+YLTYEuEpWq3Exr+rcK6adu3/TuDYd0XxBOr0LUjDa0GAD2ev3kLFfiPORf
mrXLs30JBv23pGEzUx7yq4y1ARCP4NcAkmo3kXQa/tt16imaiga1FaYbc/3nzOprYkCzBfATC4iP
MEadnEfo9k5h2hbhLpFDRslUcIKMrq3MdtPBPb2BpW+EzWgDYF9DuXw/pZ9c1OuTYOzmVqNRuudy
skNHTsH4uSZzGPumdI+iihrM3dik9A/FCc+4zkxPoGK0ZvXLIoYDixImqv9OZP8qB43rYkIa0pbL
nUQXGZkC2U9tKfaTQbW7NWZ/SkPnUhGGcTRFG5RfdCjkX+tooTjHS8DzAxjPFreH35VFSmvId6EO
Hwc5eM8D++EAM6rZDMVUlB7p/Dej73GScdAD4Ld8jSQeRlZO3qGtys8PBVsLxCnfgklMJYLd6YmS
R0FAhuLT6N0eLgzicFGiia0FwanmG882ck37VTAixkJ/kY+I5ifSz49jrcPCv6z8k4d65NdvACxx
F31S6q/dq/Ysq1FgObwTm2ioz/xbA7a/2nZKaajOkLHgtD8KK7CumY5V0xJCmcseGAq6zrTtVQws
WzCPlVqdGYLQeGPb87ECpsVZ2n+lCpEz+C1c2cHEzeyjLsIRTBbiBNJ3NHUO3WwB6eTO+ShxTvu6
jHe+EP62iTTVSZ/Jo7dB5NClkkey32bAItPLHerRxqCyGYimKgJ3wVtfxyKVKVl7uKySfZ8pEbZZ
42voYY9nH2m39noU8c9rBq9BaQE4E7nHLd5FawYB8x0OzRa1VVLwobb47RPnxgQOWC9eLWh+Rq5q
rQLo6JqPXjAlmzaH51CW6++fct/hBmI6wjl5Mam2frIChflM77XV3u+4tCxhKlCc7IrefE7JivRW
4MTN1w0cXNH3jMb+tu9N4JmYGulLzoOzreWVD4fMNLuHQchdYR7TXc6pkselEI2qULj5dQLvcXEZ
UxWwB0FmG72p3ilviO/SyETednLjzDOGMlrU3CUD97p6h1Tg3KQEMsMepKRDzRnh4Bf71EgTlELA
HbskdCWtyJFFSwMhOAjuBGvO5eULFeuvcVJYeu7CF0OQozXcMkHSs4Caw0mmRQ33v9y0h+2KDold
Uma4S/O4YUDVJYQK2hnLmtyB/rjuPuRNoStqE/H7nwrLENdXHOgnTjMqZJiLSMiYwGzuX+Eyp4vq
g/feAR4EUwgL3VR2LIkAaTpJ1oh0DVULL3OB9YpC6OLcLDiXV5ITmqNLiOyzonLbdjDqYEwg89s3
sEVuFtOOUKvjxMqbTZdp9ELd8H3LUKYl59SOVoTHh1lsIEOIRv9a14UXP6eJ1cb4w84KxOFiOgtL
SB04zHGHuKDqQbiY8TN6YbZ9/2Ch2GTCfI/nBRXS8B60dWpUcETzvLY3llujzLGdwdxqkmeqgrL6
bLYA7rH2AcojeQK/6S7XckPwXkAzCirLwEtewhQBMqS+LEfPHsj6uuVMTxKYNZQlD4pkZQ4JWWNf
OUkVHhf10dyzgL1wJYNbo/2RIYHEdXxj/IZLqvx1wt2xAWOLXXtCzrgKgmbfiuc9yAAHB40PNd88
DgdIvZmcylBeHhNesvUL/DkZu0AechEdnj6xLzT2bvdTgcYB6TmX84rEyYuVz/Ahd1Zdi8az+VSP
IZ9R7SJJJRE69GG7AOHZt4lcSwIf/vuhTaEpEe2OHSfuzQ3AKqQGYHFwWKYU6QgFq76/PELajPNW
frTGoQl9do8zXRgyy214OCaNyFOl6XIID08zZTHByN64qoCGynkxLZaZyo+71otxW7Mvx9Fnzj2n
OUenUJ9JeotVEceQ/O/sK9WEQRyd6jGrFTC7jEvF2Il5YVsmWtuTWgi7ahIZfKFJc7qcFyTI3pZS
E1kLWN46cgqOGcikLls9H+F9hi6U3V6y5TlxtgAsiGjIFOzz3Nx303dV/p9NhyKMApSl73ZbNLkb
xkqiCnSVYApUMoaeID9dL6lU0ZnAahBDwHLyfHPpOk7zI7/85WFVSe5v2SDRB7e37SWCQJwTdOJz
HXaojikNURsKS0A2208DoNMZ9MDaZFod9m+7CGyEh0Xuh2OphCzO5JoY0K4Oa8Wk/Uc3t9cmUtph
3CfhvR7m7RgjTNO4h5QAqGScrop8zzgsV2dyW2fSHeflJFzoEvlyrPo+FSEC+aqgBIIJT79DmJkX
8KbnMs3liKQX/q03tcvNs2hJy6rMU0QvqWOcIMj3x1Ri8qbA0bVK8jbm3OexhFtA10BjVkvDojbp
3UaJOnsw/FwzfHHLXWjoqZCSQ2o6/nn7+IRrDoPHxf+i4mrVi5yr3/71uH4CIl0jmecDIY+EknK+
+NxaNdoqhavVFSBHVkCp2bjV332opx2SxqX2zSsvYmstnlALrGDQRs1AF5oGxCS18hbOKiZk8P8U
T4wBgp02jGE7La0wLI9ut5GkM2km8PwJ3nQVWDEpx1NA16Wt/+5tx3puXdZ21FT7BWNoaD0UPin5
blcvaic5rIhRe1YI/bV4PY0Ns76jZB1+QsZNRKwdp2ktfvDxk6/4+6lJtNInYPf9vw7Yg+xi/OrC
n3I8QuXSEGgpBSTjbM4yJKWtMo9ONpYesFdvqBwsb8/qdb3Yscydx5XlmOdnQjxYZ0epu/xgBZ9S
F0TmApiD3webvNNAVAFjLD6N3ywus5F16fRqeuilqKYWLMDw7gcwWNTOVgHAHGZ1Oj5sR+OiL//R
HGT/HFYj9vWCc1Fgj/7+33ao/rp2vvBcv0uVfEMWdif+WbpfJXpqWlwRr+/1wKIHiOq/QnoEVZtk
ZOl3avlxYrkqNaRs25eJN+spEOC6HaJQKEIm/bxWZmDd7GhxVQ9o8c06tNyROB6e8OaTb5jkUJ3S
NX8D0njYcLpixPUlxdl2MW1YkFBMNvzmhoB83aPnHZOZiotbJHtEZEaZJ//mTD3Q3bvxT8ilr7Xk
+1P4JCfGR+/9FhG0Ga1o0SQBqAWxz2CT+Hr4p2btomhDx3JvUF7+cXl6bEuhRHumxZsf9G6Ung/x
tXxLD6WyiiMWEaXpRWogwop1AjDE3dXTgqn7EartRcr9kX+ub/UzDDTi/HeAeHYKffxHK4ST/TWE
DSMyvW9vWYLliudgcjjCXnR4P+lw6/FfDRZqRMXNG8sMINywdSdW1lX9ElM+pAsDWH0me6d/G1KR
rymfft+z0euz54HyppkW8VaPSpHLnhyMkq/AL1vhMgkLn1WdJdiF98TXf2e8b2p04l8IjjQoxMly
a1O4EbZ8mE2hX8WIPdItuFc/XZ/wGkXTfBJLxg5S+wyAiw5/8eUnGLOKsBAIy/zCsDkY+cCAAtGR
NLIwM6AN074JZRo2PbBzB4H+H9zjHZY18EQuHtrJCv978YhZyRh77lTWfOXlbzLork+Ea31AXIZy
5SD6O/Wx7Ns2IvEM9bKDNOWG5F+w1gKCxnQ1PmybSmQWq55QeWKGJCjZ0RlhjTiRrlpp6MD3EUIo
aLz1hE9pwJTFgD4+VHd91ZScYaeyhXRfa2NpWSthnVvzNVKY1AvZbxViNLadBcc+5fFFHnceaFKe
AfrZ3T/uYQjG0X7RTi+iIlhNKjv1dhxPfwY0hkBFZRJJtQtULBTGGjTp5PUgn9FL0hKQjYFaYk8e
elpjDF8lEqIDhz7WSG5TwnWpXGcPD74mxaVfHVNI7nRdG6827uqu+06MtFn62A1ko0xwA5sC8KWu
0P4287wcAm14al8vd5q4JMt3OuiDSTIScIZaQIaPMP1/pIwg1zJgAm70V36CqkHJfF+9E0f6TT64
i6lsEDPKctxLinUCwCQIEhaZE7X8Xain5QVtzj0G9SbiW9fd9CCGm14JpI8LIzNW6ekgfAWtsL/h
IEUm3qiGI41jbEkTvP3pm0wdTsB0boiwBNclSRiuoVbu6uCF/ZorcDK8dapoVk50JIO8OTFa2oNZ
iaESyYznLhHVTA57bkfOJk6mlm107kHFBk8xbYscMEk2s2NuMMuaXVAMzJovZlJBNaDI5hESLhYB
i6ap3fkwYq0VQERakx+OKBkukZNihL8lqkUUFuVJ5IbMgfh9tUR9cuYFw+SpFVyLARYQSNLcgHHz
VWzqvrQq6vCe9E4KVZLnp5yVpsAEbuYAKlE5Ez/MzzqA+GFUMq3FJ3iT/YPZonohzJZRUOtW77Ou
bjtCrsO/dsnK6UbzENdjW8ecq4gYNwZg2SVXv7us4yl26eYhhQLhyQeJqiIYuy+QuvPD0jwPvHdj
QMJSjSYNiVUhKmUGBzmYBTLTl15AM1VZ3MjnUoy4mIkTXNoJS3jElIuzvJvUwKlSeCeoPcqV3rUP
qO4++LnF0ix/wdJ38kb2lGc2KhY9K0kYeymMFzPPYzZdsT87oUFUVGmxi6YYF2j9x4rHzKAvlJrc
IHRbMuYKRqNn4G5nOClE8Hmq+WkfEuYkWmby0JU+9BwRP2IJmUdcbg1FGIYJakLnqqNOezA6+Mo7
QUlk02uErPAp9mZ4MQD2gr6bX8v09MVs+kV2q9lgGZMVDoHpE+pC0jod4yfawCN501/Li5T8ivte
kOGw1nTY2JAOyD6luUzU3W/C68zb3hm26ProxgHVs8VxK7aqlUNnX0NCsgpBHHfg2TNmBBXLao9o
AUuzqCOCNPevgO8HyM+nA8Udd0sYDNLn6mZm7X4/dC5l/cywsPYsWx0cKrhxBQelrKl75Pgi7loy
rl2gPZWEaKs9OYAs6roqWU+SWqFVYyDRiXgpugwcmge+WvOq5O+JjHxhQBS0XR7QyYfGnBY/1tRN
1zvllQbdxYBGT7Xk+y1tLFBLT9CWDOIrHgrP0oib1sbgWAkf1p7Ln8c0xJk4CrnA7WGUcSoSE3yZ
8obzsfKLPj3aJl8wM5jGMvaHm1lY9lEWca/axMww8D7cbPG90ILsrcGuvbyLcI+SI/bI8L5h8FUd
hBGJjE/+MXc5eEFWNf0gDU6IrVhS6DEsuMPDpKZZfdXstwDZcHuc5wxlzmopwY/g5i+qzL8N1bVA
NVUxaaOeCo40mfAaLiGqYokrxQUrPOh6iHm82m3SuY0PUU582G7fjmCLoffc746P8O027w9GzmRz
y8cV0AqE/fA9MgIxqnWnTlOHc5sAA0vRo5s7Ka0RAys0r7FDPs2wDpi10ywW9kl3FqKbblW2MIlV
4uV9zHEUlKGcKhxn/m3NPN2mVFA1exqvTJwMP+EsmU5ZfUcn9Al43RLH0Kn/s+G+ro1Vdr2N3XK1
5f1gguVLsb90QKfCPPugagHnrHV3YeojRcaTWUDHlsG/UPvfGQKrwmaOGbRB9QZ6Qxt1iJ8F0629
2Of9nsms4Tju1gpUfUmcxF6ZYV6B08EQsh0AeCTHpj/f4b/lNYV/7/9CIIvR3eEfNOq8WZtK9hm7
eYWS/0f89ZtN5C8AjZVQuM8NVQRoYUVtBn/Ql0d1DmVgOxOwwhlC/BUuRdTTGv4I5u/a5m5zvDG7
OzBbQCOCQV1LQe4/AZ4ZTljLrNfOLm8vfJ4m5kcCDsHcu6rdohlZ5u01V69znaN5oAXCWmUjOJtF
byGhBeMtLJ6ft5tJDaKObtV1PBRkZTBNey7tmv8BSm1onlaI+fMAIB41P6z4YkktEXegiso92xKx
YbgFr1GhKazZDTQn5fKXBlZftpsT0+pdpsvN84U4IAkHvdiDQ4wWrSGC9dmq7/t29bIuvabdYU4B
k1VB3wB4WA4pigPiAgDOd3FGOQbJl/hA3jqybvOfLvBo0043/7n4nqM1bnaTRfallBDbO/UODnG8
6GSD6MmCaA+XzYDMkxLuP4fhT2JexMAi/RQPi2iGkoMY2LDD5e9FQrH4B3it3fNAB9k0+lzbJGBP
oOK9qL2I7j4HMgMKyL9yS6NYpH/oXtVpW7cdvr8bBHqWw+WQwzlOCZcPLFTK3qh1nJChpgR9U7o5
r4Gh4+1zuYvUYpU6DVaFNHOmPrFrb9c0RPmbqcW9UKFr61DSoQv+ZfvjM8Y4G02JcAx6mu+KRyYq
JdZGdtjTbLk6c7BN1IBEJ6zTlmnqY/BQyo6R844JqvHnjIPt19VO6AbHpFs0qDjTcHhhlJm/tHc3
EOolOEmbKf+iPglTSURYsGokJFMfX801DOt8KE1YGYycjOv/BPwdZrA1p1TbLJA90EyfoAMTJXMM
M5/oSoBoQ/4v35HYaBbZUlXBYs5aojK4JmExS/VsbzW1Vpk2jQdLAZCRlAlBnSl7Ihxe1QpvuMIe
Z9MkYSpupbDKQTOZ5HlwQW/NQYXcRch5YPwQHqSe3NpwarM9IE68wzLaS62Y3GhRBqwTy3qlau1z
X7sIvJQnmVoZhSZXW9sVppDd/7fDUMOvtg9kvzkffa3Qbf6go9Oe0vdPi9su/nJC44CscQ/3miWd
fKpV4DYomVPfQuTcDZIFW2WyZKB6AzlkAx4Xmhl6j7LgYaNmpEQSKcBuWNC5CWcdgaIJiqR0yhI9
eG8Xc/q2y/U0oozOlakxArYpDPeTYNLm55/FlNOO63keRBKjGJ/1XQmRY1SnVJCOBV2KzcW1fHB/
72DXkM3vS5854tR03qRe+HauFDPqgRq1hVnXCS35oI88BJkt6Dxic3fH4ST1vcLNpZXfjM3dSR+v
JyeRiNCBVC1zWomIwghdq8NQhaugInehHCEKc8DyiwOTsX84JyGqO0ylvNZg2uMmSxM1j7z29Izv
HUWFrcd5CWxp+QHLdD5y0hC3p4dn1/pOnq7kwqHi7BEwff/YZOajLZxRqmoG+UVXlWIyw2H3B57z
oi604J7gPgJ+i1z3ELZm3fwVow2S7CCabdL7aKn0AhT0zQii5B/GW9GK0cRIiA6yqKR233OA/zBa
RMmBcIMk+PZz8XUbUmrgEHkJIBh0kHGeQ9+zxxniGSCk6VSqcpxORCw0mwhrJ157maKu1704EyHo
H2qj/dGoS+IYiOU6WNES4IUGtAVZs0S18+QZ0sWCCYRsEcsNG5iRkNSBWcF17I4CAdIEjQAYXuft
IOAmfXnvqaxQLnBWyd1P1lCvqdHUVuYE6rtlKDmUhxZOYi9cXoKZqzVG7aaS5YSOxgOhoQ3ftTo/
vfcV0+y0JYwwXtDGOjWkmtZbvrc309o3mLAuquZLQ3QTG7Jo2NjdBlaP2m/1NXSVI0+bp8FKVaJD
ZH5dNdGESIxIy3s4tiNEc8ZHzGYh6x0F2U70Z6yC5l8bs94OgtfGUtxRBzPDe/rB0CIvztNDcRlO
lY6vJ9+Z+BNor2S6YPiMprWbWP6JTU/PW8vWWLtG7qY9yjiFrnIDDSyAMiz0axsQqGfiixAQ0PEM
TiQL81B+ZXcCP3sQORWST+GoJtXL4z8bdJlHaBOm98b6ul1NbOvH5ZUtp36pD7bRy8ZAEby13MmW
RV7iT7FhgarTcXtv9XSwNBDWgxDr0CluWHhFyLi7d+VZK/yg0Y/EDiSsL9O+/P2l9Re1J4FL0Dos
9cPy1CkmURk+6llkYNKyu20BKbUcODeZMiNOhrEDbHCpgOazSTjbIeulrke4z7/HbNTaqIBPOhFC
tJ6vcUb5VCfzCGc7on0X9VXU7/6BY3XaENq9S4nECgb7IrJGEGJBAkI1JDXu/qLY8R8tnWdcz1Fe
5L0p8iiztK3bsQJjl5FM9qhw1YiHSTFgkktHBPz46fdjhgzhqc0Y57qS9sIyYHbSxKh57E8Y9NW/
fWuvvXAdVHB9qsj/ttdzEq9Vw/Kan/50Qxtm7lo40yrqmLCOzPEmQ6Jjv2eV5cWuRNV6CdxJ4z57
oUksDORRCuyzByYtiEd3GONd4vQmFV0J0hVhF0UUAnUHrY2kDO4A/Rt8gclowuW3t6VZIrj0xOSR
xOB2WjSLaRrsLel7hzeVtZVr9qOu/o7yZVeXgJzCpNLypx7HqZ/+MyYB/HO6NUFppSeIQyz7Wj8T
nbpWf9w9m+/EtwRIdppoAEygsLz28I0mM7otJc9gfwfuINIX69aPomLH6A02rug1SQ1lCSqf3647
WzldcO7D2x1CU9RgnrcDKo+iTcsqtsm5y68abZkwaAGa/32egB89HO93Q8za3tnBtMVSSwlhfng4
ljeFQpA4YIH3N/ZnZEV3o1ZmWOnQZOHbgfF+WZNcczntSA5FBx5MD3CbS5yU1jAY7RNiU5oz8Ryb
soVyXFvxn2GyEL56L4184gQDXjAe6ih9sj5YmWx+6+0FgjbooLUQCff/sbqC/UmR82YttrHSMgAY
T0briHoHO4bZX8l6PGLJMgbcvFyhvgt7eFt8TwavKFI4Jil+z07NHoqhpCJovGgm91LY77mc57f0
3tExf4KPG00nsUoemxVQhWVzBqPMD7Xh8mm0aEeFrI6HKKv8MkCd68SOKgxme4jCikwLm1cqu7DG
PjhOVxS2Y4Najev9VlxZBj4APFT7bhZ6jVvCMCqWdu2rKs46pVPl/eNN2fxLP+LariHalLaZJMHd
BbnW5JiBh6JyieHV48q7qNzfUPbK/X5Erxe0mN4z3fck9mDA0V9CcZUkSMSoP1D+noqGSZnuxtC0
e9TtlXFh/qBi9AeQvPnsEbrq5lS0LWUX/ZRfgmVPa3lh9CSXPONRKno0UyPXiTtVvrqn5OFS9UY7
nXUzwWtKR/NWWiHDSMrzE1/OrFL3iECf0E2YQ9CD44i8bhztEdSidJBVu93Q80F0sahNYN9Fo5/r
aRutjqItRXo9Ml4ymrJmAkau6F0am7+gK84SO3/bQl49GekNhRGcoTq244C5jtCYRx0+ATY8jwEZ
Ycjnwzn80jXTNwxcv83mT0UYtDgS4mEq9YFYgYsg7TPpEsJAz7NyuguL8e0RB5L5GdRRlmxZMuuj
G+8GM9OAI5rtxiYOM6x+6Bnm9lRxG5lOyGBYhfK/xDuPlzcvxJbJTmyG/t1T5wWC3Mckmdt77IE6
d/k+mLmB7uytrCPrSUJEkW2ir/YKhft9+hqAK0L1lFyS2fmeSrUZyx5GmkBBuMkdsxlvpO/cTzJR
Jx1uky4cj8LxT1ZHEDsnHKSNFvMbcoZ81VIHA6o9+UanO4lvDwujn5IQLdx4AG9nUoO97vcylvpi
tLsYaqOCUipYyOgi+VoqGq9CU6ZwlvcIrOpFQbjmWTkoOscaT0TvXrMNKMC05XME/SJkuLIrWKSd
rf1D3gvbglhROqINOGW494g+AZIeUwNa4/thTXAdEucH8cqg3Jb65qi5vIiFCmVGJqR+ViLmNl4l
mv7bqSjFBZp6Rtsq1RXh5A1cXsu7DBOE4T92nO9C+y+s/kMDG5vdKZKePq8ptqc6LMsqlq69XMZP
+JD3DGnXSGz4+OLA67FcSUGrf9v2b+3C5upRTPPDinB+gmbm74vOaGFTxpF+28FSkYu5Ovrv35PV
un9icQIEcu108L3Yv9rTUjjPjGJhy+aqVQ0s9wAjMWuv6CoQeDxnjoHVtqc2upRSyaGp5aV6nshV
+2j+tn4pZoKgT8+ZQJT6rdOBxcCg8JeR+Y7Eh8DQTuDrmngAETloAbfLJLRdwZX2pB/mP7/1GcYc
l0SvD1ClGNs9PItZTCwwAWy05TBviKuw7nWVdXVmg8xBgsvnF28vwp/9BoiiHCoVxCNkzgmPzOfl
P8E4o9QKip+4LOoryMbUijWEpC5bWhy/YLyYQ+kqhh9u1UqvO9gkQE3bDFkpjLrxCYWW9d2NL2uC
ZWua2QiwHP1Ukr9eOtktcInEVdgAsYvsfXOmYFs+U/GPinerEB/4r2yJaueibJI06/dxxC75cuii
cbnZQvVUZw6bobgclD9PHxPTL4FhI/AQ2DDv4btzANctmPueMsO6kXrXJ6ZbLvcnxoOwEI/auZV0
o3uvHqxRHOJSV3iQyP49H+llZaIn6jm/ErnbYBbr1LQ9279taR9y2jNMLc2p1ILoOX3rA6td5PJy
81xk2uExWaBFyik7uxL5dKNN+CmWpFSAbGSmVEqBrG7uA4UQdnK1v2KBXcqxMiX4qZArqk1smhgN
4gyycDtgEi+kgXwTkRM6WjrW1Cb3Ym1ow2NF5tBSpmiUuEZoTq9kIOYadB5fkNpPp5tirvTSWMBb
OmUilKI8XH5ncGEpHX3QrYI0k9gwFPui5Oy6nCyYavvftc7yW5sAqWoQWdeyARO0pVbKu+EudnqJ
Dhv2SJ0lSxqdo/KeQwowhmx2Rzpiq00ksYln/tWuS6lciZVNGo74DRE/eDfGKmLZY0mANv5ZfuqY
21YOh/Ej75N6yQMwQ0kaD3nTDIJlIOPUbneZeEkjkjx4rDDZex5LnO8FElEpSTdFSBASKXlH95/Y
CTvZvf9MboP/bU+AkXDFehApEwqTHhBS6gnQrBcp8Du//hZ3ThzCfJTG9RLjstdLgWdjcBaB9/wH
j+tavN/ZmEuOT5DgAvjYqUgsQwlo9bTtrP3CzXZxtwHVky1CAwFF3PjcrjLVltaxYEN7QFjq28px
MLF7et1bj8NTwWnrFYBSi1PJCpZ0gWChJOhMMr5cBaJ388yxAJjwnKZgMkksa206xISyfjs7hCIZ
cFoa7tdAp8vShQuXo1c0Bq3Fuhu/Ec7TQ69JQylt2p505ILIboeb8PUa+s4ztwzM8ekbpn3LI5tb
eH+oanIhkIHiYqaMRGEF5LnEXUjxs/BlRbJ6R3sY90uIhFY418GX1c6wJKRtlz9nIEhi7xZkmIPS
6s5COK4triV5GNaOxQCByoLx4C9vXeEoW/LXVCeALfa8mEnEtHxt1h8PTPP7LOxTXy2XKu66e9fO
sTrqWMfJes9C7vcXFCQnLTjgWn0Dny804F7BEvpNNb3cbi/p6YUC0dh/24Anb2fbXCE5Bb7NwDq2
Q3MvmzKFXtpuvhg5A4hPeR3zRID6Yio/8dJ4+4dqKGA47dr5uhu6Az/ITIyKpuufP3AH386sBnV7
crt7M8J4lBudXZvZYqQKLafZKB50uYwyMwEV+duJ8mWPq+7mSQvtLzfwa9GT5/alM2FbdjtteWsE
ifIzbbLeZ2GDlEwygIdAmMHB6frWVpmOaeX4GcFu0r9Ok8Y/hLQHAmU8Dy+jiwUxgX3EtZljhUWQ
yg+tyCgAzOKoJ0r1EmW/CYPB66eaGSuopHHNPgoA4NhYqMfSzq5At3Q4NmjhVfSNJgYNwZYwb4eb
Lf7fSkAS3048Lh2qs3DXMxoIdD8h7XPVinKofP0R266H/mAEXBmDeLMbw/xEi7a7KRSd3RUBqmrQ
cvZSp+oF6Xp51yMGs4JCJAMHUtR7rS38o+uR9gIyK/ZfAWSSWUG/PgLMBzL1F8IYWMoBOgX5ZTLk
xjWIAnYxQbdcvNY9qnsuD/54CG1MCMmE6YTa0kRvG2nPezInAgg+vO2zJK8vjBxREvaWs2jvL8Kx
1I+wn3lI7P1FSELIVRrmBiyUCZ/OR1X6uiaYRzu0CPslSD7+Ip1gyLwcqri4CIHlL0AJLpvStedx
N54xVEJB4EAVzXVp7R3wYRLVVhj+eRr8qNHSMKSn1Sk14dtSdrzkKWUhfz6hQtP9FHlQSyYtKTHW
BJTU8IXqbzQ+7B3cUhuT1UCBWqDZ7K+WcJtMyOuFOZfnKNybzYX15g85FJRCta+IBZshWRq/y9KA
z04dQBEU5gDtpLi1ZD3XsYe3yXYCdW/6VRnA3zuLhxZLXHaLQbQNRHaRSUCVaOQEET1yTmfKe7/Y
2CAv+Y4Rl7zjCOu5NXEo1NC1i3TwSHzFKxtfoNk+13bdkVLWKc0qexFkRi05ke/4/Wj6Vt1qBb/0
DYWJMn97x8qV834fiN2yszS2t0NJ0c6uBCLn9W8W4eAGmwR/PEWV8rK0rJdHX6vdzSdFKMRsCFIb
Sz8HAhQ4AzGr5ZeXEwHzpXmZcBvOUTlDVcmQmd5maQk7a2X8xoeDuMIXVgmPTxUmuP4cssuSB/tG
tKD+0sd2htL/AwI4mB97wLYF5VCekwOPQ9Ux3ZMdVArT7eHOhpgvHb7IAY/EzTZQb1qxh7KvmB3p
u6dOWX1ekMdai8Ux85J8krVH7sz3pmIRokBMi7jM/y/Ukr44gf5Hs0ayPegxH98g2QwXO54e/NSk
nSW2StKUVN0kcffwC/AtcceJi1zjtK7RXtVX5gfdLu4ehoF9dVrVDU9qU2UfXUPC9dk44yDdfTL8
7XKAsdi/K7jfffelxbb5TDe8w+C4w2p5LkMtM+Ld/BvKPuCFCFBFQdU4PkPiYLOjDHpRpbkQxZP8
hsDx1Ha5VLM7A2KrlDTa6El38Ny7ZrmSUWtd45xDEAiAbl8DV88W58yq9bHXmPE3DTPvTs+8PcxR
H7O/5e00gmaqut1tGg8FDZ9+Qr8Eq1FzcwrFAliOm1hRTzm0xubOquvoGR6+/JLAh823Svpl9XtS
4ETkKYRa9oaX5tEAu8l7zeY0jhFP1qQl8aZ3Pup1pnPvNNCq6F+LYV0DviJMIsKpZR8iB3aQroZq
kisK4vqBj7TmvGQLlErqABFshWeSbJqESzNO77v6scdvbAW1dcDTqJhnaXJmisuMSChtg4ZI/NvY
lRvR0msg1Aw4d0Q7a+6+MlaQR+g9kvNwVESTpjaNRvN8O2XFb7UxJfkb0f4B/1nCq/zz1O3PrqDY
gorH+8wDPZXdP1u2GfTZmiiyRJ3JRj0V6MxBV52KvP13V6otBX5bNGQTx+O8fhe5dzuZVqr/XleZ
OdwRP7LRO2KhJck7Dg5tdE0gJCpxGfJQ9P33777duE/cDimb7UiPJsF4LnI/vt+7mTvtl7CpJOEr
y3YQkHE6NYxsii01oKUaF/zUeQbRzwMAdm0HT49+Tx6NgE9jy1+iA1hHqsKHQF8quAtB8d8CSNRY
AVbvn2VZjwV2lagU515QU47H3z15131yinqn/Gk++MR0hpWNpLTYtGP9x6IG3t9Rl2Be+e7EfTiN
h1gcZ7en8FGoALlv6Adum1oU0dU1FiCfC+XchPFYiPXNisQsEqTXuotsWcd/FbOrklvc/86WDtWc
qMgpLepfWwLbEQKN+QoRwm1vb6kh/4kdewGv3VyUgqxFk8NueLnl1e2F9uN2H6xWOHYMiqMo9bk3
1/KT0zs+S7bHk95NvQoNzbQemR9fbnyb3ZLH7vDf/lHWUHfRJtLsd81gmQbF7CLLRV+00fJ7Edom
rcWNTL/e9ZiWkCH3nQN7FevQK+sqFMem1XPWLjep4OM1Q6pym40qOkEU8IgpbhT1VGPrEDEETx2o
GVe6/+mwmHk9xlZz5cs1wWg5Cg5+55DQz2SuvcoDPe1K7eSo2cNXerfeQkmwTvdiqMR13OQQwUG6
GLQvW/auf6UiL5xJ87X0ARJuVe1n3As6hAW6AW9VRrnRu/XmfpiD2W+dzS5HAlvbbasDxCkmRgtJ
8fBCQe1ya65bJUsYct2cY7sSXDgcB3t53gFXWo48y095JsRouurFjsA2Ru3iGXyaJuQXlmVoo/u/
5zpn+vAN3X/KNcBUe7GvyJuXBUe/vP3nBodt5Zme2bLBS1dfHTTFvVcMzEsJJimx21iwpwz2QhtF
6IqOy0CFgtLkhboUHslQ8HmGIDd/fdwK0RZio+nPtf4w2pVLuIH8CUlvU3Zy/aXYOASZEvChZZtv
Vqu+dmtfqBWRY4RNIWIVSnviq3nXZ5qI3fp2AAKU9SxH6B56OT2lCeSXTkyUZQB+aJ9gP2Sdd1HT
cf1IY9e2hwO0RnLmJJkkz+QD7otY/d0H3bJ27ITtbiixXEA1Nh20JugjTyXeWxTJ2rY0z4oT8kvz
8CbqC7UTcs7KXD7o8kLEnhCdBtAaWY2BLQ7u8Iujv9/8p4Wk+TiuTVIIwJ9M0NfNPfl5lF68ps8M
qANwiQoaLDvkUnOuqJgpESWaKOzhzef5kgm9ABywkTBFTnLF+KdoeultVS18Ra6Lo63UqzlWWpuV
6CDutJhiISD/m+FL5MTwTNM7WNeFHvTFK5SGC2ggzHyFRgLn5P2slDB/nFM6vwbPNHG1NkH1HRbQ
n8ZjTCSvLN/HHaHfnaaaBpz0RjmpfPb6CjydYcqN5eNBJ6hZKcF5nTG+e4mbVgy3y5l/2MRlRBeC
wyNESzSBOtHr654rJZ4XPnBhu+A03XQQGZ/NJeSzzWVot7fCkOoPngBdkgGtaczZ95dAHX5JScWE
n4Y+noX47+ruAY15CjWGat0I4FVdK+sPgfGdkPjhIYv7TkxkyDKczO3zMaW8gw082vVvc9SO6NTf
iZNmnYPsLEmereJcFcSg3CAlUA9kliKYVYxeuVK6/iFCetZUsuv460yIzdmQugI5aemkC66X+R+r
dlnMTpJPq78FAB/cGQYlJfS75JqdqEOU/83wS6rndgWv/a7LY3pdvmdZDlBlmId3apm7MukxUJgx
iRJxabDyx56fYMAOue3XEkB4Ru1QFOck4ISlLtrZnBUUwfZPVZ9D6kl9vklvOAchg3WAEXlnCscf
rhL6yzxZRySBdOzrlJve5XC4CKWczogMa3uLTpy5gn6OlWE7ydpaKRqxEINgcD/zRa5IQhl5XvL9
rk7ZIX6flSQwX/EPPOMuMdHzSdznfBvsEwCZRFc009aQPhqc6xsf8+8w+vFsxcWC9HcJUo/eIwwv
AxKYqTrWZtXlTvpWzrYiKSWDcFqI2RmNcmyTCuDh4gZH8wZMbRdQrATkKprEY2+a66m27HtliYO6
fnS8RQHXmibgWYAHhbeCP8XsWZPMsCYS4JVHAas9g1inWmjbsqYlRaJs/+YJekXy4LRSuvVjZNBR
rEuK5sn0rFAdMPfcDGihvOsZy96YvtRSYLVjZ2fNHvqJPinyLBf1b2EVmntpAJFWAqrUVv6d+lBC
JFGOCVQzpY0ZsVYsR9Jdatc7hH7PZQ1JmsmjykwnglxQXk9XctyZhQqbP7FQurJ9uxlnZVaAPyvy
JBwqAXirQpzyZwCQPAslIJNmZaJNDpsjSrUx1vZZaRvMvXWZoeZsGKHwGt5ivaW3k7HJ44yoDSV1
tOycE0vt70W6ijU4xiuxkeTUh1hbZ+A+mXMDxlZ4sy27csg98nNoRfDPPNAAYjHt16X6K5v9rHC5
J1I+ZvNCIazjOvzcLk0urAm4qAKbpWYCpjQwImQi9Rov0lQ/3Md9yyi/T4P8GHJIWyieDy/aly1u
9FfflXCb6FUhdMgVv1Rn1hQpwA9DGiEzi3nbu6cmykWW9x+trjIHeMx3bN6pg5yTNwsZwER17jyO
gd4RAeS1uR7hWXhcPtOTN/81GTnVKVgzzoclg3zwKQP2E5KF1m1H57pzH09rQOUa1m/6q20KC/Dh
8ZVqYZVDEDJKeUIZ3FnjAPEhPBpeuu2jYPS5OHrHNVKydabj8AM849Tel/JjS8OyMEPUdkfFYu58
mPESsk8sJEYZitYEn+3AB7l9CEqkOpbkWTBuVhlc4BIuPylQvCkjuaiW2rnBkLS6OgJo3HhaHO0J
rGizTVM2+I1h7Znuyubqx1iQrGZRSq+uc+k6Mg1RZpX1QgKs9asfIthO1zuIlDFX2HA1GHpUB666
dQcbTfdOLV5gWKuUeSKN2VtuU0JOjmy6BroIq5hf1v9s60NmJxgG2b+fH6bC9I3IblOig7hHg0LN
QYeCDLqNDx0BCzx1OaeHoEmsVPG1i7s7GTEhEgh0jboN8LXBPUrEkY3J+onsssRsS8YIxRb6jPfz
Yv9mfys3KWbZPsbdO+3LczCZLeDjYvfQ2xLRsP6sbzTtghozCxBcKtlawU0dlO9Qp5b8ghIrleOB
LqrcsJQhUOIDUeebHRfkMVylZ8vLJ69Cq7Z2hcyK8BUU2Er8wMViDoVP6AIz7IhO7l0i5720stHr
2ceGfYsc8M3Qbg7EpezSuIez5Is7f8sV1C1hzlfG3Dl1I1pZjX7KcMzmIkTTGx9boKYeAWGo3Ghw
WRYE5b3CxNLZFUtcuf3JfZO/Am1y5L+M978WOGlhki7l8ljqmPEY5vStF5jHeJcfgl4fdqiYilJZ
QAvmkSYPPRYKSNyPlWzuu15KvGKkSgDx/ymFOPrBOj8P0yNcgaurDr3p31xcj9XdnMhedlFuqYy3
tzFQW+hpbJiWcWM95rk8zwZ1rfJVxn0+y+TBgoOss8UTIRWND/c5dq6WcxcagcudHUbSlGkvkiag
HqrKz689ycfmCuTwV3bix1qj3XeLlXxtlD1DKth9hAWedaAVHnsA1s35sWQGYxhPvVV+D1usuwro
6OVtz6BOZwssKj/WPWP84AcxWmqe/HMVcdZ6wx8rBexocOuxUOt2bNbD8+K5eQ3i0Q4uKOXZJG3v
6sIoBdsOVou6/ynpol3goETQaySIUF7mLM0WWcpoEHgWYj3CocAvbeXhkvgg1QijatTLDX35WCoX
W1gjWz3+AKJTYfx2hDQ7Ci1Mcumeqcr5bXFpA9p38bwQnqTPqh3yGnrnT18nKS670BeMN571y7qE
IWL/GPFJIRq4LgcmgFjGJ8gOXBDR24PhxaDvsiEUgd8PmQhXkBDp+RoP5PMnHLkD7wm48LE5TayC
HVlIBF2WBSrNUdocak4UjfxP+9rOUpbOEbSHSgk4t3HJvYq9ccIlmJXKIz4wxDJm+5f8SruFB3Ns
4i3mhTSa1Pft8w4/1Xkdjqz0NnqzHVBFCzXPAoytCUk/LEMt6nnOiovxrw06CXEqRrIjrBTrou93
sotWU3E+7eq+K/aYSNmyagj5jjm9Yuuv2KFkEw5Bgzb1m1Y3Eadh51jYzmX879UjY+MGi+1tXi6X
N1BjALe2lAmgYtkUjUed8zTXqSQZCNcbw89A17kLrDBjFnnXkCfs80RbEt15bNP6j6+AmX7PI0dx
xlRxUxVcC4v5F/A8EIEvY6fMwC3v6xjiIHZxC801l6HRPVLSWmL/Wwb8kxneHU7yzLMn4w7pTGwR
fN2/omkjbxKxd8XnDlYurA6aXXofQO5DAo6G5+ZoWeDIfff33kcj9IXj9sVhv1nQBElafRw8O2Ol
Ug4TIMg98zQUHtj+pi252CnTy5b/64mSQysunOhC8g3Urs2tCjZpgWwFe22mknoRg/JgGpznrWI2
3xutmyyCrb11RxxnjA/DiOPVM2mz1kVJdoxYdH4eacn2AXk454OpvdP7Txk1eLSSzXDZ6HgsYiRL
cA2p3eakX4czxqU+ldY2MnFj+BYfF6AQTKR1gcejhNgsPHebIdCknrtysXpJt9dvbNGTnFHRV9uz
cHHmIvBCTCGhyrbJZYVgVzMN2ia59owT0Qj+B56uFxl49OQLVQUdOxwWcBfn2sHInEgsfof32QI+
ILfCcu35XdUjcBUd4VDBnxYDgD03qyjlPQj5pnK5SjpkTFiOoD5w3+t7krj6k7LPRb5LXakLgLMx
JXDaJw3r0gSrRePxZthazD6dQse8v4j2r1wYM7Lxas8HlE2p1WdPEBcP1/SCj+TXvMefzvTf2Kha
kun2kIabXNxtyCCB4ODxwyPs0hKgWUbRwOZFcp/6Dhrect3caN7oxLgEZ4lXtik++jHOhAlRs2zD
08DpOnOcbdUVEu2BfeHhHQRF63pA6BfveY6o+y6XtR9v23ClH3015f/g65krcl9C2RQcvR+W+15K
FyZgUow6ciG7fei4cNNrEz220IjZsob3FAsNfERyZFw25b2pbfnT9k9+I+SGt2tBqMqzr7tkhj60
/dFNHn/6mXT6aUP9TvwnqX2jbukrUBHHtRY/V8u/FfZJAfKoPBe0w3ifVnWWug8WYVX27spwittu
DXaG4/uLhYvyFMiE5DsBFcRmm1E5YcoispV0DIoUdnIQqGz4l20ZcNfpvr1a7MKH61i7Eqhrs7gh
EqbAE7LPXeqols3btnMHVU7r5oTXhFIFeVLxEr9BdWDgAePMClEiSRY1N2mYU2L162eqVFzanNWv
xcZQr56xX15HVTOtCmFl3bqJ+zr6D14Gi2wvTAnpbPsnR0Dbbf54TYSTHa8Yn89euuxN//SKViGP
Z9KQit5u5SZEfNKlreAUykNbFi1/XhluJVsOhZfCeF+LMEtQSSDt5MhjhpIf0MzNXJfMsGc0RU2G
pcK7UruRKNAZyglur+t87iygJ0KYEzb8gu4XqY5zYyx8EtPvP/7D6iZqmwNo1nbI26czOhO2Vlg3
c88CJnrjY1DY//txzuqQ1fxwMAB/TOspckrcdE3atBlgtegMw6I4LvkKL+W/GN4imLK76M4uFiv5
QHCRaw3j8ij0WEHDnh9GY2rM0kh2tpTVysYpa7kL21VbqSTz0EhjHUfoaR6bnY7rsm+LU0lz59VR
YQcvrAF6NCDfXWBPPe0/Z2oiAD9Loomah72ZJQvltJ9h8dsKU+Z1FB7qralO18ZkY1nOMObB8B9/
WjVSqXO3o6pg8KWOe929AeNaq9iFpBRRphVLSwff3bvJHjssaRHbIikDNhgByufKFxePVnq+czbR
pBkjzA89jLwL1uspHwzWANcTywmyg01H220wo9+CHRL0aILzbdPm6oOWnFhvY73fiQ2eMynMcsOL
G3by/YVV49jxufmcVIzs5UhKDs4v66KbfnsK2+SdLGkr29aBemnZKuwDRSNkxVJ+JirDHAOGdHbG
UHxOxN9surzM8go44VffUN69z+P4YPEaL7qUtUQVXrWa4cjfOz+NFgW3pvGM2ydE4wEM1gOa2m8t
PP1ni3jlmL4weWfhWUtunWWBGv58AlrhQTJ7nAY2MHL28RgVpPkMyN7TasbJTArSZRa9xMWLrKa0
FG+ik7rH7h/uL/PgHxS4gkeKa+RXPZSI5wpx/Gby2iBJzSLzO+xKpC4COVpfdGkfeel6ZFbiV6qZ
31B6mkqsLlIbebrRkzb8+fD/lg4x16gVcqcYGa07B5Ds7WZGd5iuavf2xOZZ/wm1/N0FUn6i7LW7
DzricgE9N26MEhlbqBgx7R3nELhWjVFaQywHxK7iaDjbH+3FKoy942cawigaM/iv8cDTMWqUjgKG
A9NJqG0J7xJg1Y6txnEVIyEQaeLucItVzRhj2ksH+IT3A8PozPLTiZ4c3UvjnJCqEyuSdvXL5krv
ZDYWdX+/S9kxfOcb1rUNfVCFz87WYxO2ceqA2rgBkp9qt7I4rtWUpROXB31Pfw43wLgLWLzo3TKJ
+bCYTgoDPcKwUCqu6jUqlgOef9FADQGA5E8CxSKNQgEwpq0y0/Qp2zb9ZR4+e7i/RCEkIb28WZeH
frvjaBiZvPESWjslWGP1Jlxewh3S55MLehHyQmvajhFyIEG8F9AlgUGKe2bRkZvhjWL12oOAKnQt
cC4yJLWF4LsObuSpKiYUIK0y4UZqRprbzS66L/xsuOqWNgqMnhsGK50XmM49xa1u75KmXxtzsCNB
JChWp3/jiSjEfcFIxKESCFedLQKCvJBIC/19Eo2Rynzr4QToVueVAxAnOElctkFABm8Onkav8K9j
YtsbfdwpExZEqZ7QlRLEjljBVoazte9fB+YThAADUJcrSym3k6kv9NKlA+DiijYdBZZcq/dEowV/
+5ni2KgjIs3axNAh7yoMv5iBEK8HQVHJ2APtT5B3GlALcl1g8lNU6hbMsD0hV88koknY2HVTai4J
9iZMHMu5btCPC0yNk8xCkwCddKi/98HrqGwdiQeJfK0NY27AKD7HdyyKFXT7JtSboRuQflTfmbYd
fqy3DAwDXze6Sc1ArWSPt0dG9qwrhmDeT8+PA8wPP2H5tZsEnZpDKgo33NRcpZcPJA3ufGPO7J3n
HPh3vEaZGGpJH7ZUSVgvJ3lFJqnWxuvaIrZZdvtoHd5ZqXz4TwoIHujs8j5AY5nP+F+KvctpE2Sc
xH5NZW/Aw3XAtsPJwAi7iezBsUL+qdodKcJYNC7rFwwEdqSb5aOW98p3qv19/lyfHtmIsRyha4+U
6flgjA1FgHcbWOlZpAbhtxrzj3YC2oZ/TsaCJ4o2/srWFqN8o/pEhS8eJB5yxkmswVlreGUT7/lT
GmPGypC8Rq0ecF7mgzntCUhrIgPUlULKAPNI2bed4S7uCPzBIgyIBkouae3mnCUEDoBCBupOQhWV
UOnGuT97Nl5tpnTavVpY1QPeHD2OCyZpda2zVXJ1KqDzdJDqFCTBueqUhatWvaRAD4HX7ysWfQvb
0TFswLZ5tNi27MJWmAHrK/3ZieSGaehftZYWMaA7Rz+oUg+08DkoiHP90bSACZzqn47DGzWBiV+P
5Dt7XpjnQT7uZGn7iTIFqHUHUtN1tu1BHE0g0Pw3fuB61cm/ZQ40f1N6x0fYZbCkT34xQwnylJ0c
+jr/Y7tummpaHSmZsPvv6pJ/fKPQfH3mEkBbQhvzmLlquKZsGhuSKsXZbC3/sBaLAvrcsKxBENGW
CkRv7aSEvI5p6nUaJDJoouQpWyPoczz1vXHznWe3ev/HRSve7kFaElmz/vobRzAWfpeY/ust1hzH
5BSzDTuNzwz5Pa82fYnpaOKDZsdxKuxIeNBVRTyLPhfuA78QQ5kenUujatTS9CorNGbGGSMefAHy
O6RHfceg/YSuCrw2gzjrIVfcmFq4UgNZah9Egxbu8ZDl2EdmlUgOveCjCl64InZUbdNYl8cmT8Pn
pkdGLm5UNlgYnoF7IMI7ZHWDh2y16WDF5ikdqwCM+jvY7dQoZPReMoMtybSwd3qK6VH6EADhWPdR
ylq0ZKwy29bVHlwtD1kPH58D3FGz4kep9oEDCNcUTN661UO/VVQJdUpxdNQRW88BSMbxU7l1SqQK
KNrA8kEpCH+xTRJao/Refe60nHyfrjR7sDmUnm+jLFTqTFtaK5gX/MwQitmykZViib8bLaASwtqQ
2/GAgkE/AIXVpfwdbfKwyNYcWDmejOktDi4B3QuQaiPxSffK4o5uuYF2U5omGtEpLYXJcu34cyEA
tv3pa7+hGuPcagx6ZRZVNhZOCm3q/ZKikMljD+KT9uTBPNCYRbM5EUnqv/v+hqZDzwpvMAR8VJs9
B6YobdpTC6WtH6XGQvKbNlyBblV47Ud4+sfIjQkvv35CvkrfepGlrzlC/WoLEl01WIr8IWBEdJ+2
9uK1PCfiRlvbYpsA0495YEDxT1X3r2oyFdzRGSdW//35nQ2ZmP+vYgkhBPSYg4tO48qp+ZhZEM73
uHTmBPSejw8fQslNkORm24JGY3PLv7AGyHrVBYSl5TyMPZci72KmEkr8i5czt7bkv0btcv1qaZaQ
IVd66tJZFWl937U2Rtv7c+VYCJD2gab4lhry7kBEYSwcy8Klb7fLarnsdp2FkD0nYOMyeRVHZpev
+p2zm9N8onETMrPmn5/wXAxPRpueYsSkAyfSbl+YAo7xZn8hCkpKYB6YsSpPb5IvptWfF2PN6N48
MXhumZ4W8Zo4Nfv8OnK5gaz4yNO7tyTeld3gz3mfIHKEX1mnNS0XLwg+hUkB0kKQJKczf9Lp+JKa
SU3Rn18c9tmjQalzZ6jZze9FycguKD7VtvrLtr9I6+H53NoDJYYKSBshu0Xdh/BWmouJeac9yBW5
Q9mwUQu6HNR/YbulcawsQed/Woz8ULOedS8mE64mdGSTEm7++HAuawoom9UgsZ+eTHxTXE7Sg+Zq
wj74WyWZSY99w9AThxjXe6N1qtmVkWpTnJBKQCX8SuTiBmzx/DJUv9/Un7P4QOD439yPwV072GSi
/MudAzr3fm556Gz9HJAhfYvpa5HvZGUgmgsBO5XlYSSqC3BASsHQcvFhI3935IkZK9qFaW1edzFF
oH1WqnS+Y/jKRSvkH2FO3U9Xw19y4+OZGdQHdTzOqjgX/EznbBL7tYq4oqk/wH6gH+715WkMisRF
QE1PXXLNUesqLHH88s8P8pvv+lzZkrEnDwAAl85TkSjO1y7WjqZYezaTPFu4nBobXmA4PPlv4MmX
dqwPA2WzOTobXtwJ+laikUgQVpF5kkM9U/H0CrVcBdTErxB6jbk6ESx2z9ULWAzkX8kukANBJycC
bDBqYKxWHCfl4VYeJICKZebFXc7S4jyuBFE9MEhozsbMcfWwNT1/nUF8d5UpSyupTlCQmRm8y2Hh
F2y/hz8Qr7uMcZpXqAkt8CfpeiMA0/qpH3hBU7qwQq/l11286Jr2JkPFrYtZpQmsbDQ10IpNd8fj
IkGkpixW5nEKoWvJS0Tat3sEWOqK3WA4uwT61KKL915mXptA77tol7ZJ/pfrbS4JoeFawOsGt+C2
djZtQ2wN0SI+rz4kL2oXn5IHbAopDBVaOknsWRbMJQkUSzK7Nx6mHbiktitgYdfC247fcfFqlwYu
CdEkvN6fSRbCxcCN6PEv0ucmHYWdOO79t1V1R+1XJKyHHnijkvPeWh3ZXUwBF+vJYjvXuWjDfq7Z
Ivr76dmU5OZYfu1pWyKF3NwZau1fT7Xd4Kn/kIS1Ty8loZjAeCDV5nGLK+tEmdrtav6noVFa1SHK
2iqQA6Ctj7x/zadrc02K/RkmOxunb0SC9pzKibC6JA5zjORXJ7VOygXrxtXZXNpQpV9VauWgfb2S
sSC6Vv4QPLtKNcSUUjkJAlSqDtO+Neno01PdF+tNllT5Bpan7DK4aqRRohq2nXzEL9C7IZbp5gXX
5RDcRhFsMJ8ELrNZsjqhFB4GkiqYlUoVJBthH7ZG/lox4WynIYwhDMw3bLhOnklZK43RIZUgGZif
mdVcamMbJ0pL81mWLk3n3dbZZsyQ0E05MknCYvv/2NbccYjdWM/m3kT9jiJyykDR6LYXqIyTRLrD
P8Tb6blu0xZFP5ldkE22blAPtF02EnAd0bP0kpiOi3uvYUt7WFzGF1MybdiG3YgFjepuP060KrYF
VngrKSuBd4yhK0GCc01Fk2wqprKjaqQF83CwxnZzRmAlfzfSafLLULuwKKCBEhZ/f9TK1F1nk+aX
yPEEWrH8Rkzsu8h+wWXVFSNP/zFRcSEoGGfP5ezVTNTOQC2s0yLVSquS7manATZtjDznNgCSHGaM
pEX9SasyiwQOBGS1R3du8CPEEjrvOIKE1F2iaucCL+8/M1CCqHRfiHNqQO/oNknkPeyVSJiFtSlo
1s+HkNzxlbQZMHuaGNPq1Lpgw5xYvMG9OVGQvJn69+vwRk58pseGKxe8+BCnGN2YvtPXl1HLtdEY
C7/rTq7l83lRaBdb8ZQcVfd5at0bMySoNOW60EgQbgZnK6amSJxx2+D+NUNbqWJc9gz+cKoYBqvR
iPa8Q2Ir36bUCp7FBaAskwghl6be77xn5axG1uW+Fvc0YcLOrouBQkJrfTZyf6U4U5Br0Ye6EztI
vo7JJ1xz/EQN17SEwbMQWom0y5Mk1lowsflhJ1o68SB0h1db4zpPoYl39pLo0aczNwwrxDg/dO/H
/obglGDGUi7Y0eyhOT58yfUOyi/uv3agqAqRfENYUnIrUU/b5M6092RySklmWSkqcEYlJg4yP9ck
3tvbpkAxIvROqWDdtviB2O5xPZ/YEQGnvCwMz4+BTK+uIYO50C2XG3dKCEdxZgHxPgYH/K7sRwBV
4oNgPbSSMK+x2P5WdDA+NC1f3bJSW01zQTM/B0MkorZM5PhRbSRWJlYsEaOWEIA0PlUwmMGb22oU
zZVtx2wWOhe5mGxph2ROlNhNnAqTKJYX3xeeu3jJajQOe3Wkt16/R05T+y2+ZqpgIQ22bi0EAH3J
7WNSCR18p/Sd0snXjLGbSo2fCNlf3meKVhKBUuCFrbAZYmviBbdpRx+roqy9nK7YDB97LZIB8SQ9
Echf0Wnzdp+jKn8s2smU94Xs8UhJr41y5NKXmZ3OzSUIg6yapxvZbTVLwpGkMbJBjl4ZC7FK0EWM
7wmQ/gz9fNBH+H3sg3HdrPh4g+wZa4qYaXI1UHhJo/KRsF6FXAV8IWEjeprECDH3DFmlUPrwhnOT
ZUYelOu2wk1KvV1n1tlH74JpTjkUfbW8xyjoGpCvNXWMSedn0OaNoAhlrIcld24R/yF9mv0w85A8
ooma/QSSi0Chv0OPtPy3cCqVbxzoMNi1OyvIITPHCzK4AYYHz9Fjh5OswG1MlhRdpE6nE/tsaUWB
4MbZiPyxjhpeygDkUnREjdAE2LVZF83Xvi0xhYUMeb00/CyVnBxvmYOiA7Nd85YdrjvpTZ/E+2m3
lofGHkTTXKXoAJVQmhF9PJYq/R7VeW3OI2Q6+t4wqWQyhbeNzwsDKjBE6WD2lJsQ7C7thQXsV6RB
IyL+n/OiQaYK0xB5Sgjq6wHQMxAcnNdoz4faySlwKL/1pQ9tP08bTSODXKRIwXysp7Zx0SMECXti
CDWNiP7ZBu2S1IBQzatnikw1Z4/bkv4UBT2s9oydBz6QnpTKbG58AcmJ9oPhlORiOYMILiTKD7iP
RCNFintuyKFI5QJco9gN7QSIiyfjyB5fxJLHvq8LQVKiL1svp6uRoqz+YOlYtfC4sIvEHN0ZYURy
HWE9x0yl3yBv8w46UQmbNfxThvmclf4rJczgCnjrrNJvKScv/eVVmFBoS0ma/LxjukMAbRgLHU7O
fjGB0SVTCDb9RaalAmk5JthXR6eMaLiQ/5zKAWCM+9wrIjwF2+JCzItWmBaerl1D49q7Nl6Nw7uZ
mjX0uNJVyceJJ8gmlQE1xDNx35Uwo1T0do/QhKt9A65JJ3X5Fi3pxawE+LVrwGoqlipGaEaf/92J
Qe5Mgyx9tv9/at8enpBLgSZDRwrusev+wl+TSWqw/zk4pRbd+dS5mHvbOLxdk3ji2T8O7uTH2k+1
fY7swZDg8ucFURSzRUv8cItXB+o/JFOdf+zxzUNAgeIUdgMNv/k8Px1MvCOnRClOy3yb0F9c14jl
XlvGwVuN1giSt0Pnafk9gPG4LgOS0ldkKnMjdTOfOXGbbItdep6aEHpdhe2BGo8huwrSHbCN3+RP
yE6PegAh6hHy38Dv4csS6b/g9IK3MeV8n54ejYnWyby9wymRD0p3Y5QZNKHQnVrRma89tUXuo0D5
BVluc2ud4VL6o1UK+cqUqPFXXSEzQkByncD5rwXMJb4vPXoi5xcv3sXsJRjDdNU9wf+kD/0BhRbW
wI6qMjs4AYeYtLIdRqqpCOIqZ1jHrsM1wUSc3J2eWaNudduzpJVIcQeRf4vlp9YBh773mtHOcRYf
WM9l9uCdqnT9fCZUuShd7V1hl3ivg/BYfo+mIWXc53EzDlQ4xs9d0KxLeW2+jSE0zCsna97BcBUm
H33KUWckr8vAdcICLQq4RvEnevJve229xGuQcHoj277DXXXnVb8lv1UpysT4Y1pASr+/EjHi6hwP
ItZ4uQDXT+jI3Xi/L6hYUyuG96OllLDiw6xiXN/XGXFUAhuna3ZVlAIDmm9XOofUw6jB5Y0q8zFa
34UpNZcOuDC7jy+9bCpbn5/Iizb4kUGdUaKZe7vsK5ccFNHcIFlVyp7RI2OWsXboNE4JAKBNJvFn
c17dQj0SYSaW5dXC5RbSpAo1ONWToHoDzTtE/TnLn+DnmnnmS8n4LwSl2cUG8+ZnWVlEUIKb0h7N
jEOSrwjTrGdepSR1SDKTRY5Z1c8ApROT/fO5QTT/G83VIoVVAAGJhq3P1tzwGf0E3OwsbwSJr4tZ
wauW+0PlfCmXMnpGP65LQSrFxePtJXkTdDHVZqVtVc3wJkbWN38nFrYPBJ82ox+FrIwSh5MHUvXy
IF342lSsD+pwi2baaj9nJupsVfValU1BZclmchkGh38bHdOGdPAZwVY1z0Lrm8mOergOtQVmVad9
kk7lFUw+Cfk0y32fxz2nmSuFOIlj1+9qNDWRFZkoABTSNHpJ2f3xTs2NS621Zyr6WAYDjHjtTIVP
38vbsEY6D9R6Y334zFgAux4N96gffzfo4R9PVzuHR+6FaX2kX+xgL5GqyFrupqNoaxRlm5ud4rrR
Bg+6mJ7Go1EW89iBkrA1lIuf8P6Q5INbtaUFQyBXZIl/j81BQXLqE4Xz9NH71p0SbSYUu3eom/nE
7LhkWL35IoAxBtGAV/VMbFh7xqpql+TXHF1QweRcASr6WshQainS4QHqeG0gjE9a387Du7HR7jyW
4ERmJ1PFiT7ZPdHJVRwyafPyTS3KNXdgYpLVu3f0dIRkL82JmW8RWNTyVdQRcb25KymMzmOpNRLY
1nqGNYBpntX1cs4S/eo/+BqZKbAuslQ3QFBpobkh8/gOeEX94DUs5sIpux/noYEGzXoesj5Ekbc5
2WOZhZz4NpcCiaE3B8WJ95NJ9fF9+QdqQ0dWUY32P/VLwiQOMjRu4s2LP2GFFc6D+OQ1rs1bgbCb
XeWL6eOAbkDGYjBRHdh7N1IgISFL/DyjhW1xeAaOTrnM1dffmFEsrCIolZMWWry5v+btAbTK+7l8
Ri55dC4DSPIH/x4ADOtAtfE1Bbm3mPXKXRdrbt578j6FtGzaqBkXxLxqLAcjI37BFNtOe9lTWGph
BwsXxJBhqNK7WSQ02Lk3wtnRXd3b+yINNMI8DrTIu968livzIgianJN0GDzSmuJWIreXfgGngww2
ZDm8IPL1TovhfmF4hFApBXK2/d60IQlISVlaS1V07FjkYZqku2+5V0MiQbdnD1VxrM5BWlbFHrIx
R4jl/i1foAwsyW8LEht0zJofXEfxFSpwizYb54p1IQS1eIHqv3mjQyXFGyhVwASwVucJoNS3vfO5
mLKy1M7J87MPpVS0u3qNiGxiv7yfgMeJyMHnh5WyNvP68kjG5q9OxgnMX9+z7xEIXP6ugMMGQo29
X85DUst9JfHDKQcwVTwNJgMGHZYoE+yU1YyXhAuP4XJ/T3gGOsSLGgh/1Bm77RQbfax83hrsMm6y
iWUv6PqCRyOqyG21tis7bwKGOb1hA+MkP3qL/iGsYmO4EOHzeqEnjN+NKAUGIbvUL3CfrtqKXL+2
iGLJl/EFkhWn/abLpNXoMzkv35Qaa89dgLzkPdH4E4z6cE3YZ+7YfJwK1CUE1AqRuoovPViqAKwC
u12Rm/pZbo0JLppiY/2jmVrV6PfQTZ1+XSQ1BghEhARP0oDtfZzNDnFlOSBbwUPgsXjZkJRn5urR
F1RoMjsVq30xk+Z5ZOqEH/yDd1NaUOouMPjO6mRyQearLa4mZYh0VZPSWFUTYAsjSAabf8xOwUbe
y3zuhCYqapSJgaBLOp2t7boUlcMPDm3ciqove85vuUJOogNmzbf6vbFiHwrjUlUtQjN1XD399fux
9Z/0jPmmxbYqNxGD4V4+Vsz4Oux66kZ3VGrR1hCFzydez+pi7NaS+IY5zB/IPJ6kyzkLhz3BVp4X
4kqSTuvamlI10iVSGztaCER3OkBTa4gnlSpZjtM7z64Ucv4T5v6icgwELkADfq+XjhDfmvEuKibj
lFYToY/4dx/UmRPFfsWayChXCQL/kf2Xr28nkluSK5HaBPhTTc5OtKMZPvtD1HVReXbUnjyUuG81
DCVIWGQPco4cFtUlyQne4z7uyYc2qwNuCrV+hG/8MhWchntKW0Swj7qDsj33Q3cdMicMfzxOOA1x
JdUxZU4lBRTF2K4t+9p56QG4WjZD0b2MvtpeRQC9FYWVteLE3Sa4miMFGVqsgR5XyGdkqQAdYHel
6G4LGEi/EOfq08nBesKr0vYHFD32snMOuI09lD82R0Sd4lIvPYtHZRVgnjetmtFKAKDe4iSyf/OK
BDxMj1wlddoKsaFhRzB5znp55hfyJ2a5DYcjno1MJ/PUSKkpsc5C5If8Cptzh6wylEavHbp5zps5
OqiEMAP//t0/uZwWer1GqP9Vw1fA8bKghQTLf6uyQwKhPuokfzD9gAyvJaficrCP0DktE+NdW3PH
5gs38Wl9T6enXjp3G4O+i3+fafE9AIckpU9ex9/GVub/KDKaaee9NFdN6I+agQqQ9tsr3umFPo8e
iljr4X8PtlslL3FWeE/B8lZh8G+K9FKNzvy16w0Y6co8IK6efFOglMlgb5ue2rT9dzTBTthDO0/L
7Mi7lgk9mOLw9X5AJi0IXO8XcDDF22P96QN1AIo6EsBrNNpwxQYEvcuCB8shD2vlZiP6mF7a+iW+
5PkdRLDUaOdlkk0iztmqSHBYbmCDTtEI6uxcZnk6fvM6C4fSBS14cXnPisztFQ0jaIs0SMP5KfUV
mZ1O+JyzoA6Dg2oBvNFXaC36E+tjxwRLqGtvflQk0H4bIjYQgdwpUInEzejlhKz4juARt+GAjiO4
ZUmkjnDSkOsaPMkhyENKPssTfkphKBk7YMqxJ4oThivU5tloFzmezUAsO/6QujHrgbm8bnMc6Y3J
IYjWRko4SKGi9OChEapDfOWKtJU421hsyS2/pAVbGtjS1/EkdDZUGlHKPdhS4d5o5uxZiwWxd0Ai
UUE/bVf3ebWoFGrDx9lhtCW0kDl5asBgcvemdpse6Koi8MjrMHK5RNCBIlbq4eSosLbaiaQ46STo
htbFZMkGFzDK9qdCae684wZxS7c8WiENNO/z1R8FSqG3VU/w27PXLrz5zji1WCPmQO/pIZmgE/p6
oODuyg+eyuiztfREgT3kNmWSivcZQEGy/k832TdCAC6zrR7coO2L3ybHn0+pNDBA8z/CSjWqKQQv
+Twi4cZNkbZGONc0hoNwf3t/GDKmkRwXwaLPnfRCGKHdHeFved6fV02YvF3bVpsKJWUyOm0Xw01a
T+YYk6LEIu3eZvga1fU2QiG1e2qUmNcJ3GLJIoHbMSbzBRj4Zu+8Ukl+0AqceGwWFWmbVXmGRTo+
cWhpei9GvsJkdO96QWwQaqNsrl2BGo+aXWhScSpygw7vZOxPTEqeUZB4g1f89RvzyCqzZtd5FCTE
Nw8yDS30mvykYosIddPYzbNTdIuAgYz2OXzUBb7H9TD9ZNQJfDPKWYFExs6rlnN8B4Gjv4SNjIgA
wl1dFYcjH6sBKhukame5KTT8X61zMOAtVGawWjV5tt7F6qknCkwXfY3kQ76YnG+VBnl6fvzpXIRq
dqNbmRe+ZlycYre9z6qz7cfUDTVZS1Vv/3J/vRYJV1KgRJ9pmoI0cAitQGopKJJMqFsu99lLozQS
rNyP6xEYn3t4FCBMBDoZ2NOIUZPNJlZpwbBgS0RrrAOR4xjk6I34NedlFBio04AUwoFpPHZk0+gC
LTPNZTxr57qyUg8Ta2qqkKA9hBYTgl+cE9k5074oWGn+Ofe03wp32nizy+2obRC/MwebUqhFWxHN
yMf+/YZePd6AX3vR0Dccnwzlrc6emIKG+utSIj+icNoPLxK3ksXi9khkAbc3nmFmSYz60vgxyg+V
QWyVrWq9tx1ruJdbAgiCb9v0f7bcttVJd5jTPuPpHJ8BkicytmFLJqPQDMUWOP7/gRtMvnUUpdN7
CpR5bbR8hQXGSET0WX6nikMC+M6daUaTvrgGxCVXNavSJArW5i2QR7myIhAouv3uzXc41OMc0+fR
TA8A5/sRuYFm7YZKVlnv15sjUgLCJDZrTzGX2zJsxQXNF4zAD4YQwPBLkY3Gwpu5HN3Rr4k6QSyu
1i3dPQ8/MSZknYtYC6NEyGzrc3xh4yOU92a0nZVEDVp4tiFpRRnlUEnPMn+uAVWeZWI5CxatRdEf
jft9XY3WxlJw9iHSnWwjU21zxotS+eWcKLJlwZrTib9vputb5/VJu7cR4a6uUIgwUVP+6Im0brb5
ZbD2IuBY6TihsBKQCoX71UX3lfBvN8OMtC6PHDMfnVjeL5Jh5uErzxSF883K2fPRbxgvO/BL0MBK
Mmty7U4BuHbIWSBeYfNInKZghSP6I3Z92NTfLeooCTNMrgcce+2YEhSoGFCW1ZoZo+VKWWuwu1DO
uiHEL/RNQJBAwaFl/Bcsak7aro9ku9AAV+pMZc/iIjtLWCXKNpRfmE+KG9vj1eo6dBVWNbUxmc0k
GLxhoN6O5e7BDNIeQir3yuqGa0YHK4s0m08QUmzd9n26NHmnEu2y/n91bF8Rd2kyFa40SgAU5CBm
S96ZmYMuGRVYX0+14sfCeynw71AtBa0D0yneQ8S0D4X00Mob2b/OzA/8XHsrCHEbZRoLTd757eTh
xxKFQVrlMpeGcLKi/LHAQDJaWHA4UC/s5A68yfoEdJw4v2LUogH0bTSg7S97G9u3nMRLPmt8Gmv3
s3LQ3rTYhdAG7GhaupTu9X53nPEU32Idiwsp3RB3ZqqiUHtqqvqhj50uODmvxJNHzTg+18547N7I
0WU2DgkohuMOhr/oYc2kqTwyFaI+NGip5bDtCcS2+/hbKyCACclYGBWzpO7GjbSNmpvWQDBzckR2
THkyt4I75qw/GaZgWRZ6t03DT+hZ/JRUCbbYksuSCxGkvO95K9VrmDi6DZX6wEpV0eUnZBMCvzrZ
tmzha3HUnX5xcmovBVxxeTBNR8XAh3tEzG/ZFe9cbWksf9ZmY6nY7wMdrCV1YfDZ7n9YPCEmDsLp
FUVK1OdDRxpJTyHHSbjWVLcAMn/pW/nsSW1Q2tRXYBRTeQgGUgMVr9TN8oWnU5lfYO9kq+8IxNkA
d53A9gZBWNLcJgEB0QQdA64XtcS2I2rJ1eOpPCer3sVpTyqfMSGQCNNnbKfqlJdFIHbVGWlltFpx
kFuaOP158jRYXDrHnV+u9/XAgRAc98KoE98wgS2k8I5r48At3VHW0QudRRwA5525e1q+FoZ25AIj
Sgq9UsA/soyLimuR6xRscbBD6+u3/h0Fgx5eIIrsCyk/890gEJhg3tD7p7zOeoSRSCC/wulVwjjy
eVAC3P9NnkJGXjH74HwYdF2QJylNa91IReXHAvi2/OFj3ReUi/W3FpKhqVbsSDJjf2W1Twaj3dCC
lY0JrJ+HvulGwnC+lN0Jw4X9E7FgN3AZoWb7h/VUDpPEgqvNZl7DLD+fGixcrXVAil4AiDzPcw0x
M0cHxwQzo+IoQvUVLCQie3HIkmJQWHvudllrszGz6fvZt3hMCRyrQoRqG5KAYtcuM94r5wJhY26P
zYnK+XMSsOhCriOr4nPIhC5IxN2Z9CBZEwgUIgkO1/YbkzJSU8auxdq961+Z4tz0lyv/9fk5gdm8
ntq06AC5pE/nPv88KWzgfJcNl+hOMJqi+bYb8saYg+3es9GkcZnNfTjEG5xmdkTBXln7GCv9a2kY
OWAYCPRmGlkEE/S1wx1IOpHaYsT/8VKixuW0xIyPTcW93ANOdbp7VykQNfRXnH44oemEIRmiE90n
zWj6jxcQhNcNXAZ5W1jH9ZGNfzCM+zUW5FF+ko/CNXtAE7LO9rO4D31URiUn/8KfA2ZpwY11Z+gF
SnTIfRRcMs1m7UqeBE4V4mYDKDeRRsYnx4yBinfek6bW94XO+c8MGJqX8kDwoFzU3dKnSzjLkl8u
jNPSuatC9zCUn0N3PG1aHVeN49rKzmp++TixVmNqg0HKfV7fHAu0062qt/qq7dro6ZFSzToARXS7
IN+h78NOM/zj2BxPGc1Nw1cK5FxdQrHSf1IdPTwouH4eqRS+aAvAe+B6ZdRYyc/yMxb1PrYMFfHd
SpToIzOaKC9CKyZix0l6rnyTpOTSeSSj0SY5dNo4t55gLZIIrQIKhAaCpptw2jUsMqOjIyJkeqfl
lfn7bPg87XD6OWth2qtrIzo3U1wifIKQUwRwa5dj3bZgtsElOetEqmO83JewqcCxKXDDecyjK4xR
6P6KpY9f6OpbcVIojZEaD4aZdQkIxrnbW+2TNRQAhsKFV7B9AZRu8TJcpkAq8NDSyQqxVYKeXopH
LF10Z8C8hQwyc01CKhwhX8h1AUZweUde2g2oqS8BnfgvpfIyfu0X9Tgi7l6Bzo/PHoZcPTwkgkVE
hxgCU7FeomJw8ZnhBuCxHEJcIz3CNPQsDaNzdKD56NhOej1nq6EzmNbjKLA6YcswMFOl+DU28F1u
fi2JGqf/irEv5LQmNChD6AZp4ycQDO8a+5w9rQGzqrcr8TzOyKSQdjPnqcw0BO5sVEVM5HAbKwx1
96RZEHJf8Rys5OBJ8J2yIC4hZPFjuY8XdhITTc2NeYjbJwXns852BMqfH5/TeG1xJ0BxLQFppcQK
9IJK3kozN5o6G/7KkExPXiK11/LVbsJAlc5Tme7QNOxW4yI/7eZ3aZZc33MTRC/JryoDqG9rQey3
W00fEPacqBQy1e8FWpbDRGX/qCKB0PzLY31JUb4lqyxcZ3cpKF8JAoYS5vU/7EBXLR2Xjg/8U65R
8pNifXQAixykt9/XCt02dDaze72zvRyRZ2IPEMgukA3pyW3s6hvC+4h6DxbZanvHmVHVc7HWPMAL
lv2m1d6r81apybBS/1Ost2/EU4RQeEnJaJTpU4j+5R1SnAXUQKah7y+qPU0WNr2Od1Q6YI2vm+6W
AAe0CEKo3sHIxIztZ8ofbtyjcnlMdgE1M5y+S1YAxAbrSCIDzxpZ07fiKVIP97vRet27LJh1Vc8Q
sdcLvU/4BwKzMgU97NArPTeM25RF7Ae7flCZiKQ9KsNERGLdZIUvtVKxJ9ZYS2xBiRptCFDIVS8y
6VtWcrqIePwV38lKSGPIPDuOq622lzZ3CXhiTLPZheFEIz5kNFe03eQHSiWVNREn8hSP9If8sSFs
e/IbPtpWON3q4lQKvTUwNjbJMGiyGSDkMU07evHNd/DdW99icfqhonTRunl8sVJ7tPyVR73OHsOj
9rDaIkF10jC5scnnuJ0nsTkurNhyAkrsJo85Tw1TFSvl3Yq5tXR8t10vtACBfIxJzquc8AYPyAwH
aZ0HMtz4j9rd9QV5JyQ4irvuMIShk9zdq5QXm40OKXUyk07ESoLVHHgBUd+AwEdR/0D9hxTXThPn
qFNJpzXeqFPVCmF6Hc+vWXCQmnf1ic+iCa48TVp4vYVJMoG22pV5gZEeuBpG11gdokja1/s1BY9A
p0odbzVdkPCBJNQXIcgII1t3B1nC5ZE+hWgS5TRRX6vyudtLlqhIgvsdJ4KtjVkhsCRd6hjMUu2h
wUUUcVnFjvfYmMQTWfqDb9EDa1dSJl8C1jeV6QIsL2M21rZllzA92E6Km45k0JJU8yBR1+wFDS+Q
dmsNm9UP30Rn34mX3XODilDE/BSBPtbSEpiRUBZB0mlsMlw6xuSMlwGI1niyzQiP8y8iEQ3bE9i9
Uchq5PHr7jOXUlqoApzRPp0294A1NFlATOcNmfP68OtjvCTiNbktwwGfrg+treHD7ceWtJJFmxjT
qZ49RStQxR0l3TwckrnFICwqSyiTvWmaXRzwuVxJwvPtWn8kq27AHH4vrEtKrO2fwxcmm335Fd4v
o6Rvl7j3Ab0NCtzVOf2MhjWRVcAwJUwosK20VLe5P/Rj/nqdJUZxXIkmIpdE/FjqM8in5i0nD+GM
cUsxBpBkRqABSF2b5h4MNJLstPYQEEd6jo4JDLbwgSpA+SGPu+g1oQEKoIJFUb3hlxBlAusN9G5O
yVIrGsNfUU6+1sG+aroL5uXNMV1e7wWURpCoH+hhPlp2shA5uZWqTkWVq67TtEswRaRibAzDZrP4
1p5HgqIoW8CsaQ94KZf3BsBLgI42PGqc1zaKWx7dwwwB3TNl07wvXku5fywNu02J7N3+HhKu2Gyg
mlP8PwxTkk2M/xHdQl+4MUYFRLBGxkmdFe5YtjhNJXzpLIRGzQI5cNam1nZzNDVVAFGNzmqv0lSH
rW5h+ifzzzk/29Ex61DN+LmXny4YQedQnKWSNx5pBuh4n4/6CtDYmc+tikRfDzfzhyeGdE/QVjsN
w/KwOcmaPdIb1u2KX3EDsmpkijr7wWrqaBzEYgJGZALM4KOdhMzYMQKCGSmUw+SBoKnEFLy0WCbV
IlZ+dA2jIHgb6G2qp7hYKmEl5BEloeqgeiP7Xyvrm+gQEwR8kmzSpXVS2eO2H2v9eRsb2qgRj3Zm
azsYLd3yODG01Scp9UcIvW5kUrmoSLUl+FdfiRb/sEG9tK9+bCxHm8ZP0hDxqVO+euz163BqDDeR
K2AZKagyAoS9CSnvMK5+bBzKP4dfM+cKaB6j3FpCZVLGCGYzA1DJahw64hDr6/ZMRiicM7IVZJ98
UFhLQ6xY8+3PcXlriD+2u914laZwJyXyMOxFaXuynJZQE089rM6trsFIvWPkCqwj91lu+b3/bEaL
9InKiWBLb96YedohNU3vSNQwFBuXbIMZcFfLZ/MruEA6EqRV8WaUEC6zDE6aqTTJJ97+hbTs+mgl
zVVXiFNfBi57TGKz7F9AAZ9/wQAyUFQ2zomyBt90kFwKq7qp5yB66BHgiTTHHT5L5X443GwF1ZGs
mO2cl8AA0buLyD0BNxwE+tYNP0A4itOMavm24A31/0urfy8pXpJugT5UjGdzvvIUXeOmv2Ax4/7z
SQ4W62JCK/7CCpTu+RKDXRkoXVifm0z8vrYyUAuehLXFEdsp55OaPMjMwEa/vsDyFrebyVUHSclF
rg/dOKlLh83iQk4vEim+qwrco2JhaTy5GksXFqtWAG+9W4Mt758hAetglHNWoTntIINw1FFG457+
HYk4lD6SV9Y5m/OCKiIMGAX/Yd8eHtNXL0ysDDoTFNzsUAFFG9tvpLAQ0DmhZZOsh9jh3Lsi2Hw0
j7i/l7BAZ58CkzsWsGS+rZsqE0Vh0v1o+XeO8qwtSzaYHis0yc7QY9h3glE8eTvZ5oBYwAIN/tlO
vVDe2QTTq2E1g5UfMwM1oALD+0Ddiktn9ngOiTv87GFIUwuz7MwpmQI9udItGn+TaF5BZDraCJEs
1NhXtMQV+7q8L6Z3XJsbOFRN/HgThZq+qV+JEy+pu2ou8RhGHOdhWkAyFlzW2zC4tnu60QOiTr9k
t9IxYbLpQDeW11MQfvjZF/pffsnHQ0VpKF77SVjSwJOKKOOiNxVeMZLV7RZq3DiHCPckV+c0T7ww
Sti7kWNb8n2Eb42361d10aFRuToHQAoIIC96oEonodTrG6mDYLVmPi2HFEhppVqlpx9aTZLFi+5h
GY/om3/zcfLvVadzCUX1FfjZ6MU5NCN3Rb/2u5CV3v509YWpeQ4DRv3NHunSEW2e3CUZoqx9O7Ia
7IGDw4GkgD/93v1bawyA1a7JjLy8EFJCcL2prpdi4K8rlFrL0/T7fEnbd3kjxrnKIsRnJuEfhjsV
us+fOnvyx7qaNVtxDteem54YfLZDkY5Iw4ZyIv4LcbDBVHWTLVQhemzPwokeplG3MNhNL2c/aIKl
dji+fO3rD7BDAjhkseaH3UhKJIUPRoee0ktVNKUoqstwPTmESlKwBdR8WhRE31PRWR+VfTkdjl9p
dNmFQhjFVBIQrJabwZN43wlXTtyFEMyDjoLC9VyM0fVnK6n4ITIB7QFJ1vmaG72TXdoS+CUmiS4s
5tfExaydYQfHK/48TR8QZzcLXDJ8ws35qFdQKZpitoburPgdaFwC89MjGi75bPAQFsvKunqmvje7
sFFGcItY6yZL9JUx/oyVUupd8gqs3pXOQQh+aaU93ez+gua1wSYFYGNzuB5Q2MPyeW2Wl9Ce4ehp
W5+YsrqE9nki18nXQv3MlkjEcwV7N+sw8WbXe11ogUSgwtSbk3noZYqPfZkl8IhxVXgf+Zc284CK
NYvDQ7Fg93XXoLk2KUbizOcm3Ozipn4S3AVZZF9bluKzF8tYV9vLs5bVge5l6IaqRGKTknLRIf6u
lDSLkWypxM2V9SXmTGJLPW2ERpeX2A7qa1WLR9sumQ+lITnlZtKTZlzc366B8KKXnsiSMZAc6j3e
ko8r+zl3r5wLRNiqzTbMegf8wguHPOGYvmsOxLNlOmXCg39JfrBJHhxJuFrrm8B7X8fmWW8XwQZT
r0SKwPh6z4LrXEIrzJ/d929vmv1yMVD2mURnIdATAt90SO2jKrXzse5H7DaPmiDuIqdOrVhgt6PV
cB5DMn7Jsd8cl3v9SGRdzulkt/Cjy4LQWnQxkQ9jeiVheUsWTC/fLajT2fS7A5tlGRCXG1E5OYSC
lWFMeuKJh7astoM12998g8EbhiqSB3LuVafa4fS336FTc38gEQCep/6FreU8T/gjk8gV1fGp7J4P
6j8DSaA8ceQ7V544ZwQXAIJsXzv+7cwpnpQF2jorHGmj+HJ8YgjY9wwjGh9AWcSO2AYRLCHW3c7r
5aKEyYmduzvN2S8IdKRhyf2lGCgd04LlbR5GTr+WUCsQK91GceH92gEgLmSclqOv7SPxE+xtbUXD
TW0mT5bRDRxNK2yrKvbGXokKb2M/NCrdaI3r+Y0c2tLyaEYf8mzC/aYQz1aviBSB16g4TDo5Hecz
Rl/3ZrXjMJkvfa6W0zS2S5R9lFtMyFFe4RevPtaVjR09ehJfje8tCx+JglI1P7WDr+v/8D/s8/an
t3cDqJYrR9qjHwqEcqvBmGv1AMrB+xCWJR5+gErfdy6vUGRKOvfDiP9bOdFnQgU/zOYI2b+DMmlB
1v8OCIuqj0Bqt20xzIKfuTNlB7Pj2s0AzobMueGLuB9LiLzZMHAKiTtMx3QyXuvJEe+IjUCvMmr3
/oIjFkR2lw2IDhNSCWzWFYeKRAj1ouMlmA4HANPCbq1eMHo38nJ8agJMR2A0J0H5D2cwRt8jfhah
G1WU6eNl5hJ642VDoQgrtp9s+aanEnUarPVyVfyFxhm1IPIL23oSgpt50DuLF7RKK/k+isGaBVux
IAJmH9MG8iq3w/AtP8cLX97bICwx+3/oNu5MdjWrExUFqZzxnoeu6I/NvSwLJ5FxPtHbUGl93Iix
yjhcWdsA/mly9SB8xH4sZbIEEeNEDgAfFWttoNPbWvPq0yBnYarsqkvr/FeP8+/okXt+HnOu2qjo
RO+Uv1uQD95xjNHMGIoBNl3zkwaBKEaSPHm1G2M/ue4Zn/xqNKLbTtTHrKw34jupCvjYTaneL9KQ
uvSQihePlJALxy+U+vsUtUrOErauqhDcc9X2v6+L04FblJnAAG6nb+g1zp2VyjMRpsqMhDxMo1z4
onX8cJ8jTYE7hfNhiH4VcxwuyAPfrb2nkhMq1debNfdUW0PfO+cFdqgzkNKJyor4Z+oEgs+f2XoF
6FBUOmF2kcFAdN/lhMRV0XiMsST67phEZopDDuXgYVP6qUQTHLglmodcgBOPOPabBUXHXRttKXFw
QRvAapJqM9DhEEht+NWxoe7QKrlZSZgyP77z8rcuuaKMU8xNY2lRU4d6tqsdPnrk9U4y4uqQ+948
7LYNWkdFMkzeGKhJAe991Alzg3pfFKk5CyVBZ+SuDOcrDEkP67yiqwvRRBe9f6Vg/ufkz9JoFVCd
aQTgmOKhYbW+MvA2ZREql1Ezm+eNysSR9Hvrusi9cHR1l5ixkdm1XY3j2o9sMjTUw5r3JbPf8m2k
kD+1zZB6OWHDUVEJWGSE1dOxLcB1Zku4n6TYioy7vOZd9LpAHk56EBRLbxBT2wMK7FGjDICZ53lT
Ute1mX8J9uhXqoonVCXTeGqKThZNGhCGyUo5ZMNLRUycOvdjMky780VzoYJ2ejg/eD7CK2bhYnXR
9L4z9qxPVhEbm76ryeuKHeYCk9vsPrldwbVKRBgmuipgndv6m1xL7ESmjQqzSVGydMl3yvRGKQ8C
R+/5Fli22tluJomzkO2InGmJ+rXWZxxrshXQGwHfk8u4cY1JQCH7GlNZrLaHSk3hRJTpt4soVT1l
JiusFH2WMc8B08WSFdO3mMckmdjE/mQ2/lsZMnpJ9VpFCqzkpXpUCaoN7uHheK/fmW136Jco+ceY
CKjRQvBwOTZ9LUr8Tw71EF7HhmwqRve5XIIkihlQVPtXRUFqT5u5wNmtM6JQG04lU+cbuaSkMVDc
f17RjVaGu2J3GQ/gD/2PmGuF9U1CXOVkE1EIr+ako8HYD5TqiI6eTBuQzV85y//oLn8dt+Ni69UO
qnCEwr6J7MX7UMmcTaXkSdm3bIuwv645nNsPI5zi8LtHuWUoSfYr5eYZopaSqL8CaMaJaqHJq6AM
6EZUPAZuZHwD39cxpxfnBZ0VzzPHmEJU3iHdZ0G5d6sP3gqW9e0ZJKHM9LBObie63EhDeT+Md+Ry
0htH9YyT71cYSYX2zypwj5WlOuE0fv5i3gvgyUsZfbYmjsA4ko48BOzHrdc9m95RoQD2Fa3ouRgt
xKMnZFwZJvtn8yDOUkSrLptsnaBHinwswhDNpeiNjaGFfd4wHHn4IF8tL0u1TPy+P4TUZmMBX61z
IYdHujCT+T94HfIdfC7mlBhb7iazeOtMPmWEbu9XIGHqaVoX1nQFy9Q9b2QSLhFGcmJ71kvUeuUl
idGqB7nzrxl7V616xmEBf9Ke143g7J5XUQYMmEDhtqS8ZUQtYZkhc/Cc45NDb751gxNQj+zNn1Lg
uAT7+povqDawWghVWzKQje3cAKMs8+731WK0opzoRlKakaB2LUyOkq5LOMlJcIivDA+VBcvlrv59
bVE2/pRw7Flj6Hbeqv5oCxyYwgEp4j6qjWnEslDMN4LBNrwWwrRcqRTTwfOzdIQQ30y5c3MvwtK4
y/4+HIM2gzAMiIBxgwbKl3dEvzb6B+/pKVNoIssMVQbJcti3DNnl5Apdhje/WKZD9gjSfrgaia9B
tInjQO9kQWETwYPmzgKEht9xkhZaxsQPdRhl2YDTTk0QB35jAmYk002R8b+Qi2MVgwit8TL6dsqd
xod0ZO8o/3iO4pUduEp2FjBcdHEZwq2WnN3FI+VuwXNnvT4194uJ3ZgWr5hlaP1zlJpa5jL1UeTQ
t+xTw1xQnGreITQk6uMmuT/y4mtlMzFMdQPfqpO5yMsY/1DEcXERNeeQgMeo1iNZmpd/QDcd3vR2
nj0+Rhu+mmcUtAmEmkI1VUGruyX9Qo6ImY9+1EvO17HyL9IQYqZtUhxDQNGF/qgooaF258tOvr6Y
7haATxtcKAemOPBFkH5/5n7Nt9JpR8Ce5EUaj3YH3RLtu83OVOyHSxPfB/NKcrLSf+tmB6UpR/hL
ijuHLGw0bYKPNdQCBd+Ah638QyTXV26KubzHGi62LNaTpCRC6TWLugucKU2gb8bKFxHK+sM8IBfB
FZ5WoDdIwKro5XYRBQP8pY3qgR01zxEwidunb5cQEsbvc4tr5zI0RZC55Eh0s7Tm2ZCqkiNTzejz
v/ifrvYb2i3VEEc0ELeqqF5xxez2HyHm8rTUWTxtBgMj/j7l4Zqf4b2M7pTbbItDhTvpaoFffurA
QmESJCHdipM1kuvM93KoPEVHtwiMMyEE1X00x8y5NDNEkmgv1UDLnQGd/EsIX8f18v3nYjDj64AF
zYeHRv3lyeS6GzVr5wD9W4AYuzIOdasNgZUhv91ceYFrSsUSg3NRmO++3JlMutX5xC5qV8+M7tmP
m25sQIT8T4uSVZqdJsfldX5peuolEqF5E/xi8EfGvhx5cBjfVUivAZkv9BPe+a/3OhnO7rIeYDZH
T4FS3LF6HKSXfgLmjPirhxFCKd4cUu3Dz69oF0JDdMlL+Gan7uEuWz8BFCCylcyPU5AsCKRfc4LS
nYX+DbR5n1ibHvYfI83ed9HwrED1shSEY56Qi95rXuIh1qnrMB8daLR/GO5eXOcey3KAXmshUXiP
wPemqouyBAVu0ahcHNruYvSSHM1yVLk2KorCrzJsEw7iSV0BZ9rDGf1nS5LxWvKRMp/TmPdCF4Fi
x2jTrfcpkD+QWc6vWQpVmYQC48TeApfLTbfMzs/7gDL3iLVDOUS3n8N5IVymqFw5JuNAQPta3pvF
ts16daGE6awoWEfZ3SleQtIDV8YltXP49l4MbMKnqKn3vrtgMqa+WMMszKlq+xXAHImlDUWG7gRI
1ZX8t4qdMyZUrsk6qMy5l8E6SoymArBVM6t9bja2m5Q91Y2Eia3BoqZ5qCMIK6tMHL/1PDIjG02G
g95lopxEKCop+suZ2o4t8JAdy6ySYi7S/TE/p1B4Yg6mop1+gYQA2kszrKE0lIJl+KLBKcqXov1N
2EQZOIqWf2lDGzLZfUJcVges0TLlgJ258Se0Qc8CWcjjUAS0c3zsXVie2XGUWsMBOwws8XM5jtff
ES2zzvCA0KPdAMa4FeGTkM1wBDZxn5RKnnxvcI7tAVjScnRHdEzAnwSrft955bmazZZ0a07SHiT1
psXyX+Y1T4v0U3vPAwMeMX4ZOeFI8ctzvBevFZtaGXkT8nb2lK2zvWckMyKKunYkQNjTB5Obf6PU
70dLh0BlzfYoCsZWLkAfk0M4JYcy11tfdf6a7hBQSHRnSJvOVe/8dxIGqr633Sq8Zsztnzs0FtPN
BYdwtWkAJtjBNg3Gi5jtuZ7q3Zove6NUz4kiRgR654OCtYYpJTPvozEvVdLrOqrXHepdw+4/yFq+
ESlS1qoaeYc9OceEsKuCocd+ZYFuy3SNYHcH4WJHF2kwQ++/Ep5kZ3daY1IUTvNaTWTsKGqaHXpG
QESEPgwg0uzEw/OfYv+3AypCxh7SVJvg5hQ4uaSIc/WS7ioDVGaLMld9abWfT2hWPzEmcGkepYcw
6JhsdwBu2PyBHewt4nRgT/+u1u0ME7V4ljkQLzay+8orDfIJCjOh3NjtScp41uhb4Tfm5Df//x50
m5XPmxnELa5UzW/lbEeppzIHQUDn6mTo4ifR14PF1jiDs0zmxIQgeMm1zP3MTw6d3omTV1f2NYWe
xVUkm79vU+xcbNwK7lpnhCuAFq8o1SSwsobqIHY5GJ7ciC0Bw9qEXkn2O3a7qTai4XYYGs0+wXSQ
Vu+uOvMKETQVkCfw3+upxOarx6jl2FaZJDKuKY1QI0N7A9YLZjfzZViHkrtHBWdHUtgl3P8RXe6L
xb+e6Q3nRvr97UMZx3t4rfMafkXSkTrMQc625gw0NKeszIYNqtUKzxIdUdb2KNmzJZrZY8XbTYeG
8kRNB+8mP/m00qYo3izdNvCwvT315rTVFc8fHWfCjAzMATlefEqf+S5VPNDbTGcVWlcucGiXdP6g
FuxVcTHtAlB5AYhSDVue1AkMxhH7es1Uc4lSXDXpwvoQNQL0j2Vg0rqvU24+d0ygSg/H3IlmZmn/
AcyUr3ViwElzik5/VZiuUn4np5UwOJk5aPu070Ot87SS8fS+hVIeJmQqHGZMBpA1cmUZhjG4i+wZ
XRWv3K0Nx+cR0i6vuBHpZ0p0mBalKELQDDwDCoYtBaxfUJyExge874KiqFIZLb3JydhgnwBW4POM
9klA4b8Xa5qUxA2P+qWwMROLDv7fyVuBpkCZy6BAl43n/Tr54xv6bxPG6zA44Yetb5AdoEH8jVuQ
l+TE6Dk7kHIOyi9dd6Q9WoP4Wc+avT4WIm9pzCxvSp+TpK15NwpbhqIWBWUYSBCNilH0gUkk+wg/
OqWQtkl8WWsxc2U79xwgkNTXLSHdKGWPvzjDFS2MNDQ2Q89qNAROFx+gbs59kKgfmrEQvPSici4Y
ucYPhaw1odfypWMmncbUzp6wCFlmItoxa9ZIGJoyPZKimYeml7XdonQZ6bqrB4Gieqb+1Hk0f2J8
1LHp8fEQWsVJcYhaFP8dFEJ3IpO2cGT0Kjig42s9UnjRB06cGM38ckhR3VJZTOPmaHiEN7UO7jKx
fQOWsV8Kur0O8lhtLy7Lw0C7GvTkEJLFQUwXJghF66Sjx4NaayQaKgHSeFk7Vdpz+didvanj/33E
vHkYgSxhtBMZYMDa++/StflJ5ruRs3q96gyWVeckOgMUo8+p2O2GrDsFyg0hwn+Bnjx1paLFXl6K
7p7q5oLDUvYs0iNj0J3GUyy7hsOFP4uEpwCfK/XR6aI7alDIsLdUIksejzctSfjXWJ8WYmZdYKPV
S0ul+Ioi7KhaVKUv6SDKO4Lf60JAe57lJWOrTEiUM6yP2XILDuztcaoKwtDCzgPEPeIJgPw/P5EL
N3btGh1HDaj4p3QiheHqWbog3zfhbwjnfHNcbbFjCKVg45JcZ9Han5uZmKS9P8eOmmB0W35uwYG7
jhd9pDNecHfcAn7t0/+OEcR2345I4py+SDQgaTXz9wT2yZwTq/cqE7J3lTuFEWI2eNAJLhQvZDNs
7lk6BPLseEBQdDP6SBGjjemd7XvkbQg5qeyuMGHHSSIN4nSHaZOENg7cDn16eqqa8NUuUzgbWT66
JFCxbchiKViUcpOgnHIof8mV2zLRXgpWHsbJZbTCAeL5IxIuL0dE9Jy9+bS//9++6e0ymlCIHsVw
CTg1B31BYUJE0A2ZPgfEHYlk0EVmTXIi6RoQvtojX0G7p4Xi8HLLpwvz0I6IN41GIvdDK+USfrp6
mTPRjzjZYkXMNVG8ov+ITTCpChX/lRHgaE41U1yC+Wx0XDqE2bN4zGues2IQk4VesUIc+Xj9BmRq
bhJ/dAV2ykXBctHLY0y4VpPEJnQMRG5adZ+qdXmT0oijzsO3zpvGSmL75/7oeydEHoplB1H/QwTh
K3vFHi9Q8L3WB7ByRPkqxWoNnnGmzGypZzaIOU2YklQQS3lQpROUvDC9wjQL1MDcGcmVspEtk+9S
RBq/LNwmncl8jeXu58UCW/I4a8Olr7iEkQ/O0jbDhuu/CZRTrh2f8op0RPN2m/W7+OkprnAGIIB8
LBE/Yl4zdmLCWXdh5bKfiArpYJJlFnDLWaklUZMhwf5We6ypKGA/d1bDM52fVNAiuGxc5FTvOhT6
Go0qFnQhg8r+Z8VyUj4qFP897wWkyNx1eyh3vtlUed2zcFBvutskc2hLuU8+GyqLAyv50uM4RUqs
OLccM4+C0DAchGynp+QI4D5di4ykCHWZJy2qcckuHRja5gpaZjSuJ3vlTn4fc68Di8hA3gcSyKu6
72lShQoVRmpii+QkdMO19/s5c/vdc2vIyPNernov7+Q+jd8/CmK4CWiyS3rn17JFYpOrT/uRvbRG
AfFrbtiQbbdaHYWApEROh72z8EPgS57wlJQdEZjfK9j49nUg0Bemkw82XZaY7V8cSswfneajChOM
Rfp06qgOvkO0ET9encr4uEMmShZ0+RUWvITYV1FRqNsRmQT/LIRj10Z4RgPDd+9u5lm9yFXzjOl/
opq1sietsnXG1RkhcItnaEku9c+pKqjnEMM+ACfv3OXKmY+qAeX9FXH1dJeXs8HCyfogGNvF8TDi
3Mr8VICWuJzwJpQRcs6Wgazj8vUp3ExgMeiZiQ/zx2H1bI7heoJ/5SS0EPviO29EdjyhyRzV2LZt
5FH/85Z4Sys2H9nf8bdwFwd7i8A29mtCtjtU9wPGN6H+GlMqORCoipIz4HpYzYLNWFuUDa5ku6Bu
0ePnlVHfUmxhxB68nRXNr2pEj9mtnrSiIBgXBlWY+h42hJpmvtKzWUuyHlrBcpbKT4m0SI5ers4t
D8IMzATYdtnK9qg4sJBmpNMgBey6nGfCz+BHkzJduv4Wc7Jxij/G1vL/ymRuYQxs7iehpuNtkU/E
3hSyxTpRYiRu5u0Mpd2wuhzAKizd3qb9M+Y0J1IgfuGif8aaZJ3YO9fowcB5d1GtUrtlfrfKUp48
dFeu+7UH4FAKo1dqWzb28tEvbdDCmylBtiJsmJ3/QxqJahy+gGsXdRtoREvO55bphpU5MLICPPdO
TvKBmejyk1HoJ5i+5D2GfSzX/cbQqs5BKo98kx7dbns1a2saDwCg4zCVDOQGzHrfwq/xzBNpb4L2
kLhnyAjqiEeJJPx045G0WRL9PRJYfTwMPiZ5lFM+mzH9ELF4Df4CdamSimiCHrP/ZA6X3x+e/vGM
n1YcIG9ZHRrz4HdDWqEGDy7FoZfhw5BcxijCFI6g4cQ9T/Jv5Xr4ots1XNjxlF10qXrDgWmG+4dw
hCx2J+UHDVF+45Y55ZWUECt76Y7knW094dR2bVa5ubqi7nK0P/0w30AVgo9wMdcRobDAT0yKHLpd
vPDxiu9EY+T9+mzoHjjAS7wiHoswubSxSO7pS1bgBeKEB7rxIoyk7yIFg/3r0CztdsNCXi2W+u9W
JIZYRV4xS2HAu/rTmP2VF40SycML356V+sBRBxNh5fBnsJVw6avo7bIHcoOGIwcydCu4LWuaiTlJ
J26sj1XPabsekAFUK06LuHzmDFnk8y9BtXbuAovYBX5xo0AzCTaWfFXc4pHWac3xjPlLSS68K6WQ
qbPTDQBbV4j2V2gQo9c9pAKiX6p/KiHf9cG3u7/aUEgbJds3mKQpxx6gi3c3nA4xDzVUpJ5gz1Qy
eGv35cmr6yQr1o4krozGF50WnTSEyhzPV/9ikxDoyTlCn9N/6jj+5GQC4Y4kkAVj3morRL/MHiFW
Ppnao9jbOcFRj+dmGnqDRmMd9ANYxFwFuHCK+a7V+RP+3uUkONeiM2X3d5ttmLE94cxB7NXtpj0/
7O+9eKvweBQQN35T4U4crsCilxHnIDCfmj97P+3VF9J+nGfGaEg+ifsheeNY/Dkrz88HjVEydrvp
j3DRRg433jFaHwpzlRmIeJNpe5hvUHV+r9EDMUkrJA1g4iYR5sMg/PVlB4Wg298zwa3odcNHgz8D
zi8j+JeJOh7jlBoJkGv59BTX/hy8Lul7NgQMTvS2e3BXmXThLQwarM2l8JMNW88ijD3Vg4bgEFuq
Zk4AUhF8lhvvVnVbdqh2j8H8JR5ydgCUxR93opQ2ipYlxYHtYOVFTuJqcn7ht1GnGjSfqRTSDEi+
gWWgVGuefQv/3B+0QNhTOr0RVR3paoQWIQn9CqcWuMcDxOuN/XPyR05+FplxDjshyIhOYh8cHg2Q
Q0HxcqQPxMIcxEq61W76HTn8eoGj07+lgq4/T+TuhTSOgMFuJBMIk1UP51isaM6UG/G+01Iff67Y
bz/KduYrzdCSVQbgoflOL8HDjvMKstFMCqjtypoMRc+Lo3bkxfMl9elk2kmOge2NiS6gStsBFq6W
KHUfyqk/AIdpBR8VkRkdvbi5uMyj0kHzHUfiCpAOX77ED2zwmjvn3nvF86yRXiJgZTEzD6eHHf4Q
MIR1PDYfTWDDx8AUNb6x5e0e3iehf/E+QrEiNH1hbKLHoHKU4YGS9GC1Uknq2OPbIoXNtRXDRIF0
jJxxlLqm47WkBfh0xkmtw46MT+BCJw6kUlH5aT4paiXcZ7AXEJdgWpmJ16QE8lc3h8rQitqPP9GQ
9qsRsplktDgXyKGmEYJmYeA8+DR0a/v5sGucNx1m6GKPlLybjeav8qNcKvxWXQ4lmCYGEpCiHTl0
EJIdz4/y1vULX8AMirss1xP0Za+XzA0HccI3BUL06UixKbyJWeZnaU6dnDbTVzWB1pfLM7WoTZ8d
Vj9X7a1figC0RV+2cH5JnPgqecLslbhHxH+3Mgt3WUSYCtv3GWjaKAJpkXYi+gcTVpASYP8xSJvV
lTbzRqhSCP8GXRKYY0DHY09sDuREDSmo8rztFFS12iXdEh1cm34x29p2DNGJUeTDWLZoSfFY9fd7
z4OcUpCYfL7ErmQSFcGGUXjcEhhhI0gEhf7wEXEv8VIwx+HNadUwhDrBswusB+Rg5lIwcyJ1OAJf
PCFgzJHKbDj4S/UDOu2cCJX20OhdoOFdGL7S0IlmDIzjwe5kqUJXtR4aFAWG/saM/brMhkTSsxa4
ikuHaMaZ/EjpqjO78iEs42klZgHk/XZ9vmFAXXVLyC9evf6y31vUEkDPhQo6CefU44BArqm+kCgM
1CU+9QgGhpytPUWbZ6AMXUZPj4zReQlzno9uCYU8QqQ4d2BZ9jEE2bOPxN0f/wQjLVIlRd6g8IlY
El6goP4LU9zsAx5/YgCBT3UsS3/uQ9y4e5+kElhHVvktrQxtu53tt6eEPlDVs0E9pEJY/4LO40xs
/3gaLjgLw9MIOIQq6PQ4t8WtWhrHcHlNeagP4HqtKc5qdX81VtlDJ1Dcfty6lay9rbhdGcBfBcuB
d4j4tGm7LUJxClPzyvb6FlcsTTJdUnAfrcrhquFHd/Cm/y51pporaZlnMnD5Ll6Ns2zP6t7uBaNG
/EZ34s4z0tFjzxQkdoUR3fwOJ9a/MriIOWV9fsvEFddKyv9Cgeyr6MvcWZIEFVjNGntgB6bBXUez
7QVHtnl8cG1+pTPll8755gbs00IJWN8UOsGQboR0YfbsozX2pRokD4NtdrdPOd3y5Pmog6jfx4fC
0LlNy/GMzIsN+T4WBrN/V+aGLZhWtWBiio45gv4/tdYUNFAtPjeDiVIcf7CiiKcF1FbDu5URP627
BMAE9Q2vaF41MK3ZdWC5MOvHD2H0NHEd/1kqaqlP68SXKyziAGMK1fPTBELvZrpcwR63OIr7Rvvh
sh7N/o68yeYXyn/k5I+p1v+NotkCbugOiTS+0ypq9xbtfHTvviUfQ2fh/a/nYt/xciYI577+5amN
VNPlLLGxR3QzZalK19AV40wGyaX/Um811Z2bUED78ovZS1GhF0iXLAvypSkzwzwUaNLtizj9LsRL
uExmUrzPVWSQDlRKrs7o+U7qWDcUy2RFfQ+Kk2NihjOwoJVTOdWPSH7lLo2GdjY7vFvUY93KKoAq
EAhxQ1RNxAtw1oVRpBLLYEogxvZqs9ndoSCQgNJ4f0KmCvQQ8ICDNQu7aj9OVe3ukgRi/g/sIoOE
YRLiIth0SlCXfh0zX6W/VllDN282i4A7EMrY8EUcAsU7VKJ5OZHOpVCjalaNIPlyVKIkSRi1v6EJ
CMRvWMCMM3730BZNUsH5MKRP8q/GOJddA5jQ6WIJsjaH6ApGkpZv/MbM3L3bi/xHRSfcr91tgfKL
TkyCCRYzh7iUXwzWFdRt6AKtp9QMDnWZi4BADkLfk/AG+Hlpmw/M9Jl3phFEh848Sv0RFzGmCJfM
71h4lnEMbsvnZ7gmO5LynGqVz3kG1+pWSdcngnwVpUTqDvNgD060yUi7Y9psWpHnGySPT4yeWa04
TGV6yg5GEqMSvOX3Mg+daIVRbgZtSfwr5NTs/L8ruRPcHxVWK+kJ9LVZqXrjroJAxMkwOYpef47J
8k6vcaujAwxw264pkflztY8XwpyZ7QF1DstZ+pLkcBlkKFggd+W8N/Plp8rcXPBAfylu/OTuE9EG
0XZPwjVDfMmZauIJpltmPxTJTw2w7OBbGHRU99CNXXO0LUSykZH7zVQaVc0Og/Bn1kgJL85+8453
4SwHm0OQde78fcW/3jdqSaAfV90v/YazOB9wzW6n/0Ii5lXx1PkYKeIy74Y9KI4A10gVFfBM/hvT
zehkTA7nZ6klkK3Y9Pk37qJkw1U23q+KwB5z/eGhUAmGxbawbiWBzFM+FV2iPdkFq1D5KsGIUTky
u2oSTPRK6S9BoIkwvyS1wrEtiKfg2ub0jBMX3FURG82BzzdNP2x08tyNxf+VFo6WCdHJ5GyGJnow
3lMMEkrLmumljW4fqWeGv4PZG0FjcPWOHrCo97DfI/9Apmikr7sCKSTF1Y1FPcZS14q9uFZ8vU4N
Vhl3/hZn441w219+OrI76ZVKIqvuS+TLqOwbn+N9kma5FvFOpm8Ojact6BZdmhRNf90hzyc1wZNJ
d7ERGyAJQNGPyA+Amtre1PLsiHwcdA+MqfQ2+q/V//6BOLhnEUnGCeR23XBIIQdcfawVmPe3B09Q
Dde3YMcvhnxbd6aEClnwkTn20C9tbatg0npiT7s71Xtdz6JFBw3nt4WP1bBXQtogp7tUtPRNGM1H
AiuD2ewy0JWRuKOm5UoF4F7mem3c+xZKmn8vWjnUJgcEYZN1BdeVyOFL0oiDpji0f0/2S+78zK/U
Y/cOiILY5NcdIR/MPhMyc3J3en1xfb+ZjuTrfg3koV4g9BzIPyOjaCPxvqGNe42GQq4sOG18WEFO
9kzykhOB/P1EFx0HlAdEY/v5d2IRWru0RuuumogjCzH2o7TGCXlz6klBBUPB8YXND/AtyQfgaPDz
IRRvddFm950RHZm2/kX7zD54iVsAF16F3qezUvlumlA6NFsWKX42eG51I/5+HOCma/EpaqVKgTrD
aKqysxmf0YpuKkJQhlRVc4pDnL7Y+c75IDy3NWI2CoSxcGC3egvgtAC295QLVTQ1NBTdNBYVTB7S
BTpUc4rqLj0C9W6FSPWmUnNz7/noCOq7DV7LVmxUNKY4y4fqtqyxa60dN5BnnQbjBaWxOtW0bt/6
jW5eZsX6/Xh18gQpEC5mTtfwMEiF8+8IBBOp1GpMhHXp6JP8wuBNy422X1IfaUVnxGW5naXHq6IU
cDw7ikk8BsyU0jCUqfC0/WXaSdRwbvsmbET7Y3Vg7Y8VJpvHaIVb1YwLMZjC5J5OKWPY74WVdITp
QZePSRxrWPkDgODZTKzUNN8b6GdFyOxzrAZWnOC0jDvP0maACohKMh4Lxe4ZIIgSyL0mAqiq0HQH
ZYoFYwCYmrW5xflk+pT4DZ1OJq8IxnqLGmclF0lEcaywszASxP8oaU3g0Wzrpl/luFTQY51NOSTD
LhmSAjoX9FT68AxTq/wMGCOsSIKBbHkuEy3n4egw0iL0SNtBACJycHPC+8WZ1UVlJTgdHG8AaUAe
RLKqwnYx2YotKNsPV8z5arlPPbhW7/cjdzxv1HY9we1ZLFjCF0idqaNnWgT02qwzH6EuiYEEY7qq
ob61f9WdctW3ezGCAnk2A3DTmX+Sz95IUFeBYX8FH6kjGFF/JEOLjbXcdh2xeDrKXk7AEr3XFGyL
5iWTmFZiMx0Is1D3y2cOpeflY1m6mq9aoWqDSMNUle3Mkjh2XqhcYfnmS9Nc99L/WMZMJyqtfWJb
5qMilRpfaldR1Pc0iP6/SAN2u7M0w0lbqhcnc2l3bTNhlYIXcCM4VIQklMUK/dAot/dDCJnubK1d
uyCDPhXUjt3us/nqBnNw3VZHgqXGuCmbTmJRVXwV/ynKZRH5xtzjq3OLtOe7DbZHjBv+vM23YYDc
/nDvRpAEyPxvzkCJ2sJNv4G+XGegSoezv4e2wO6iN1qoraTTInTjufnBCJZGx+/rDWgMwJB0oysd
otWoWqDWIqNj+rIT2jBheT2PNEg9hfdzD5fPYSFKxrST/DI/g4GotoHVDAMudeq30dyO/kFG+jHU
4eYMA9ZH1St0kn7vvzwjxsLpZYdTUkYWISTLlCWsW63WdXrkYySKB0o99cdnRt5LI3RpxmII2KDB
WQ2gpMR/Zmfhw+DpGbMIpLQ3xkCiW0syDM4umELhrJiG3NFU2vGycyOypR1NbPKP6m9lvsUYvjak
FJmULRJrOEyABBSMZscx/VR81voU+bJUjnhnALeaTPEcAYFp+KDXf3XJln8MbuqX+Qov9BnEbtfi
JHDpjsWxVF3SFpDA+rr8NbXj57nc4jpzpkvDj4spwz6N1a4r4cnFOwNWPdEIljGg1/Qt3aAKRSdc
9KC4Yew2FaPgSgcGcXhPIoyReCSIS7ZvttcVlgf89/GDv4MYO6wy8gsfrzMqBfBXtnMfv1bpmRqU
aoPgTG0jybjXJ/SL+X2aPvew4UDuCEUD8UqFdbr3ExwwTP0Q8sSRUhUTIW7PZH1yPLyiswP17vyY
qkIjtBeb7YdjCig/rslo/oZlsqQyhbj9Uo5EntSUsdJBQq7y/N6pMAzqtG3TzcNUqMH7ZaZIPmqA
Vh5mXwpWI09baUpI3ggrXEX1ryVEbIMz2aYHELjhGVOfVp4DzQPuGX+Z0rjMmXuha4ZCkRw4DAvj
1GSwfw2zQMCDX3pFpoI09mbCc+qhAT2MI7Xtc43trD+gEkUCrk1rpUcaKPSt+uM7dHBzvfvRPkry
njfqq1nr7kM9YTVbBm44qgNnyv4piSgzDz2IO6e6c414y3kQF3CXvRlF4+B0t7uu4/yB9PogmF/L
jDCqJsBKSkBdTOHoSe/SD3/lW+4+OWsTaEgK2jTvlPda1+Us5IxVOUDz6uisMDC2hPVDnoXKoxnd
l2o3PnQDMxmsJEpCPt9ne/MdOkZDWw6rVQMR6Gu/KD3jKOmTfxHo4Tji1NIfyYQ0s56BG0bj63kZ
/q+w89WFljCg9rIqlqs1wqjPp7wLk0QOmzi6FJXGDKvplt0do1zFp94ejChv+deuUKwv3QM1gtQr
s+E4zziRD2K1BVaiy1C6UlK1A18/MZiOJI4w67ZujZI3I1izZPCJn2klsL71x1xebgq4vr2A3SPD
Q2xy8lidOi4lIdl9khzsvwHBOZGyU9XsjepnIC2dgftrMgIb7eVBerJ3RUhU88+44mMl3bR7VJDj
WNJO9MpZM6nPSFZwox6CJCtBVDc43OzoDAo3GLL2Uargl6kmDV+sWKeJ49De3pNtkWCg0NhDV/3b
NTEHihxrEk9rFPJP9/fRTJyHGTQoNW9xj+NXL0TIcyTbyOkvkpl85MvJ4umxOKiDiZDZypWNzUb5
SGnu4eBYkvkU2z4oDIlryT6An+PvXpiY7+OobnZJVY91AwdTHX4cKR+EOSmZPcE8SS/qqlegLJOB
esp3VbwcdZ0K1ebU02eW7q3dVgUOI/B3AdLsZtth9rG7by8vHE/WsopNYNOzxnhgjIS9WSRT8JKH
nPPkyz5/tW7du9hrkLGQzgBy1NY4smUd7G5nfazMFxydMFwbHkq591CVlJ8dzGoMM045Xxgp0IOB
9jLgaWvW7AkA0mh4iAajqirVHN0Gj2nmuroCuMbeqC7vUrQVO8xohFhmByFKesla7tHUplsiBXje
KBlQ8AIFwB8t3KzXPedLpLAuUgawfCtROabR0Gf0IK3kRGwMHMxXio0GzzKdbFQ6ECLkxghDyj1d
0Pcp0rCxhJtRXex/0I2V6jtACgFcLcuwtLnPOFdpgPFogaw0V1PUKgKwKdbRf5eZUgtt+8gHZqZp
yLIrp7wBeFm+DQhAOrw6RXCADiPk+HG9dOudqtVFS5JZoqCDVXGPWUYzn8GPbd0CpRYrV3Bfj/Vv
xkNjPvSAqsITkWGGjYdrpxN53xHG3T2ysjGwu9pxub4sy2Emp0+pzztHb6wQxAvQPSwPimAeHy4D
IwoTo/1xhTa0P+qitEVT+AhESpFlwQFI3ALbP6Vi6QCTapkV3L4L3ZZIxaz8TuhYXKKnvUdlZFe8
tozf3Qe79vlza+9TuK55Y02e52B5+K97Yfmk7y7ACstedbMIw3tzMeMg3quIbv0nL6ZhFJw3Dyad
uOaN6f7rkg8v6/RuoCkveBrd6BDYvHjk1irIDC9psB78AbNS7Dg9p7qG4NYZ/bK2kQ0lJv6y1LWB
O1jxgksmTMH1UISCcZA5qMTbcCgu5wgn+4qeorUbwactt+8pbwll7w336cyI67Q+EhIEemiwV7Qm
OXYopKSdnD9We0AHiFfFNmtfV7EudKG0M2/rt3N2McNpC9AW8PPyJOX8YK7P7XWIbu0ec6acfgB/
FcFLhKPDoUXe6tHdd0oUfMlpBVEAtAsMt0sSotH29epTS4uRCkOIupui8bXULusH03D/sV9y3f/S
k/2RAiDWTwRscTXwo6UNV3GHB9ooWjt+7evH4Cbafonbtv5hxeOGSvt88HtJohDOEw46hL35mJZp
kagaj8LOV8kBt9ukW+14CI+t2UmkY0cRL8TaRcIYf8y7MFOqUwJNda55Jb47hi9ZBEUCwzfPmRTb
UjNEXjo7qQf/cPVrvSHoyQZniu0QJ5NTjDfi3dfnyrSji8HLFhS828z56ctWJ/PnaBZ7KA7KjY1v
u+T9hTMfqBPFQDn26mkSck/yDNsjVlBxgmt+Gb1+9NrRcdEVMjbMrFyFqwmrSvVdIlsY4E/rpndp
//I5c20wW1PlxxeCNdzxnwo7SZ0miAKsrrlbjLdoQ2nUbcSrIk5gWp6qGYb+MReJbMmLlEaG70Et
om+vFZy1x7EwATbFL06v3yPJy+lsO6ipEKjw7OvktigSlleFw4yV69pWQkdrlnzkTybTWPMLOdo7
SAusY+WRpHucWPu3jojeeCSJ1Z3b3ojuXDmamd2nZxz8XoJDBVozJSpvLxfbNgo05I7vTe7U/OUl
83t0toQrY1VOmmwyxj6WLDuT3quiE01cF0LDdTRGxXjGLQ01jC0EHpSOLvIhs+1v/Dr60y0HI3KY
IHwUJ12Cdoej8/rD36ZtbWBl7t7JiZA+e0RuIWJ+tinIHa27w7/Aoz2KsPCnQ+UGBVs2frD9wuBH
bXBk8ndjA0t43riDJbgnXXfLCilPrIS+M9bymxtJOcSAGryFbwUsbA2Ff6vlN0xZVaUbhtOFKkGk
vPgN/HQSo598v1offeQ59/vt7fvcGg72D1ziegVKTEFNNrfQTgsIu5MPvFcb6jCudb17m1YkUGtl
GLdRG+Aia6peHJgEusE9J39WvX9OkdkjbrV9Egl8ybTSUWu6zz4V5n4/AZaipWsoNZBqrVPOtYYD
e4gM9jjOyS3Reu0DTs2lG19hFi8ElQs2CMe8VbHjlFun1jsArmPO2A9/oAwwwCQX5/1NxDYlv3Ve
G1DqOJRrhjFTQ6s3yq2wlsFLXGNXYq9EyBzwTS4xrMQvc20M2gt8E8lNoJ8O39C29kWRQsHCLoXA
OxGEED/pcPplr0g6xREG80hyDN1DY46YdFKvSvN1y7qu2nUO2Ucpcuf9yHVGG1DDy4c937/Aqkmy
9xXzaRCX3Y3cGWm/vfmY6yGIusiwhwK+l0qqfKMlYp5nLWyniixwrS5vSXJMEVvEtsifSwxV7+k6
vRvRybmURKmuT3PHj2lUgmokqG52mi38hsI7j2XEwOa2YX77P6a6APd3KzYmrOLMxiiCTafxdxRx
6IrP7U0NNQBOWVbvj2d3fK7HBhtxSlJDl4SgodOk9pQVE1l5sG9pwlcAkb5G7j8GnEJCDVahyfld
KJcuZs0Js3L8Jip/2BT/0AgX7Kkk8Sp71W9pt+5lhq98nrUaIhQvAE/VMl/kyObsriKyUH366ugP
i3HaC4eMb1szQ6edHW7X6pDobwFHeoJJupsS0k4IJzQAENNcnDZnFtnauhIlAGpqIleALpChUV6w
UdR8zYPL5JOttt62rzUO8B7kjtDXOJvM4VBKBURge0BzlDVwTB+H9YnwdVfNuAO0IxSMiZyypnnd
rxoUNaO4LtDscnBqYJqzMx42xnewgBadAXpELhEgcPhfvBLQ1Zcf0uPZLH1Tr8KtvZvlxWs+478S
eZ5/eIhNw71QJdk4kuhMqrj2vZR4xAFSWU6Twa1vnvpL4zYyhdy/cib5xmF9Iqz4qSDgShjZhZjh
AK7fMhyp4CvrnOvsTz4PDy8pM6H+5nBhEblYvFXvGGgnBNRSqHofVdtiVEz6NkA7ponUEKbr+zNa
u/f+//9P2d5KBjowkMw16i3HEm4A/HKSaq9u0v9t30lsU7sWphso5ZF5h78b+hwGC0LKremhA79H
2V244csX3XPDudYhIiFxdgQN7oSPLChciOXRXo0jdYO+ZsTgb1eI7xbCE3iTwEip9vaHlyoHlKiF
LO2sUnjV5yVUW3feeJZMkfoDKrsI6fEYK6Mc2rb+JJBgTf9XiiyIF5AEv9/37+mBjgpitZBXovXu
t0hswgJDj6v2TY3U12c+IImCSA3kK2jQUJH/IFp0vZIEG2hLUg2hPDNamZOaJSVL2sWgrqpkCdzd
1tkQOztC1bws2cSy0rJea68/r7vxwnYURbO6C9dT6YJTpM/Qmzv+tSapxEE+JY8UCyKudR6LqUOQ
zCANourkLK4BCODhN4uP5HTte+BKuFFXnDg2ozbWCsExWUMuEcDezdM+oum/d6ZG/FlcLK0Qe8l/
SoZZeSy6TXsH+LImm70KkibH7vK9GpaccOYzjX6BvGq2uHSlZ4nmtyjH9QNNsUS8BQhSVDMXGh+n
5gU67HjYAw79EupzEd5rsJaXF2uD1psIWY1J7gW8ynD+/6MId7b5+VIXLL0dJZToN+GqMQCZY/Ka
4p275u+lcm5fhK15cNMhxfZgAyzQeG5/ZIgz/00wsvKrP3+rHdvr+rIldssNjOMUFX4Tw/ZspgA2
oxpQ2Xg4iIBiT3v46F3FNRsbahx1N+oqyBNkeXFso2tBmlYbfd2xQH4OiP22mtNFOhBEMZ20qhta
YIzhEAzC9jM+2sPg1RAQxgqGaU5FnKPBHgbYd27I20NeIxjsbYyt46YJxxkx4bKNQXAH2O3Ql71m
iNSyUWbdHIVQgtolanwwxMKnbtESPh78q/PuJX/Dqw5gJl824F6naS7p3Q0vIA1EFlX7Vmys45xP
5tAcY1QgNlm7nEqUAOLa4DogpAATnqfWfsEzEb4uHRFG1MMx/JJj63RExZtfYdnaJucCDtnJD7UD
ulzoPb1WQo7Tt1b4DYvpqqHPb7DrdCatz1oKTpcjHwJyZe7G9xgJrD3tbLUSbSlMl1NjxA8hmffY
W45wU3RbeVpR0qBOTS/bI06miGwhChw5pPWyVg0fvWcUUsQxOV7wd7N4IwdOcfPz+R7e7Tc9XOHr
nmgW93Gobv7WovP+nl7Yjwm2+5Tf6z+7AmsTgIaJThdqcoV+w68r4JPmKuBHPo+zpCj4RIe/IGfq
CoQs7bPQbGnkTlOj1lOf1HHjMhqED5JEcFqWkxrBQFPW3j6iuKCu9oqsaLSBrgE/rkISCgulRhUj
YBg8vdr1FKmDm9I433kkS+bmE79vakKl8KdVrEn8M/uirlyOHhpItI10fL+hVzlSTtK8thtRHzHg
goQNdGso1DtwThzgwnemup7wSWb3y6O0PlsV1MqEx8vdYc4fYMoex0v/kRhgiMa81wSorgHDiaMM
SFLGNVYkykjgWmEqMIey2LlKVlCPEuVL63gxGoVZQcL7NQcoTA3QUjQherde6qoa/zpEs7jelp0t
xfEDMyKl82ZQYqC6n4jtsqrqC5IA9SU8MpP61Vof9t9x3DFJd4px9CRoQLjjTOSweVXd1b+jf4vD
OcOqAff3Hdax1F9DwoxSddf7l+CJrbZrWVBkIIJEp8oWDWeeaikf1sJWVdBI04fgfGwIxsQj4yRT
GwnW+Ga8V4wQ8EwRoD51TFsNt+BWbgB2BSzHhmHTkVGz3UZlUNtG3NCFl1JzBynQfFpfy5bkv8aE
x7GLd/Y04cPsneAl6RRNgHPQA0kB46B6pCH+IorwCKeDrewVQw2siqMyUSDPXU5n3ewQhEYHD+s/
svLiTXbJ7QK8ZkwTokivDKvDWmLny+8C2hagXvT+o+uDhM6LMCfuSXFYQ7HlBh+JsY8wM1UBTToU
QVZRM3P9uw3trMlzFpY8OPqRyp63NNnHydINbVALeGnJ8QSwZQvlpiQza89BfUktqXRYZKRlrm+Z
TwY/cR4TAySg3T8uy9RZZ381Na//GOW95GjUv03fzUaj26FsuTeWxQeEHna+WMNWh00lzmj87I8b
zHH2l5SmEuIs8ruHNYRF1GMBtiQ3Xkk1yzDKtkRP+Y+5l7fdnl3Re/zCLq/yrt0xKzFW1qeFA2iS
CMjRDtC5wIC3Si7TWSWibHyqV+6YTzd4YwYvxVyGhTWY+ffPsBBnyQSZHWHsXTnwlAXejk50RXDV
oe5/wzb9/NJF3/i3FEeBWeEz+0vIYsYgsErhK8Ou8REBGmGdDf+C99FtXNljoNq8d9ajw3g7WpGN
sdxwP8K8hMUCixOCbngk+xKl8xAmzMwxXgzMnsL53brwntjTtdvPLngQg1wxwRBJHjKglVp9PTYk
ZvrL9ATRyGHQEV+xVoOx9HKwIUBhtmvgLzBjswlDR57LcN27PgvL8ao1zJotB+3MOptdJUHdDohm
q3LvT5CpGgmGf1V71pxoJ6vqhbY5k7l634o0GiQe1ZMAaBcdA5h9CTmrhHokgWKo85qz0OwaNK1p
1PFKfPj/UKs/bLAbXmYYz9L3c2yAqnxcIgA2+cNw5qh6MARh7jLCEK3YaDvxsc1jc1Bhb+Nzr5t/
o3n5D9gxJN9ed2QUrmlLVlN3gclr5Wm2A0lzWGHjIZdS4/w0kxXwS3mqfA52FU+eXrW94Ol2wyYA
czqcM6COewOKCj5WOz8/jjc6FI/6+BWo86lqIixK00sxtFh1wIv1hfOlGmUSVXa07NrxDRVqrHSF
HpFQcUfvCTSygl/miqbL8V1RL6pbOZk5eC324Hg4S/Y+22n3E7NR4iXwwlMoVcv49guxW9VNKB7+
QkmurM2TeyXeHWHHNex/rQYmajWZadvaAcoQfNZ8Sd5o2VBi3oPLlRWLIqpV17S/iJ88LBeNuAgn
KBfui3miOLXX02uXAs7e9u66aNBYTCnYHcqZFx6X0ah80JU+8aWPRN+E6vAPliY6o4RSwUtLLEnD
ca7tfgzm0rE9Vp4AtzLG1AFIJRQax3YrbBNWiO7YO7URmu5gsz/aj+pGWVxQGnQKUZjsb6Qq6DEp
Xm4WIah5v2pA2GB9Gq/vDxzk9mPidkt4eQo5lqcIRgyqPxgiKHtL9DVPtovZVdYxal6X8PunMPZI
dhTN+q9tyeKaXqxWGpSTTwCfpoq6gGHRQcC2gIBKOabtotoP/tcd303IoN3nCqgnFOT2ApAhgmBf
hD3JIXbr8v/VqtgX9koEL5e+apkC2E9Ow3Z5GOhhN0uUWL4G4WVUI5Pkpn5JQccaERPwx3JurNJX
IO/qZrUU3cQb6CRyCcZJUqnh260UPa6QLgdF3a7LVLMgqx5FK7dnzHPh22ZcmuJCbvz4iMi8yFzo
s5AfetTDPGozsMh0/0OxDa2zhIkWnkZW8kCyrGUewaPJN5mampt4d+VQVJEjDcuLSY1EKSBhhkuh
w5uy/kye4IicFUaBPZV7rT/LTjYoYZN8BaiMzuw+G0W0sMJNg9pzvbWzh1KtghjX7BJSehpBvhwq
EpV/VVX95L05QQuQNFuHWD1ixl82taLCTTIp9boPiYGCMJ1I48sZXX2mNQTpeCJ2GliN7J++O/0l
moT1/MGCsyBJ6gZNrSPxAucD0/6YvMRhWKyjqOu948bkzS9UCdVCJYIQ0Wh7HPyOobFnY1Lu3YB7
z0qWHtKr/123uAudpRCbH+H32T5eQhmFW0K6rzJ5V5ziPb/1PgoGadaIN2GruOwHU4DdlnxIGEMz
ua6L17qa9HeI9bMFSXh+t/qzC+HPxMnoekCU4FfNvexCSElEGCuMjLjEY932UAA8r3xGnHRQ+bVu
NezkPZzLQ4jNvbfcJThIvBh8ublsC/FexM6Qy9Y5XHulTDgl9mz9vOSXsyZD0PFqflox9ilxgLip
jtv846TlGnffTxZGquTL+6qdcOTL79K4CG10uPNKsgtLkos1v3OUXYs3jM0yp32g+wBTtzQk1hLi
Ha7qVaVfUxhm4n9t3xhtKsxtUrxj3d1W1cS4RlXbFoeO8j2X4WIGogoeOM3o818ppwbA8J1sCrtc
mCuGmq3Mt6LxuZ42RQDSAiguhxzVxRyoIFjp1Pldz4rWufW9W2fUI/wKF6Hmq7nJHSF+wZ1Mn3Sl
8nLsr4jnHzylgb0NjWlxhAh5hS40/JM8PehxqqSsIVBupB8wVGnBuAO/Bg1s+w2lPvhiA8lMBRUE
K4vz2+REZX9/IDrrIOPZtroYoDc21RFR6MdHsHcQOy6sndRtKj4B0VfPzR9M3/ayVXl3JcgxVV3P
we16eeLAIamQexHSKrLsKvuWpidUeDUpy+WvP9ctJdQKrS3SB6XT6FrnyoRCUqYZUlqQk0O7DOx2
W1yvS0j6bCLWJloCVKQKx/nrSIAnOwjUkCYhrHhAwLZfBZ5ikwDWrD+WTavk66DwR2i0vSWhD/FQ
9O2eD+49meD+GYA+ozRA7NVMGkupXII+wicylewYzqOp1YSntKlfsEh1/9nxdrp6YeCygNcEbbim
nZW7jUjcLL5baaWoE7/D7IyvB3iLjB6Qf7guHmyWKBsCKfwMidg7kjgKphJh4Ce1CXSdep3Fu1El
Lw0avrg/sJka6g6BK22wgnsaJhAE09AWRqPe9BwSocDbvClfAbGQqHCYtcP5Az8/e0xza1H01Evs
4jRIuGCGhgOMaAhHAjLSK9xCbfzlGj5KGNcgGStFkr9iTfgXOAivSH0a68//S2LewvLeyDbXrv21
dqp2vfygGGCAbY6VGE0sYZLNonsSGqDwwGcBavNsd2M7JkIHrgv/1cm2xK1X0xh4adchpudyRRnJ
IwJVsaqtOU/LraHyjjpeoL+vUikfKjhlu+74AS4/NhUyL16scMPPRdqDvDuHeKEV0hhwqCvDCcpN
gfjioLwdj/PvSlzXMn1wSvAu3Zcp8+hyK+Z3rSd+lwpjuFJh+/i+3CDPj6wsKwwQTGyueVpZ3WCf
8lO6OGAv8E0ypEXt9gwQBIj12rbmIeybeYjj09SgSFKg1Adxgm9mE6bd4jKjTW5dJ8NwiNX9P78z
rjI9X5Vhe0p5PXcSVco6c1JCR6hnqmgxUWvuRWvzvDfIW2R56f3YZg5bT4qcUKvGIVA8bXd9P0eD
v4TbgeLqYoX6zliI76doMNKWHB/1jzVcVt7vrnyRWRZo21YbmS9C9YFgC9JAR3DJ+ngP5ZcMTNK9
m/jTZ3CLT1Rj2Is5LbTe1nCuYP5yzZrzDI5H3N70EnIHE1tFn3ftqdMs3dllYS3mwLAw3nk0DGIi
1lWXtoT4SobO7kz+Kfd043wpmczOzXVQpefqSD07ID7MxufNQbj+3X/ZemQm39N2VMX/HYZWdzpL
CpKJAxtibQGnIXRJfJJlmeyTq9208eEN1d5BoK/tptFh4MJ0McjDwT9EkSA06+JuQBfGez78FTut
XqaaD1TqWv40+vvSzWP6tibPPZaZT2TP+G/8vuenCsTrbpun68XkGk4QoGPq7jvTQr3HTfbkfd88
mrxVZ1nBtYct7TsB6KIJ8my8rdAnP5Tbf+ASf9XMvt7J+J6v/1RkjUjcCt0GrQ93lgYZe+iZPDrQ
YAkS6ftQx+kSsls/6yITt1W7+LhOykxl/glcFWpDBXi7dYxz8r6hJ3zIXr66KyGPKioVAcpchS3r
FVtKNrWbzhWMrLNE+FNpXBBnCHv4I3wOQ/u1lZofKKYdA3lI6cLgwTC8944AmYeRE9XK1jKzvu9H
AjRZW2dFX75wYnM4IIi3bHqL5j2RUBv+m6fgG5A6kcmzpwWBKgV5CJktDjr1P9bS5Odd15Igp5wg
q5xN6JUJoAN97kSBRuQkN2gnumXI8PAG8OEV1qSoc9qVy63CsojnXIGQgVjDupiTSmUX63zmujrR
Hviy3y5cKzb2QSVhSSAgifVdFQunKja0FhcmD/Oak0k3U47OBpgUOgMbAvsswC2WhI23mF2XXrkG
jj2/U7vPrmILgyOZknm/9veKm4AvlsJWtMjBeEmj5NP/331/bfR7gwbJ2SAFtK31qwT9z+EusCoM
+V9HKx8Sco3327me2KpNGQEMntpJgUnSQ51i09Wdxdg3iqbU0mRfbxE/IYy/YtMLxEw0BDL9CEjj
a1UGFzWlRFLWWB4tEyffAIwF0905VCTX2+c4eFRZDrvSVp22ulUu9UMBPKZ5ZWpmygUOMtiG+RxB
HwYJh+GlKGyzvaVGbwTEtn9vcGENuyjXtt2xFii4oD4iV8b6THOye+QwA/XApqbYfpXvDSyc55NN
VY2GSO8cSIADHk3Yq19K1X2Fd3BanwBso7wlKYo7YABKR7175cydhz2Hdr0Jc/qbgmKnC1qH6NVq
WoQiyVKVo2EoVtT6pDwvlEr0J1v4mHxG09fDQkv7GqddT80ukriXm4g6EvRfFEEz8860hLh3s3xB
Pghwbh/OASn5qxuq5frLxGM9R7sYCQHbxiNP61VHxSqf300OVJKWQMK5Pd/Vyhf2CV6Os9hHA7f2
RkyyJSxb2q+OBByEWdsaFbRad/g0XtZB+0+ze8KdGcQU3Ke6UiqNjfVyQ7thgeATWG9ve/JG8mlg
aDcTGELZe/9w86YQ/m353zTRtF7ADCCLlsK1dWi5yYeeuZNihUwtKLjMZivSojYy/uzGOz6QuI+m
UDYQFziDStQtLo2e2Fc46c/D5mg3Iqspck8zIkuXx+9r2kFp/DAuipj4fS7wkmUwnB+MD6AUTX4u
oXIgKNnFbIV4mu13NGcYunuIU7xBFBAPUemEQ29dO44ddA9sJANyadznjP2MH/EN/TeJ+DRXDjwz
uwwPEofLSMZUKGenuVrXS9qP4Xfv2NsWbmwj1IF6KaOCDMGje0yxVLAFgkUhqty58h8ZmCgBus0C
VIUavy4mYYwk4NNTZLrl3tZFJABQuWlgYjJgrp71cqRqInrFa39SSNW3IL4IIbmiG8UsQ6QUgkjn
zqjtz1iteGMw957HqnGrRGV3Wu3fiiDRmQZYlNQsuTDUkf4/1hHvZhmXD/VrXDgAeTXa9zB1cHAG
jKCmjnrjzpWmzCL8q06MLTtWBaSOMKLIesWCXGAPccHhDEe3z/vfb9f1XoXVCoU99qk5LDlaoRVz
gB/VRVNMswHg3N5U6+dXGE8/9uu8EdBvj6/boYZfpEsQ5Gh/l2seTVK4kMwELwqkm0Icio5LVmWI
tXJR12utQVB0BrfVSG7cXD5dawrWmfrzbdlMG67YMa49ho17ubnR1JiOClPqnauZ46RQ8M+eyOPf
PxH8xsQcdy+5P5ekscy+9eonF2FmLFKFao6cZpDWw7KGDY+ucauSQ8BPe7ok98xuz0yjC3Gx3BN5
mvYq3KqUy0v6oCXd6h4jk8nKWvJTmnwGKJ2Puc2kz0DhbG7xM5H7neMfSauXhslHqORtR5LQ4liI
5nGVBS/6anSXkuIpM0DqORW78sfJULjmYfEDQj0TTPlwgtal/E07nC89g8XYIh2fbpwX0a02w8+s
gNd6ajf9GS8STPTqJbGPfVmea7EI/Q4gDTZJ13OsdqmosFfO/xabF9hq6Y5ftkhzqUKFpxOmpERF
I9nKy+33JLd7aNnBkJdj4mtMfPc/G4f3skj9sIXQMgacMuncjOxIl0ICOoU5zItKO/3q5MmxPchJ
Pqiqhp8pr7KIlcT4tZYnoeKuX45LN5hOckCvMokVuAyjDChfzSOCwa0ykN32syda5Rb26FZZOg3x
otZWmxPJ4zyL0WWKi8qTOmfci8La8radijTDYpXCGAyxtr48563dA7r4T78hcqnu7+JL/CIdgRks
imKqwwNrxqK10j9BJ7gtzh+i4MMHpwxvsG3+CETjYjaPWy2R4IgSJT+afcmbt5nGrJ17gZYh6los
+OQ2n4NGCV/Klvz9vVZbgOI0pZly5EwRbQqondN85atGvqndyXj2VNs7GKGo46754e1hu8iajlce
wG9eDEX35LGHnFuFujb+BfqnxLYNFL4iDJypzx1zDUUKIfA3by1y8pty8d/DUWYDj/nHb1vf6WvQ
xuZpKyDm2TK99QdT/+NUtmB60fjWKqHZjlc/xBprRtVTH0aVPubABE4yG7tQVGdAFXhQpB+WaZ0A
D9TN3WsEJxOdMN+K20FP79xjiKtxldLSryYZ44p9Gqii6mhVczb5q5/aGgyumzg99ZRWiQV1SELS
007Kg63I5JDEqy5t6UE26hqbaijY1Cv10szAgczqF8ohMbwULp6t716RrOjaG35IZrh3y/L4xrB9
3TShUl5MDbh8NLdh/Cr4ReSK0yQ/WEBoibfKR58nrMecJIBxNnLLX3+gwunHH8c2zdtldUpti1GI
fypSnQbUU5CZxAE4HKMdupFw6nW6roF1V+M/wF0scObc9GQkN12PF3cAV5r8+RWBUWqJf0D3QRNp
NaAgh/JustwiivQpcMh72Oj5aA/pBVxxRMEhYhMCDmiFohd7JCKZFyNAs4iKvBU74CoHVCZ5ing+
yiYcr4sekpEcv2yRIjlPkfIle0cKSqRuDwIZkutnC50SWkXQpejxPpYZ2FTV0Hj83RszJT+0V7kL
skXzDnCo0E51TuSGO/NgHuV4GV8COdh9B8n12Z2y5z9JD7RkcFHH8nE9FYODKeGsSD22wtqmTqHi
/fYnO97O+rHKcR1hurCj6G7LX4T+iv9g3RlkvntNzzIKzEnCT0HuDFH5QMYUDnlSEifdrlJpvcY8
JqRPVV2Db/YSDo7y+80c0zgFOQXZrlHKoyYRG+i/phIVsDxPDMvtZjNVuCStldZRJiRMCO/Kq7m5
KnC83ceKrE8dbcXowFy0kYlpTnbaXL1WRFeaaPESBlnXCB18FAd5WXotEe2qnQXYELQgz+kQb/3/
x1HVnQDzYhH9YH9RqOPa3Ywevs/MuMYhOh9U5NWT9/cIw3xC8P8WYJmwz18ji1MAuU5e+iHAQOxk
i47nEC9E4bdeEsFasH9khgJqog4NAi0E14D8s4Xi3CTrK9fyae1uUDvUerWa/pPJw5KuQ/9/F9ws
GgQHCCiN/iX+VEaaKYqrq4IpSfUCzU3Zhxtu7XVUeTFsPESFY9z5TWCrvcIWA7s+RAd0cjiE0E8y
plE+QEO2brihH4MNtU3Q1aGmuatoMTmk+3cRSkyVSXRkXwWWSvlCi5PN07Zsv9q/EmopecLpqHri
QI4dqspdL6V4OazSKvUy50tQ3cMbLPPOXnmGdI7gXJfzn56DsDAmFr8yvqZXHIQJRWqGwTS9SEGS
T7xEX7IrHCKmz/kM4XCQuD/dLKVniyJM2sfNGA36h6PzWX/Qt5Ah0ZlsuVeliG94JKR54uKPgkQm
VUBzOYJOg7TsqJLD1kU4swE34LFb+iFOiQXCS7UBEX9N2xYyEWUrpSuDELQ271tfLl3ATOfwPs4e
lDHUhM2R6UDro1+QP2MvjmpQ6S5EWq7XoTah9CLd01ZADPCLPO4oq/QWaai4HpLgY1So3yszXX46
ACV7jTgebddbn/nUeP2Pd+B4YLnZwu4JC3AxObnZ5y98fuyOwhS7k51NZVQgmsmA9sCtPBF9hQUQ
ksHv9MbaIhOWhABzhtbu4S54gw4jKoaEI8f50IXxi009wiwRXmecw2LdcQC/Q3+PuVHXYGC3gXkN
t99GseZisTdDIAxU9nzgaeokBj81jFSjaky6n4pFRycxqVFtW85sC5CFTLJ1Egf6ID70PR4ghyhS
8YUwXmej6aMlzGE0jF+IGyzRngMvk1VcE3YObYajcS1x8DodJ5p3+zycHrmG9VsrwO+DdCPjV8cw
a3GQ8/lO6MoumiVCgULgaI3WUMyDC+7FR7z8gGOC/yks3RGpopcc9Hi7NGIuolon4pOg4jZRg5zM
wfl/Opzs7v5e/AYCp2BS+EoBUa541/hBqSn9UWN4waPStXMda818tfK+mhuYNeUGcg1xozMF370b
Rvl83LMMwVZIkKjLCIPZEFoqYAJrct0Wu3QDRMdluKPNjHWhq8N4VJRf6aaavToQ0COAByzOEArG
H9CVUVvVCXXgIR3SB8xv959u0Y45oejugLkMXo0LJAsgQIIAKmxZQJpgkUvFXPlL3NVevyv1GrfL
nzg95repA8ewELyDr71lCt4+RyJkqCVYa3X+loeZXwozbSPEYtbcjJXVuw4hN17JQ6sEIGpkHBEQ
fuwfmBtG1DCeKUUoZC2q89pti4u/P/t+KFD9OtEAoq/kW0Imow9oQzPRUKdEg0KqL1+KGcX/ZM9G
WQqm7LkXT4LLEsITA5N9Pbv026DZs2V3H9L0LxT9FiZVpy3+QATUE2uAQzHwgF3JlN97Wqe6lIk3
SeLz64zP2QyGaw2QSpft16hF6Lii0ivXvM5QaQvIugzad/ucvUVrgKk0GtghDLsK/bU2amKkEZOy
g8DimmmLMUe97C1bH8ZsqHg3NMiae+ZguYuRyakhyduLcR7Li4c2cys0qdxK+a9qNUW04Y+m9WZ7
8xKHnOsRR5WqL6iQkj1Bhsjnw8aQ34+dLhJzMo9bwloBZXy7Gm/1oaOB/kggGo2bWFiQltaImV0e
3vn0u6T4o5HUMtSYSxp0g4UJX52Jl9FZEkTTpx3Enm+dATbrqsFCjG+5WmmOyhx2vIiiks+1pjSN
TzWybGnFqWyJDA/uTMcbjzFnRE6Q+HlkmgskzFlB9N1MVWfHYeLK8dKYlLZDM/53Qrr6+1j3lJKC
SOH8jdtbMEeGLkbOZBBy0MSny5nDzkJHmP027sb8CVOXsUrjmJk9k4L++H15VDbx9hgBsDkz6wqf
0Qb5j1leB6nDxURgWktoLUK/lDr4SDk5J4FErH4Qr7uYh7k0+76s8Y+msYLpiuor0uSeJV+f5Kzp
oTH4zt6mzaEZTck6vd0gSzTg5ChORIVXLPiPkZsfKN4HCc/P1OnvXMqU0c2j6tt1CnFS3Nkiy/Ly
Q6rWyFgq09wlwSHCujr4yLXLnzhpptSkVuqKC8dBbAN49SqLUue0qMV4XxXGEPo6VMIUqYFEg8wg
WVofSl1bV3re7wh/yiu1UEdHDF5HR5aLadNFOYYVgUxduQTymWlYYB1Fpv6TfzwwFEn7QihlQx57
coCm+s8Z4hAu4/lBqQvncVHAPHM1gRlghNxvHwHC5CZ8Kr1+a+qUqY23R7++hD75hQtMNaDs/WPd
9ppgoU+wBfM3rVykwUk+HEi85neTiQBlJzD9z7nLS1vSySkumZ6PUPPTYe+5nVCubuB7B2z+Ho7A
hDFlVDPjJYfI/m/hsbii3Zf/Xf2UwQeFGu6zCAvW/zaJ8F592ZE64dgJlGwRTGpyk2+TWLzIEDDM
1J9qBOriXAe2Mu+FYiLpkxhk2dcV1xGcIfubv8Uq8Pcdoq6jxmgqSAa2CCTrKEwalZujR7UW/JIh
4J90eG0AYJxt6mMQFQGfsW6ppzpGJWOBc9s1eYqsiVYhSkHQit7rwZmAx4N3tDaxGel8cm080iJs
SxKyp/OSKFHuonSHHVBAXPjAzOIfuuGAQQqeaDi+ll/W5+dm94wWyS0iF3FrPE7anmw/yMXhztiY
CU8zSvCpymraEgEEGkguHsfPmip3+A8rY4o/zLorX28EdaAobSHDs/TA5GOstTvUEYpOvE+uoLWK
7DfMHv8UkWGZKfZYt44Sw5UQsLTeNPExkYqqIlyzG8fQAj29RvrQJgDY04n+CpxCkqWEciFmmdma
Ehm4W9mcym/t1kNUOimoUpnraM78O7kBsl5x1ko8ymxsIW6l0GKmY3hbyWNm04GRgtuMan0l4B4R
VAkKPbtvRBVW3Q5f0RrsPfN47fblKzvPPStE+Zqn/LIs2P+XlYhN+FW/VE8Opt+lPIS6AOflntid
CYZGyT1TCirxE+Mlc+ikt7qkKApg5oXD9uHnBHxUcAC+HA2YuDfN/D6O72PTeW0L3HpbcyQ35WDO
IX+sDI0hqHfzZsBO1Bp/P2myu76pxfSIebenAlq+A8dQIiGh0i1UL+soCKa2GN9dBCwRIYCnlb1G
B14J72urexVIfXFLETlMhLIuDb0WfYJrFwdGWJA3U+YCflzqbVQlVC64LSitEQfpc3zJthijLqcM
tOsnVPEnKjCPD51kJd6HIOUODlJm0kM3tZeFoTRprLC3jUll1D6xl7QqtNJJc6AhYrRcbyBBy1wv
VzNRDGyggr3G+z1Dd3x1COaoQ65bFaAoXMjY2YPPHPwrBIpGh+NB2FKq/LInpqqO9EXRroxBYjpW
LckTDs7aycy4cpvMisHOVQx1x1QTPO1K2ESdGjKj4pXN2S6CLz+0b0uIF4i8xMgUBZKgw8rXpFgZ
5ZgY4PfJMjzz6oTSVa0+osdoc+tMoqKv9KwjmCml1f7eg4NDdM6/5NQFSQqkbsXCEKXO+gxIPyIS
RIxR1LEzYACWWGyI9ccZs29Ikmb3JLlpZzOFIk9Wozt5RA+2yb0TO1NTj007ES/vL52es+vg25Ul
jTUkn+k97po7heCjPdPAiAKaoW3MrZnq33jyAd79L+rE+fsIf+QfgcgX9q51i51NbndFsmFusCci
lRmFFcdQ4KK8foAqduOeYb8casOaYJ7jHiy3jlr9GZ/031dOYFGV7NcrDdNQLH2tbx53U/eNZZ9t
rESDC4z9+V6weVYd9PGxPeebgK8fm/IHW2M50zP4US313OeqexnT7jiMC8YBgH4x8T27tpi5pj3d
pzmvHDdo/+V4C0HqLjlfrvA0NNPAeEXKVWJ3488b3RgGsPVc3RNrq2OEplJBWrC1IFy+Qu23DsiP
chrVxiIgMS7sG5rm9te81vrDiOP6+pJiPwmepiM0Z9EeRk9cnYurUl7mK3AzzfCXVwfpAUNa96zh
yRiOUvXjqWYKciJ7UxDsX6jFdySpg9s1UCBobWg8BzvPXMqpYofGBCvHkjrX1C/YbyI9TiaVg4HF
P48dn3V0Cmvl5hwr4lwvzY+p+xS9Fjk/WSHl8PmfvDKxMJ8HJMkl8cIVoV96BMSwx3kn8fC6Oef4
zWVjC5l1nAi0yE6TZgjyGXrTQfkM0vS5Qm1CgS8j39oduSfVlHHeKuNO7oCaW2XyRGd3kunV4/0M
dVsiq8dYVuu/2WuNkvRetXMkUA2pYUDqLmApeewu4/IMF3g47zj49IJWNNrh3Jp3FOs4m+mp4bQJ
xTxEbXhTM8QfUpHRla3Q80N8G0xBM48NXfdmFFylXoauK/Iy2RD1+T8iL0n9ShV9HAJzlge+wKGx
surupeYmL/IfDEz39K/MD+W8VFTRBrcsN+q7VPQJY7pIbGFEMsiritdSRZjpSaGch5jzzKpyOIBO
qYT4PJg5dUz5C8jRwhrXJ9OLvnNgWSwkFPtd22DTNHfUoJmJwhM+/7nmj9VvBVOxNKnZ8v0qZhtv
NWT2yRYFbDs6QxiF9V45vQUfnbx6fNIMr5SWbVvsWLyNbXmFp77g/gLRJyEjMQFTxovY4wktD4aZ
ANtxJAjH6+2LOyWJCIvK2bA09+8nlN6GxOr2AwjzJrMnwL2xb6V6XX+/pxeTTI5goZZ8XjRs0QCt
9SSHH/hZG029Kfcs6n3KkVcEkX372cRBdpj3i4PalcMXD9E9zGv/NBGrFUVt1BA2Yhb+VqdJgvxB
0K8jQpoqF7IY4Zxuisf9zuP/UFwJkuvU8X+pxk9Fva867e9M7dp3XW4DM7bm/+2YlxYMPGHA34OZ
aETESQTkPMTqdi08caCIdVIPlaso/1QlKcsVrKg7hMXv4z/XRpq1crbAU8NuFIXEco9rWr+TF9Fx
FXOMG/xZzdOOiNQq5Ppo4nBEw8CL/FoE1z7Niw6aNcb6OkKLcAgy1nm6B+TqbeETIywSmT9EzWAI
6DJ2RuGkwDOGlhxUbchzcWthE3ZMiK+1Dt19vyssX8jwQBzNsUVAPAGuXlxXkU1z6zsoxcclO3XD
ow7KyA3OGTV3ICU4B4j5wjBp5Zaj2Zil7qXPLXnNVzTN3uuFtCQxaKLMCcKfuiGquMuGOCmqVSge
v9hEwzhW1zfTgSzTbivEnbRQygDtxG2ubRdrhgJQIsskjvsG4EEyAYRwOWTttW68heJDaDjvIPRr
0lCg/GnoiJRshEeLR9bBzW3zeahG1EW9WzF7spJ3ot4tZulqWdVbdL9yVjt+9Gj3V2fgV8JeFCRq
UicG2OyHGmil/XEmCzWgtpVVJQ+LobMVBB0TO9ZFxmECj5TNXkifrzP/OwZEiiPeH/qEbBLOVddu
aBNUK90KBp4sk5B8UkHr4EqCLDo9JAd0C4QUfMUkVJ0gb/FYjeZgkIuzgeuBL9OuLedm0L5H7QL6
LV+EZCaQ6mi7nhx+gKL+H/RMjpJeYr30KE0i4bUKI9LcAEnbA0Envq2RLobyL6PMG7ZQp64uFo7U
QyaU2mODtj2Qj09QMOhkOTQj3qyYBesMYiC+nPSfJSPUcHYWzkyuXVqOINnebgwignazkJKnty6O
wr30JTjvTY3AK/wMYFe84gKauhpmLoytA9qrvJqV34fGPoULFYoCsyFT+WJqBFTkjHfVdMoBqmBd
+2Is38HvPRErL359nMqDXUozjxXpCh7l8CymcdvKXt9LV6cx7wQu6gHTQZxD5W2GWoFZlp00+Ylz
Yr+em/n4FP00yxQxUHMQUlhdfzvBY3Dz44qZSjcBJwiD7gVXyaoFYwBZCuyMhL9ZZliw1rcf6l51
Sb37a6+5utZoxwyRV3Cksk3LYNc2SS9iUlSW85JmcFBe5uqFVSu5pYfCZuoshevAi0yG4LpNVULk
MvP1Ir4EpSWdUoZorYK01mGcVOlmASPSdraeB981mSH7aDNZh5Zk1gG1KgIV1DC5VRhrGnMUmVZ+
N7zKyYQzEiH+gkfnHOkoS3lPSaSAyA9j6ohZNR/SglNg+qh7MlnqDH6jsWH1JsqKTGgKdNHPnnzZ
xpZGMIh+t54VR66Opa0awUjmUgdtNEJOCOKE955KW0V+VWAXrqhWa/kLtmZqDmnR+FUOtgDA05hG
yx7CXieVQWL9yuUyHyiwHIlKnG6BvPt1u+NDoVvEAH+skI+Gv6CO8YetWhkFayDtgbkJsCPmeJJW
DvwD3ITvMQG0GmsHTFxvO9kim61jPKx/aaUQN5IhO4sISiKU76+SgrNahLkoBwzwcz97C9uuFw9u
fWclTLIil1me4rvpitjtXCR+/3RZX2W5k85MS+mKihg1+dnUo+nTl4ZJ+7/B5ppnqP1k3KyWmMyY
SyGpixifDZcepyRrfCHSEqXDDL/aopsBwIxYv+49Xr2g2nvUc1BZtBZVbABFkedbFnBEcbheNw2S
QlhFvRoVXCJeK3hHVApNn6DOBIvTQKWDKv1jfu5kyFjVkA96uiHddx6qx7Q4XHgIgEj0Z8W4Vihi
jx6SBn/XU6V2Hu67Loba8oe0CVIJinx1JDYUsFUsgTuTi+F1GBN5BL6Tg/0kvRnQWDf+OSTzYeXI
nyzOBzoLaiYFIDkY11UPeUKaKf4mioMdJ8mBvqkAZRjtdcfsTDdF/G/itC2TgWZbOa8MAZnvcmsw
Uif2fvVJj9bwum8y6RArag9zrXLWN6Xo5Ap7dRYKJeapOs83FgvHzhAUzk0+VmI0Y6lm2iDfIZv6
kYnNBpMBXf0s2sWnp1OJx8/1G4ZZIXK9BLUPYnJn2hZS03cwvMJ8bfPXy6Xb/aiyUQJL2IbGmDVC
ijlr5rX3eVRSJKelLlX4Un9DPdLtMyoF05CK1vF9xnek8ZepAQUAYX5abfpAQEM6ss+l4LPaZAcJ
wm5/9hinal67WCQ20mMiQwmeil8DmcOnYTbt/mhhwTACUFnEaRP3Ldw+VYH65M9yYXYX37CMWd3J
IKbLOnjvtTrFz2n4Y04Tx2GEjo4YBxAlVryOlocyCAtk6/J0LcXaAoK0+j75AXJmx9ahbyd4q0Ho
MFzxhaU+/GXcjH5BwD9ale2GAYd1cV3RO1BE/yR9H77vQOHI5mDYdCUvS5CRyHhyXJrFsrq2XsvO
UZIaKDATxCJgnTJNxcq+zW/teY/e8dN92Fpb6vDOy/Ng/isAn9BD8ZyLs3vbkm+rZbDFJvRDQS8B
MD7WIFi5eGjpHtiA05eLlhtWFI9k0VWyLcVo/xSY1X2L+hKzdr/ddJqmRah159zHlYhC0DkbInr/
Q+L1piUTVNaXArOqJm1ww3LsRx4Rpz1zAIKK0QUQiyStJjTMkHYKPZFGO2Qu8BhCh5h1d2rRrm1t
uU5fv/dtUkgbKb42rocmT8dNrSWwmRkM/t0AYOqIcybwHgUqNGCeXD13fLuJ24q7lhmIwp9j9lkU
dTUAH+xG54MGpdqKK+SR1kZ3kEmjnX5042OGzOG5jmwEZT/MiYUCCuyQ0L9bAgL1PZJMokPTcGAm
3nw97BP+gMA7x96BHW/BcyO4FPdrGqQy1/+hnU+E2w57BR0JgUqd+kWJWcXXntujuImbW6+66+ND
a5vEZVD/91QiFKYaJv7RWTh/EGN9SOTcGsnDIduJWPRXQunvLU7CY8hVGQHqPFO88QR4aIU5ltfv
ErWJSJhP5Q2AlU/y1IZdSh2b3aqP0DyDTdwLEK8EOhRNJ3IWuPzxMfq5+/ThIPBnGAPpqCwNfZxs
OHBYBlb184O3hWs39VysVGyp6L98mFSXRH75l3roRSEigHTx1j2ue5nsxlRnLX2qddvd9Mq8Wgmv
BeRizrOz3VviRg29SQNwsZsAvERQHacNL5T7QyDeDf+K22DwEVJiBS9soFOHb88nPtF4LgJiOwdM
LYvBRzPqmbzTqjVyoKTlnHUGEnadV81zO+6/2hLDrmlBeR9anY5GAKC7vozPHb5yGxEDsPfNz8Qu
FIfq8MNcxefCl/OhzwC4LCh9UfrIO1/RlLNEyOfrFJ096xLIJpWjMjZXlmZoTpMxS/UKE1hnhmyw
uStZRaa5dZAUQ8j8wEcL9QbmjuXBh5hO8JQ/FlAvZmbwyQ3VA7zFaQGHOabl5R8y4EG1lLUiCDB+
rYldRWhsV3J8nCMh//s+EFaH6wcBNCkUB9DE2I6Tpj0tmhVEsSRrTP+0GaeYCz5D2pBft7Ax1KO4
TSdriniyvwQ4ZbpoL/o7HS49+EMVhsp6/1u7TUu44vwH2U7SC1wnvIgF5bTvA+i6fphgNYOMNcSu
jxAhPO1k9F9L3FovMXy11N7anEHs/VMyfWilFf+9U55Fg68OrGRaEByPaIPyUCaedJlVh2GuAPai
MoumJ7OJaTZzxzAeiYWHeyqyI9N1HKNAmq2aNQ5PvLvPsup0xtrzP2Y2fK4MoclGIy8p/WRO4nUq
Wp5BbrD7rkU2QYrfInpIHYYo7J4RliHs5+Y2YJaLohIb1o1JDhsPzZfwSz0jhvA1BCjJncIDA8i2
BZFRJUKaVDJPkVkexknD2NDy3D+hSv+Coc9NDHzHH8ChuXqkmAI7m0dZjXWVW5Cca1l4dzs5+TpF
mLDDyzcuPYHR3+Rj/9P7/Gelujcfxj9biJwObCtIMlwysao84r5n4Ku0wAviiXliIwkXxE8e1v7v
vtEgLYs2bv4h8+vGeyeQJ2gJ8BjFKDLdOzetZv36KdS9UDJjUXJ/1sM1k3DvPTJQzdZjVW5o6jLc
tl2kl0PHiXEC+PQSjLlMvhQNTGNdaZ8vv5+HFHNQGhuUIvZRMeWGzQ3qKAjnaiDGW1a/cR7RlnQm
anbrS3yOpDxNUFIgoho8SbnqNaGOK1xznG+L3u7oNucgKLgg06F5ZkV5B4s54iu9KssciCZWIf1l
BbLvLABjerynFelE+BAzwkj8ST9F1ID/ivZVTdCimrfhsLRWqWRmu2Gh6s1tZOIm6dwVnDwnWIQQ
zDLhIAPK5suW9GrT+VAilM2370DZqHRJvznXAfZcFQN8OtyBHHEQETMqybVhZw4awJJPRX/x1lr/
EpSsqUBTV/w1fW3G2Uq57Nr0MyevB84Tyosu7MRl8X0YJs9P3jkGJyzwa6cX8sviVH0ui5rg51v8
aevUWY1YMJ2VudlKsYtUNn2/WSHn9eVrR1g0YxVVlTJ1Ox9kGWRA8krqaYfzbpcNvF9H8eKwBOW0
avT2L9JIiNiOuRjq447aPFhWQRmyPvH6BzI95caZ7rqHmT7cyjUpGISrekpCK7YKa0NNZiEXPsrU
hzCKUQZCWyvtfEQLSP+xN1+PK5CDaCSDxqkyRkbEfunU+V0M6MfP9ptYNl5hcSpXMFIVPwvvAyIT
lNzLKQeCoxQAmaGq35VQtXTLdN0LTBVCVNpDkGfCJHrRbms4m9gia6BiucOep2/Dcwt1q5S+kn3f
ol6b2qAqqJG9c4VLffEflb/L77sp75vFERrxCY+9l4LcCXu9BydAAVdMcvsvNfHCdRPGSex/5/gd
9+hQoi+5TapI8yMEL6kJAmoViKLM7osrqBwu+rgBwVZwcIpb7WEHpVKWrxwybGE3UOWlSCFcZFd1
L6qZic/t7mtIYGDPqgP5XbY7Lz8BfySfRx+998GuyF3GZB7rcbVmw/LSr5xXyE+WA7eFFy7JkVC9
y88PQMZFWN6OI+LHFC2rQLlByleC7BxZvCtEvZrUzymT1lp7m7+anbY2BPoh/N9jKm78epOLV34d
6bfE6C4aKySCIBdoHV/MsrR4cP5lnM2CakyftvKdOnr7VqAsdo+e2Qit3p94W+LMJ/8T7oUZZ08X
ygUb+HrDlUrwvGRTnTQzcV88CuKkPaidRV8qYu+fCRgg3D6fEA7wZEPaNBf8c+IVNKH9sCXuJO0s
mFUFBM61IaOvbluVRg9qylW2Dygx7PfIFGZQfB+GPIrXKFkW0Ft8v0eF/uWsxXx5vCJOwU8xUwPL
axF7+nC3aphJqN3ztM5i1youKnZI6Nuhk/y7NAOUeQmNB1JcX4rqdq3endbJR2UiBaEa07yizAl7
Qo77WGMKBR/3bgxZ/4LE5HATclABA4GRY3ejqsLJf5VHvshcpXxdu5qlBwEfcv8KiivwXStoeK6M
ExsmKBz2aixs2qkWzoXzzp11lYV0QHL6tzy3hINu24RKjv5r75nFjkUd161hIliWGAaHJWNWSTD0
CCCFYmacYDJLtpVh8iGUhBsJECRCOZayTEM/Sq+o9axG2R0LUizTLrZrt781yXTpy/sVmRcQBvE2
wuRjJOIJQDYnnQXcepJcWUHoPrOHCYyacBLtYZ90s1rgduBMxZePeeux7SUPR/SjOnVUXAXz4qTj
d4YpWvZMCeSZUWAxilLb0CnD7WBbWJZo9oPkrUOuMhAD1afjticgETkbDxZjFmqM1ROPfL/r+uoy
PRIGdOMGEGZ7KHWFKRjSDsV2h/Ke/rufSEH8JJDxay5ZQYjyyCNUj3XyCkDkjjJSrlQNuaYdCF4P
1hEAWF/X96SXPwHxvyRD2j2Qso8DVNvr2h6AYEEI9zWC/z6eavnvoIFRj5EXvEz28C0/WWxlzl7i
GawGRqUpOeJZI6QKvSZzXVN5+x79E5kJxurPcLfs9S2v9M0go4Fj80dhO1yxNRwBCPvCSFqv5vWJ
bpgLXJiVq6fafEIDqYSXlGHBg8pRHwJSRtoeC/mJlQQQJDRyM91ySgBImXqCoLNJ2z2W0VgSdNID
sORkuIjpMvPNZ0V2JlyIIhHOp6Lm3Fl7BS+CYabxSMG4P7t4stQTauMOaTJ5BJu9BOCS4735fI9Z
mmbMAq6/QEYAyzp2FkDBBmku7buOPJA4Z6jbgPknpnW0IilI/kKTXzzJmUO39vMQOXVq7d6g00pN
2VW8lOIy1fh3cKJE2S3t1b8i2YiDtY29rTzAX3xmtj3rV86UPenkPK66IIIXswlF6sSA75/eFZux
WidKqcAlA2Z9/0WWABHX6whpS0MUsYX+p1VwYWDlA18UV9HHwcfeLGRJ3icv4ModVrJURDnFnv5Y
IaOWTlTJP2jz8+Znb6sr/sk7GOO+YWK9PgJBpTiUGI3YgN0bgR5/6OTuM97bNCWnJVo52/eEiTc9
StOvaWG8/AYqUT6hxBWaYq5DaF2rto5cO7DlMrBtAA/o4yw/NRrNk4PciBGoShy/wXpPOtKwoyt4
pGfZDJlqd15ifW6u3FSgIaTtU/KR822vNOEPxOFSUwV6zpU49if+z6vaftzl+EGuRcD5mbBnV0hm
ZxdGYiRJEcQWgcT8vxjpnoNXDU67H4YKgAQjnITjvnELUgvIE4UQc/VHjYs5UslWCKDWXppf3cIl
PzXZSE920Bkf1+/zC7GYU2GiAH9jLglbUGwdMU9v2xmxT+tWRi8+5/r3kiq94fkSN4NxxmPhloIr
9VMlNViC/QK/8aD16hMGFjnhdDeljbtnChoOaw2AXvblh+N3f1m8ndwftu12WuRLBSqwsCD96ONp
q7I2BVh6+bLbFlbgRsPNcipQKK63TfN6VEMRjM8dooU2tO5Q5hPWb9vSzhZPFJYXY9gFtFrSmXnn
iUH6lhQC4xGt8LqZa+P8WB6FEtBbUFzsQXjxw2hZgD3YUx+qiRZjeyS3/5vTzdPfTc6MjNSFI0nB
HlyhrPCn1U//e3C9pf78Hri4xRq+cm/h9ngNH6DDainuMcbFGO9oHacBla9khAs3pfC6qZyf94kK
PprlYcVZqqsibMGeF4Sz6kVgjKFZ8sxRMmnRqEt83fXJELYcVuqdKDgi6PboE9dB1vuJgAcmZCPW
C8tAPnLpGkTXah7rAxtzbcba9I9b2MzBOdG2zFw4h3Uoy1usKccjTdrScP4kLp8lwlsx1dr2TCRT
nhppOpBvPCtmNJEKVLXLKSqFPYAPt3UKg912a5/n12Ho7H8ih/IYpF6FskBy4MZjlCIo1TwL4GgN
qo2WLGsjo939OpKhK5s/vfY05Xc6sK/OYJF9wAubxxS0njXQUFy3SFWh0+XMsMZtxFxKgD1r6pe4
JCRhuodbPZBjuw6PEmSayIRHQOUzionD+g5x4zyMfvtsPU284ivBTc7W1mQXS0/Ome7Hnh2bISb5
kktgDs4d/DZYe7h/dcSDxSV+8XKP0/5VpVLcOWvcYOejVO08R5uuaK1TE8cfjfs7LjQcqUatWrXP
3Z2g9mFK0dZZIo3cJXlkc85LBvNYR92vOQTiivTRx4ELV4mHTszms0ihZ9gtq3tezldJ26rkPc5B
iJUioKgQFRy3a/+wWeag1R2ismS7w2xlsmEMcnzuQse3TAaFMdZd9FyjvfDZJOy7t8IO0ZtFN6oK
XQ8/TzNO7M8Cq3PVbOoc/aGT5LvrNpGwfhg4ZAwAodNnxkLw3yT+DKIqkDIXNHJh3qSgiYL+WY0H
9ukA/XOuUP0bpFGxKuSZzblZ1xdGxq7wi+LDwqvkAbSS7BjEaXWwS9xefSf13ehkjByuDtVTEvQl
aqpQnVHw8HqMwxHOHS/j6UPQ0M+2/yU0WPByvd/xD3lccfuBs8WrvLaZCPc9g5b2InWBWLkjg9n6
JlX9v83ysl9LwQqef3Uf6f9mVRssZKqWemYcdz08USK8ee0OIQoYd7LcIsb0qNcPIbXroxoHDAFE
M54XQwjxaJFo7EPbqwvktiLmTR711TjbgQGH+nXQcpO+JMkfhpcoL/LGjOY3aA7ftnjauWkSPQKq
ZASwTTIYjMN2dUcVDKO/s5ul4nTOtCwmywkqMDhHzivaIDgUEiel1FSkhosj950qcPHKZuqAudws
ztSiIZ0TPKCUq7QMpauuWB+56PTMh3UMWR8qTku8MrcGh9DHtbhmmqyvrvf/3B0OpWh5EK2lbhEG
z1ChVaH2StwIhiqkMujSIP2nbWdnYCl2vKNbaK1cbIio14boWOnoSi+PBd9HJcMSimNjeanp8Zyc
OaCGkgnxJwQUX0qKxOaEv7mJZps49FNBhEh590tmQ6nKABclQm3lZiaZaDxR1B+8a7/YVOlXQVYL
HZd7awaeEsxyPo7tV9Zlna7b+pkAWpt9azyVt/P3xzZccjpj1nyMWnu7yAtxu28n+05lcZfLGS0h
B1RQODWm7BIqqu8chfEJa3cHbvJPPxAIk+nDDG7ruKh6Aixjn+/J5iRx7jX3/EAdRJ3yDXjKHiKP
aKrYy6UjvbeGgfNAsxkmmXOkgK9G7Ja5MqDjiCltoA4mhjbFH+L7HvtdvmpmU8dypuF+hxyxLEow
tenZB+6SiD86ezY3Qm9g4618rQ0Aq+HxBmLm0lAbWaV/jr1IgIUP3EN1VTCidNbNaKl5dYG6TcVu
h74rNJS/l/m0FMbwQR//vXv18/kUywR0SAJmSJy/Wn3jTcOHFu6Stw+7Gy0kgYbU166RIi1eouNf
tVqhcn7XNEa148nT6DqQY7WuCPI4jnf5opY6E2UImOgbGj+gFF+RgpS2ULJz15uFKulW2nxznp55
cCecViIJLaUMooDaLrq7mldgKinJaJy+KlD8urArB2qbCwarh5OXQmWMZiQFtYYocd7ums6UGQbi
ibCprrfSiqGFsY8c6MsETpynB4FX2+32q/ryx+oGf2kMBL0KtysldkVY4haVa9MOcUfV2cbhWuRq
B1JkSIsY7ubEbufUNb8ShZCYs5X9Egdaqy5f8j3w9S88Vsg/A90Q2hPNtKPAZJM6g5W4T2HeDfFh
91LkvWTs3bW/LDAvH/TO9Ibk4eZEqQwIMmQvzzVc5GE8eS+Nl2V2mArLPQCdAxMIavwSBVDckou5
iDtUBWq4w7iMVtbZ1RA/UtHnAH7a4/lGPDXsyTMZUWmSp5vVrHlufQ80goAABi6ab9AHPVeS0CPu
nU7ISPHERyuLR8IRJ0GrgQ/7bO9DzVPNbusxct3+sFBlvhxzWgCcP1+sNjRbk1eBTtOQc8i4GSVK
Mc0rN5EyWjZVeQm+nMVxJsEP7D8QdDOBrqiwzEQjGnry8DxplB6gx4tgbESb+/RYresiF6NO2emC
5/UBeRSdql72yv8oTPGg29imoQAPQD9kcI0E2D/iIDY13VJumzPeVu/7p+0pOdWlDGJjQyfZaXz0
CHDz0e9jC5P9D13ZzWMPx6MOTKlfmw82hgIPM4aXZgWs+7/UAAHM7JDxuOFPJ2Okjx3FTkyBPwav
Q5sIht9efQ+lSsaP1pI9Qdxy0zkhBXBNgMbXYvzNTWEOo8ZnKwqtiZtl/CmVfVC6ji6KEqY0gZ8W
m19TdBX/UegNEtFOKy4HKYq6O3384Oyc8wAaLBultc846m2qFuyietL408FV5A+V1rLdZRUWuu0G
w56jwrxLacd1HAkZaPR5Fh50dspX6KbjvKDbHENKOBzkve5g5+K/UCE9/bDO/3menuL1ARz4zpnr
ToRAVeH9m5dcXasDUaIm/8QFxUhT//ZoblHkYAikigph9d+GqWjn0ouWylzOWthTHIksrAyZ2RvI
LJqnvDdNTyGjlW+IavSLZHm/OpzjOGTnqMZpdRLOFlN4MD/hNiJj/uXA/CtmaAGeIJh6VErw6x9j
OyU41UkxoxhJCq7+yyr7ceGRuVGCFjKLLqfeD3C6gx4QLIJ3uC9kPZnGrIotrogwbv/APlijPDpF
u/8kQHf8XdPT7AhFg7gp5zEKOIoDsg+dI6x/2cK1FtGM0ApZfthKrIwxTfrkuUOSLB610QGdr4TU
y4Ep+8XmUDkUaheeaxWMBhdigrm4MsPC7tYwZs+tL4cTq8WC5hEeHU4RREVVpSavb40Pdc5kHHRB
XFErCPCrNyib38swvks2eJ8KIzr98yYzQhpP5aquHxOwn8QKSY/hQSsi9kSzd/mxNqMwZE1cyle4
K1EnwQnC8g6qhm1r1t5eiQPD918ed0zluKPg0M3pFGiQAWggi/wLCYt9IP1kXxJ7VY3KALFKObqr
66T52OAX7h85xg0wQ3G60KQloTOP3YYdUeglrV46QMNj/ict2i2NWNJvxV1DULOd1iJNLLIMPOMn
XfSNWiy7StlgJkx9wIGMff23MrjSeyHGy4bM3cLBogbSrCWcDmdWwHNlEBHI8l+do1ROlxwliTT9
33ICb6nt4uyuqebF8i/pcDRQsDBLTIrFAM8vIZLGT0dXelg8Vj4YNewXSfGfq/4J0PUdLuIFMJEo
ENQnvLwTXsiGBgbpSA9RjxwBB9O65jWhQBa8laJgaNgrXeKtdiaHBMUh04djYCwKRi9m4+lfvCXT
/DuhSDB+2r389ZTEejEuTqWSWbDaE9SU+q/hk4f8lQBYrdqLno61mdX9X87NmDeST2O5FwBVpxA+
NmSHUmtL0af5cBvBk4Rbpsd/bG0/6h6B0xDOWXUXBCtRBmXRQiGYUgGfoYI7+DkWCcbGijMMTTfJ
s07GeDPinKYDakGpbV6dXhNHoehAi7a+ycmuejmzM44qPYAsUbxnAcyBbUuVDYTUEATIUGXAvbhe
oQIOmLK6Bmqabg7xhlZ6s8rFzZseRwzNSvr7tTnluafiVxVpp6/stkPl66pbGr7EuITmsLrQr7Vc
YsX7Gq3T5wdgFzrHEESPvLXzBxzkU9Xnu/+S4f2WQBqvt3Q5hyE6j45vFDIki+V0fyEYjUuQY3nc
kyKXtbPSJQvfFNO7bF5WHfr7S7zWrnbgG5lT/AnAqq++b0oYe4+bA/9zW0rla4CnowOsh2uOEWgE
wUqVoJDeWNQ2JEIVC3pc99UT84FGnis93acg8M8SngC551aKfaG3YExAT8ziqMRFC8VNOYppdGT7
ulc+RRB7tKdYuyGe8pN7cOBOEtR2dgGgQuZHt923wc/I0R+RRAU8ZHQSdhbIw7K0PeEnJmpnDJa+
d2SEJPD3I6ODzyZqdRJ6SxGXa5eBzmCjrQgIN6vGl0OpvqEhLXl3gVPMRHqPawWu/KccHNGwfgBj
LZLNVvK4CxzlQP+i7wMgYVis1SqC2+szGKrlaenIWf9nso/nVCJz9y7mT3Oi8CPdWd8P83mpE6kI
U1BAQHbLJMkmnL0WsFVn8ElN7a1jJDKdZfVK5n7ivn2rgmsmV3KW5zZC8DcH1yHEZen+IDKHr3bK
czs+8sWSVIGqZUFfok5RZV5AUuQOm/2u0/G4aMQJHGtLdDNPzv6O7dbdMYr4u94ZmkHmQLC3HJA0
ipay2reBfiCSipZfnIS9AJVGHVJZdLDFrgcFyceNcWqNZFWfhhFy3c/uFMK6nYjEp/Ac6Xc70u3e
gYWhw5yB3rmKu3+c7SJm4jvrDk4ZhC1srTF294D2HT/KvNhTlbZT/d1Snb14UtTH8Qo3OCJBmFly
ag9R65AFS58xzYMSuCMYq/BQeYKCFQhwSJD+TzA/8sa7eGtG5AHn7x0ZdBlGzCMqqyMSCN4Z0/tO
jBfUv8c3aPPXYLGkijJH0SNFQlu22KqAXQIK0uydfq1Zr9NIAo/aarYQxTTagxxl+/wUE6A9le13
M06ikglqBiWSFm/69HLtzmymZnR/lZ9z+z/aC0pKB9REaQ//vTJ/KcSkjV/YgDHyua+lSm9IUpKw
KuprdjHS7gdZ4oPt/g05PoV+dDNdN6e/JzJkpPFdFyu2SZxBBKjNh/N1JHlEVXe2PkrIARfbWzyd
bjj6IfDawGuO9ZhemYMCdnotW9KNy3h1Fle9BirQxJrHK4nhbGJRBJeJXKv+SvkEPakZRn5Js5Wq
Dd0Uioe5h1+aSk9jtJN1Hz7kmB+8UtGIdOjOCi9Kg4zks+LNCG1aswEOBXNYlDJFxvqAWt1FGTEs
8WMPuXfVDtN2gKKP2igCHTnjJqoAhorxYV9ISlLFgRBSFQH7anM6sLo3dMAzmNGHVw73TuR5MYJZ
GIMpcyZUhmF9ayBjKbKrWuvmCOr8eF0gBWc6lbdd15BgqaZmvyyi3YmRG5rWkcwLSOL3kGl3mcj2
Uyd2jdJLSnIYQz4eRoouXLVFtTe7bcQWN45X8n2Eokwi9jFomBuoEtceUcxwVW7x0bH8KXuMPZfj
hHV+IE0gIVoWbAmvKWKijeQ/LrWdHsdryD+LXoEKax+QNTn43mnZlVr/hxYbIQs4zUEsK3xBuacJ
DpMwwOjFHDSL3ieLBehh89OAfBDXNTs0FtcqV1IdtTMj7l6ynfSm8XOkXKXrOw0FCbYn3kKAiwQk
joeyX+QMOp+3KL9FwVrPtiOT3osHLFOta+fzzewXpHakjnH86orltZxoCUnM5GJ+kaeoctCTq0xq
RP8Z52j5vJOuon03MnnFMMsBbkDAI0OuMH4w/723HEKBSWaLECibXrV0Q2n6x/sC9iyxqDoP/l+P
qRPtrOIOTjOJje9ARsBN+bMXqbFytD+UOfO/zpU7tyy0Pr/GYIyfJI3JeMqRQX0Jzim3O6KBMD1E
XXlVbA5PuHxFvT+G+1MTfOmY4l/zLy1Ul1iNDu6JCt5dXhIN9czRTTUoW+x0Lnxyxya10+nf9F/4
Jp+QWgRxWcWA8VJ3Ab2H8wICt+SU0431Or8D8/Qeg+q34cCR5TdvfSGjT8PF/a3XQiNBrOwsCTRE
MpKITrDpG8DoZoiKeRxCpi7Ov6rYLsZo4TfeHVtGym7IBsekju8yrRSCC44yVlD/V2Nl8KXeuc3A
MunszdaKY5D2HAf5Gvns22uD+tVOD9Brv04wlltCEnc74gWi9nXFPXHDFzWatjqWluYzLS27TBmS
CGFBKBZP6wzbHFvE08ZpzA7yKtBK7oQDxovw4KvRK/ErJldpvKXxggSLVi0NKAwHexJ9Rx6Y7Sak
77X6FoeyDTRCE6IWWGxJgCsiVruButStv9y1KoQPqWFDZ+Bua1UiVdbSiwg+NHCslUOcEgsrPkga
NJTdftnCiD4LrNbluURxtU35Pm5+M8PxXqaPKN1cqaRjN1JQotmh4Ux3ZfjK9q6AIXG46P3qws5d
W/RHDsU1B6+Ct/OiBngwvNyymNWTTtkbRE+svVupE6iqQXZkUP5VoDwH1kXqQhMr+u4sNRlGfJ4X
KJggXQRgv4A78bc3T9c5fJEb7qljXE1zQzyENGUmmlQbRyQkmfDaXNnjHKZy0fBR2PUxcZDUQEy3
QvEZHIO7cf1ZxIX0rgtMXZLzIqmUqVVybU65OxGE5qMUn47WbdUzo5dNj5ichpvYKxtYyoQtGKIQ
r/TDjED9bFCS2TWdXVDgHfB+m31NwOJS9H84rRUJCsweqvWzJrP2ql7VzoxlPcRIIcf9sDxuPftK
kfUZCb9Kx1VTiQeVaHlALOaduqPU+hebkZe3Bhf4I0khTpiW71qPDQHh/WLDVekMqoHuttMcPw+N
Wj0FDYRkEqxyShtTIBphnpM7jEsU1F7IXKJY4pquydhTjtMh9OooBhVjo8y0krg8Ff0VK9dxm5/7
SF5pYx/h3Xt1/ChM6oWkH8TVZDDnRvFZYo6mjmMjxwu1gLjSqSzTkq0Knoi88NGGV7n2XNxMawBj
qq6T6OXb/HEh+TbcclGP99N3gNwlLCqh0wKw0bun05WjDduuctm7Lw0LJ/iUd/Hq1nzbBhnWGLwe
LqUCsVaTVRZXeXiK9+t/561xRKJIcl+ZctL6nXApyvEFMdzePrtcNrGda32qZG6ZeSOdvOF+IUnv
HKjUK7q+GqBeU21mtVBUzikTIdCkqGGcasCeJzMDWll91NxMuS5FC4VgVHah4s8DEi5zLi2jZVIb
YvuiRX7LH/+2vVTwr5rERLB8Bd14sbJIB0i7dFRb7rJSVJFvMvMMHwP/LknoQmtcOijSLu6VwJ4p
13Qun0dLHWViDKDn7XKfdW5KaYryqOvBer3FWrQ22zvNNMTJdbBNjuOcgKXS+3G+4JgUbEeVnJ2D
29A3+uwE9gKZObMzbiY+32oowL9ZSvUFmL9MGLCHIBpX2da4SVJNmadAVXpfmgytFy0QNqHNBMKl
x0KR73CovO1xq3e7dGF8cqb+KzV5Ci49m9Ayr2VGuL1XXsKaqc+o7Xg83khOtxH3ahXVio1sEEJq
StWE2VaOw44TN2M6TUD6PuDU6Dmaz4hYC00LlRNyRyZLx73gUBZCG9y5JhozYDQUOWoeeWsNRmyj
83rvAWZK+A0mUMRoCiMW7QA7TDf8qyEPge7mb6o3SlFWAtSNDERun1KZFlonqHPEzApbfbo+XZm6
XsPIoY2e3TwRASSsfxNcj69J4smY1qW6PO8r6CIH+pByKl7Q2Y5FyB+WwDBpRNnuycxtGO29S/UC
ftKGmvhcRbL+FIWfJLMbCcph94HV+RiPLQSxBBzwGfMS0KCdBccx9hjJyQuDZzRJcZirBFAbg4dP
zfivUvgXKNGoa9z5iX1qQ6UJ8OX9i9MTCGp7vYvvsYVQcYILV8kEFgzeO2g29hNWmVlbY/uSF+YF
t7cBg3mqqW11KWyz+qThj00GVrf7MVPpp2Rli4AD4vDYRZYsEQskaJZf5d7k01j1d43iSmqtReiC
6ciO+zkDj+hblbIJSMlKFX4oX8z/tH9+UebTbXtq5QIzYXvsxpjRrzONr4LrzWaiyW++6eJxvVLT
B5BCFkB8tBkLATuuTed4SGWj8jRgWBSb5sLhAXgmJVoQ49G4eV0RqhTYAy1MzCoF8obewy3YiPEH
HlwNpedVTQtyOaGXr15HEOfYu37idnja4ZrdMq6C55uCzF3kamwAwaBzjg4GKgNsnL+s1M6iqns0
+tdex2z3qdTA+faIxWRWUIu+GVzM20xtMX6nZU7re8oLvTPKu6MLmzshADxva/y9QpXmBZiRCnyc
4cA1QuQOyOXHUZrLD7cM0XCbJOaQ6YDXMP6WpdiGYU4jlUDnxlOUD65CLmyG8mhukAAhSi40CVwo
V85JNSaLC8MeflXbpzMonO4JHL21+yJVHQiSmRN58GHRH/A0Uxkx+JUK3i0A7Okra5+cOFXGDSZw
qUcMrE0KzpMrOuviamCit6h4MZxM59O6D2NgNwrmIaC639VonQCipsg+NCaNvQ8ECykmfOTKA43D
UTXqa/1UDIUYrnFsbd9DRB36HNu/QAezrEvhuNWzgmjvnsOPQS1TRbbI4hDgdeMD6xpctLZB2MqQ
YnPZuHX/20AgqJKCLhSYdG/Y2cY4v4FVBBKKY488GNYANaz4nZz6WllPyoXKRe+kkcKcz7EhYrQK
bjwmYa7T3cSEFR4jU0SZZDJT18mxFnGmWjh0o0Ed7u/vQbvgXr58QhS9BeeW0AionS7tvn5ECPnL
R9qINu71bCT7Q3NWKZwI2UAwRSSeUhVQ+8EvzcQHdKDlUVafIxIjytKvN2hjpxqU+cR05G7s+EBc
sR7RHWvTlkRzrr/fyxllEDyXwWd7NA95ZIhuY2dkO07NIZzWfVU5EgKCzKuFdA5tvxXvldISll29
V45FLRdFsKNYcRUakpUQFzsAaHiO3PVDiHvGAGNQDhXwOwwsPr/+QMUqq+7i4gaVloXdMOyIEzgl
VDtj2cB1JVA9hHYCGdG3yMiWRhtANrYt4Xr0xJUpCohtjELZQlHJOO0Ql1cG08gCdIuxEp2ucw+g
UmMaQCI8Ijankl7l7WrLtZklbD7L9SG6dz2FLZO2J9qxyyP1Hq2hrZYG+TZngNIIvl+pqJXumjCw
PpeYperF+IrhxxEEjq85CZ8gdblPDxQeNeEayhua9nPHd0+M7iBHKiYM8ouSsXOzxN7mefizJADW
xB3uB+CyQSbyYxRGky6waF9D4TKa4POpAmWodWLjNHUZsJT5Qek7TK5t1AC1pZ9Qw6bJ85Z8dY8c
Z6DfP3eFQdR6ZjIWrFuPp10V0V+NBp7bIHHKDpSdjsfDt89bCZbp10405GsufFzcrfhc/rRDssG7
N+PkfaOeQQtNAUMPARNt+vAl/x4070nY5aTOHVoiaZQFX37qFc4ji7Pu3wG291QUAIbecVYttFg7
Kpv2/EAWhyYgtc3sl+Ha6JgNsaFOKz/y3rLDGb4w09IVesEwCgtaU7rD+uy/zn+fp3+XK5Qr1Ads
Csi0zkb4MNfjy/nPMWl0dWT1OuoDMBCNmVHmgPimSdpGmELy9ZVHQUiO4NMH5SRAnGNhzVqw3C7C
R7mDI+utExTWe2hLiRAaFA29CQ4vOxv1DAQJaQ+yYPoUfYROX4qmjmpsW7HTqBVTBTp2YFh+3XpS
2bHm3OU/B2P9zCQX1bWOuYKNBqIREazhyV5t5OFyou9wiW5efuINRuUekxi9+cFv3c5/b94OKHJG
eQHKQ1ZUnuYKPdGLOvP0WtbM64v4KQhYbOdwKpID8QyW46waEtJtMKIDXnZMiafSfSx4qPd7STvJ
oFpwJidj30BEKaARAh0WbsXU4oUiRc7vMqNqnpA7byJ+kbvO0TaPrndGy7MVoUY7IHbmtpzeijiK
+ilLtPrD5M7BWs+PafohRYvZWHbtSsni0dAIDZP7FKqezyDSRWZrpI9NgOOOSpxctle6zFpEb65M
+kerGyoo4ZAgn8Ex243oc9UMrC8cfCiL+MHJqPiQh5Nzfdir7Ga7pCLKadMYVmMysiTLiSIlp2HH
BvIMWbciRapKtuztD5YjX6KFUIeBxwnHWqf1r9rercnlNVPHT2LsZsVM36/IAcBpnkUdBGTd+xpB
XhSLr4jXdB+PxwJbSO6oFNtfABN0G6XPkdn2AjZ8FrdkYL5B/N5q88wZJDn2nrl9N1GnJ6azJLRG
qIMf+QynyKzX9JMPqTkrmb2gG0RG1oLnrHEDxSc2h+VABG4Xaco0DStVAdsOGVq/c+bj/2yKeHzt
0yjEj5cMXhiLopCAzQfACD0vLXigKrwe+MgzF3W8dFpiM4q3HiMcnzw8id/HtztbFNNwVFsKhFNV
8bdUslcl508/7Wo8vZUNTl5zJp1EMsN+hipbBEBkALr+dLY5uszqjS94SoD2eAHN3pcmLHqGgce0
QWke/esICV3Kun7NW06YQKNGWhm9AtbGTKXd7FEFCo3kmpzO7xSTmRkStcQ3Fe37T4Hligmw59k8
fAmCWqfx44FvSHr6UCISmrhpgNDL/BJ3Tn+FX11A6gUASm1KtNNKFNsVR+cmoqjyWhXqJU5HHMQ1
99mhNS1NtkNWu8K0cewBJwUDPRXlXjxnM4YUXQzuCKwFfcRGKPj2F0EXIAeUBAc3kF0P1GBop4Ps
iVxK+/1AU0mNFzxWUSdOxLN5Z3R8Brrq+e5oqrZ1HmNoHMaRm+260657S1kV+YATVsps8dhu49Ci
rGVk3flveKW78IRrCo4ft6gGUwbNtWKsiYVPiP629Qgq7MT4x35hWSf/tGrCmezuppMk57tVpGFX
bKUtoxz87KNqRslgV+YRArIRjmHizFnx8rCSccXgFxCxlxBnHywl66eQXT08MFNaukPTCF865iys
IFmtuvFtGM/vo6K6/fwsJ5ydZJl/d1dK9RFX4ETklMX5a8LeNxxjCLPYLW09VQ5Dt4hZzSwQ8rjw
anWRaIK60KYlyEdVhaGgB7HjKqZyTwNPJby8sxbS4cra+2SzFHJz2JCf+vTLEdgvYXvcFA8r2DNV
hvtf7mFovbBxFXjM7nmpG60yRqRd/xozrINAb5/LNBmJhNcY//QUsDwTkkCPSUDA6Drhv/Zd10yZ
I+pIyMvgRrRJd7NsuB9bYbN6GTGhcJ6BROkIwhwYNwM+5B1BiceOhFQdzqLAcbPNofV6IRGMomYl
L3C3s24dV+vJHSVqekYC89hDQ2CNfiuMtqkvdfpgyyS+O/xkhJB+5r3acvXIa5m+Kb/ycp7b/Ll/
+q56pXlYmDZl22L1PTk7VbV6Jzd81beFfP1aw7xj2m7BcO4GJNlSF/hMSe7Y6OvDomxy7AgXyGmr
CArPURftSkzqD6EjD5tboakNd4GkFC8eHuOKORPvtMjzVZyGR3XalcDJMGmqb1F+lw5qfCPbhCh1
g+8sGfpKnBr01E0KTfFOLM1uvLBRNjtCqCK1qY1CyUXwbF1ga5Fwz/0Xd4lcsiTLlhqvHg1sVb1k
3vzB9LRIAN7DGKiSk1b9f+CwZR/GY+YJfSaBCBUU86SgarhQ+j2zYv7xjzbY77qTj+qMGybmQ++V
au54dWctXwfW3TI4CpTYa1WTpbKMDxRRBa7yHLwvH7yR3dUNiPRypbS8nuTZfozAbbOqt1rgARIz
pr81QRuDAS28XoJyOOB6txNsTXWDWUjv1qsTi3j77jJT1i2UYWw8jnE3MqeI8ZGXsa56GW2xIpjR
zDUmlgCeGQBrVME2H/ZT5GpNIw4kW56b2YVD0s4k9BJSXelrOF8074APzbphRYvArIIhs0pGNXtV
MwuOWzZb5QZCWtRi5hTb7LFa6+X9fwzKdaCWsNnfUWXao9TmDokyhzAxpzbgNdjgHDOpvan6xjf4
S7ZFVysBL8/eLVW+Pte/gBYLBfnumtux/cBwhBO5aCo6pT2t0QBsInLNkYpqrAe1o53Ekhwwinsz
CuDOUpRaIaPVoBvO3irjTY1ZUQgUAuDF5zUdM5VJtEwzWqUIn+50dCuqd/7uM6yhEgpeJ3pgfh1q
lyB2hoZtycHGhTQhEx3Q5TQikU3tbrVRov3ukqjMKtdTsLQuoBtGG9eP7IWAzxMTUmvjBh5DXOMK
eOmzYmyTd7UJygxglLGPox8za7S/4QICMXSdfbWQKqbgdxAJY+fST3OBjvF6A5VWJJ3kafMP+cLc
8NO0IqlHCiqYqpBx4MQphWxC/HmYHAnZXXxliFBdSvh4VOg3e6OAGrJe8nUAXcHnGDpc3o8V+uaq
/iPCcItWDD3IL3LkTRugzefgCkHoPMasCQpBh3eMNH2l6naCBCckpTdNIixkTnVgd3GUnP+EyxPE
/tYh1QGMlh1URd30cCKWbiYonDb0z+nOleV03hqa9mKM/HSk6OYqgrhwtL07Ok9V2zWJyVUUlVps
nGQLkBZSraeAUa3+mFRrpzKDUmi5a7Y65UdTKV4hPSWEa91suNiyR/Jr5zuqN9OQ5C7iciZRPflF
queNRqXKEws4s8c4bYwIOsKq/7Z5j2HijvZMaT+oQqUmNFYYSwKnjcv3Cc5FEEwI3PgCHGSAi3m3
whmaLCuIU+1d8eIGAGwViRbGEcE9N+7+sQ+vEnH+dhFZIwu6NFEeeIZF2rKrQPXn7iD1C2Qmh9C3
AEACWQFKY5m+APz4q4cRrzdyOnoqd/PWNKmwiS2ztL60OZiGDyIp5Fs6oiCNdiu9etckI8z+Bm1F
qvAPVqqoMdiLDsjmFpaDFY6DmLcIjO7WPQfVb7wH7A7i81kXXFSG6LGPLSfmgWSvTy3bkw0RYydl
aKt0MRJ//N03k9xr/xtNMI9vNV2QXl2ZHE2u63Hya7OHgyLfLKiBqxKbD/tQd/Nwb2Hfo7tH/xUQ
T3ZChRd7Fnd/yb3OLv5/4pNxseUWJ08I+W/BO2aPNM5Ugc1HpwLrkOqSkzmy5dmyKFVz/5bHs8Uf
31Mui2RnwMCn8RB4/DOEEJFSLX9aSdXUMYFIilCUXV29cC5JdcB/jJGPurfZA2Jd4EM36WcXOhxt
uJQqRObK5kntmuxwuphRtO7CiMZLmz+LgK0/xCOaz+m6q0/ELvECd9jkqpsHWxQv0eYpYBO9xT0I
QClDcxnnanYRibJhOvctpYXu50OmL/Y86HgJBUFy6EPmEJc+Zvkr5zizpybxmYFz5C/xGUibH1HW
OKNc8+isnJGgS2ah8uSiZJyfxqnqXBjugvHk3ToNw5CuZ45u7N3fAZIuf5gPffx3qyLZWl/vJ+SM
97NNatIpCVA4pMSrRyBK3gpuPoULinBDwWmlWl+pCKyl4nA/57zTGqxwqL0F8Ogd4YHJZbUP/lJr
wu2Gc7ikYTQgYpt31CR/rERthPDZFV/pp2oZKhsc45oEpLpxQZ7Twk506e4xWnUCNaw+SeWdAn+B
XXQ04CQCBaldYix5j4ccF0i1bfQ72/Eny6y38TY5nVjouTneiRfSUMSU7uQYBSVNLWMJkvn5Ht3d
awcSdWKoDOLzaZEtngPCQYlTIBJAPZE+W8JzUpXmHQzbiSpH6nnWC4u/EX1bR4HanWEBwLvg6lty
UpnbVo85d6sC+O4/tME2Cnh/52+gEROl+z6aM7BwXW5CY2/wC9qvklvXi6+QpJikfWT2kvjN0Wsq
93VgaFY9KaW0LhtaTEtUAV+TXgxscrGt9WRQKpaRDCWcNJPa/a7J5Lbz5mYnl3UFU3wMP35sBkxj
d5fYTelAQd/DCeCDNqknSimNMrQ4QIO7J+FO2zpAyMtPNSK8LqH5a8a818BrhB4qUR88uBYL4y3G
1XshraNE5UTW/trYPEkfq3PQqyPXE2/XvAYOcCTYwN3wsr74MtPI3kgSWUBHHk0+JqUJEix6ajfk
ZHamwBXp3RsilCfg1q62TnXRuI7CTQFf8hKKFd3GGyEjTCv4UIn12iMd0gJkF5n5OSWFhEDoUwT4
ON6QvOd8KFvT3PIgHMY44/+wPiB9xWnxIsmFJxQAKjaVu3Gdziz1BfL+ns7g9VDPpj6TzPuhtd5f
Uvzy1YPhyxrrOuBjDF0Zcd5e4wPKc+quvJEUmmq73jUnlxbi/EBI9IcMroEPwNBRAXOv4xhzQ2Q6
KFt4tXlzhhd7iy6LBAl0yC1PpmggE0pcWIvszgTLYPtrY8BWUVaCbh0PQP8CTxAJkhCZyQlqHjff
2856qlkA0e73d3HOfzViLMnMR9qSeFhNhem2gO1RenZXKx7lFTt5JSyoq0x6tZM1sSDtGvE3wErl
q1Ps6nCdTf1N3BCRjN09Tu+xpYDF4uOSwABX9quadkyLQgHsxUX1PouPCUiOQThex3ig8WG8yBqj
6dZzv30UQpSa+t/soHF2JqMPE1jTAIwIA5+BbAlY814Qr46GYW78ov0lLDrulNRZoXKBL5kssF3L
TEB+zZvxo0u/XlpzD04S7iiUZ8AABBrBAPeCNqQev8vnAxO2QFB4fZIu2eOMW7BurUettxzsC/VY
9i8p2R/rw2NCOZMz9GCtQsJ1x8QmUClePkrBEMCjlKvegTg8EMtAkTzFqG+RzU3HYSj6Tpu/L/Kr
8VV7O8Sewy/AE230Qk/NGbbb/1/P77Kd5UwKQPWIsX8qmkza6D2zVG0LlbKN2H3feR08ZEHl1OWD
6ZrkXzF6jlWNrOkMQBx6gGRRsdEWQgGGILYFMrNwk3dnTm/0e6EexuBiHTvCi2rNCYAanBpq93CI
J4PST1qouQ39wquuToXIkxk5p+9F3pT9NyKEbmysjqOIlDjdS23KOS7l4d5Bgh6J2L8uuUGRfmUS
PhdEKs1tbrGNzTsuiu9GMJv6y0o8lBnlkS7hyI50ypt83etBx7EQVDftYjl6x6jw7zrY0d0BxIIg
dJzg3oioeUQF9DoaLfr/+cUau2AZh3s+obl1wNcRuuDROnQTe5oIuRCFiVy82d+PpfGenxfF5oqN
8qbF3QCnE/bOKcUwssfx7Jpn3ezZRa8EngIlZZJ2jsZbnnNtNZhHQlw+29Ci7WIYgQOX3fUm6jFb
cAcUKjj9n69dmWtcDPoHgl2inEIGsWb8fZ9fzbfnmzYmZs1Es7JCtApKV0bDnShjfpkEBvs39CUs
DwzQIVRTWn+ye9xF66gfGKBqqUwQQFD/6tgi/yfquxhYS90LwGkvBBMR3SuLoxkD0rtn/IToawi/
xbElYlJVrk1V3vC2wjwyMXu6L1bzeYdDd15j6v/QD5I9pUr72ruovgaMjI6PLnJYViCP+J1SOlZ9
n0v3cDx3WliQRiF+gEMJTERQcC0W8NcCTRr1OZic71hZr+2ORz8DmrQNU7wWOhLViBj5PyoaOHAF
nohv+kvotqFMh/NqrwdHEg2Hlj/hfh07SclN+LlW4yVszMH5JLGz3WeDmlA9kpRaodH+RWlN+8T7
olId8Wue/b4urexIOZFHCV76LOqNQYE3Xxam0BPhk3fbxxDADk99Qr4F3JWbe6AFGTNvMsanlMrt
KaxbKeFOPDSldmOrbvvAKxXrudL7B7osWmKo/s1p+4uZ+hR+oBqs8nWf7xZocYj1b7MDm72Lt2Tu
NY0eEG1JekqAvakdj4AbYYcnGSH+layvz+pscbTXy/5ojK4MFepIU0GHZlhu3NXR6UMO8kE+DW6z
asMfw/aJMM9/Zfs8nyBclL4lMZttxq6n3yG1rqv73gd9bYq9JXdR7OZPuxqgtMT7xxacn4FMvnUV
QG8ClIgyzmU15bGzQAbXOlLZ43vNDM7SyEb3kysW10974Dxbd4XIpKPZaEbezcZDruLHzLEqvdMW
85zLjpi/Qa4kNXL2HHmv5YBJxP3bMbMkhj0/PWxQMn4S70WNMo/Gx+hQQc85HJb9nEAxF3iEBsKn
7KmR+USJ6rNm46EOS+K4JK7EXkMPjZEkJVwQTPE3ADE5ouwPZyZ8JS1xJoYLj8I2+M2Pia77aG2U
PLVBSdgzKF92m9znQoi+4KVG7N1AOgrgFBSWQIR3ZAhModEsdSB4lBAb2f8sRkjHpDl2JokodP/O
WBLrPG359cgHFmHZrQvAF5sRP9zD6ZtpkXQm0rFFwNGn6mzgG4NW0eW2MeTnkhhRSQ+eZkGsCJ97
r81ng3dcZK+YPexn4WERSbyXdMP2Llh9gJqV2nsX41vuR+uZWr2GXTw68UJ7TQ3JyKfW1JAGKxoH
rvaPMJHOTuiZPF/rGiR2Bcb1Xq9Qm4Y0N+S+VcIzMVWADVKwTyBOQYcG0WGDU/sOth+8uisrwfrE
SFHbEj0Bv+w7gCnQ/ZDUlj75gbToaHUAwyzvoILdEHZ7C0DajY0QThmxc4Mu7iSL7vE8uqp1VL+G
850q+8scBRx6pTQJ7QyjynTGCyWZpwoT2Dbl3Srl9NVwQpJgL5OSQXhPN4WhUjmuGMzoT4RoAWz2
FiDa+5JNQstyEuqPN5ZdV0pllXjZsuCpjws4ErOzOwSuy7h/hqRrm1bxW+2CPe1GvJWXWJNgjwq4
xFjtcIdWq0AmreX7eX7yhT+TdUvUzGyRth8wLpu+Xnf7bgkaFGulThy5nrSouaQbuXwipkR9PBr6
GJ8UGpb7zFuC0Ua/VrzaSi47PfI96VV/e4hJ4fg+FzkY2szzutPabtfn8S97c2lxyxpdPpJQ7vQU
lX1jyi72C4yB2xSIhywqKeQvNK21gDFSqkP0aRRDe3vbH6vX+HIfuvtEphGsGjY+CsGwqD+4NFNC
NVJLN9qX2g551visxwTH8hMZw3wm/YYsFXzjqpBAS/4Eobm4oxqebyrkbIGmL9VSBvJRpvop3+iw
4tAQZ43XPja7hemRozbXXxJHNqmPgfXUefye86TwxwL99ppe7eCVO6+JiGbyTXgzIVH0lmMmTgKM
FqAWiodnZn0xt/kCC0VDsA0u3iwpu346TYFSuUI2oFDXBh/Rp+PMIBItbqEJ+i2EBboVA/+qaMd8
mWA7EZKjKoClDgCdcyCZl4iaRiI3RSaT8d1ce0vXorqzCFcyMIdIz1ZxBySNl0n0HL6Yj3Ujh8UI
m437Anf+Mb1NOkfVbwIp2+LOddHGFmcjUqpPMSdmPjc9uV029B69hUQRhbxcxGHpOL2wihxxtEUg
tusK+odqKys1n8ooCIStd1zn5tlOV4cMsq782L/9vrLQ2n2Zz8GGK3/jxoxYtBRc/Xjo5UsxYlOW
qlPE7rjflP/ZirBmPba0THrEkpEsFxRzeZVF9B3QgpFDKCeJCp4Ch9Dyp6VwAT9VC+bYFLjTKgwg
OWlTbg82BqwIybas3ugLpbuyEWs2+ue3B3fA5RFoPAlNjvaYXo+k/m0QktYONZ7bTf3fLt0DmmAG
G8wz+SeokrhF6CQxXL9IEF51ZSUoJy0zv7coonZ0U6khPJICAjlhlq/QeCRya65bOxOc3hnAGB6m
e/7xpHTAtVuOD0AXiI+g4Ss7unW+fsFRFbFeUp04uhae1//A9t1JPwSZlg8XczmOep0Bu4jdM77x
YLHyw4+ZTxh5dCkFxyxqdQJrKcHgMghcd4dXTuuUoHbvmx4yD8U76xJMaJvECq5ri2Ra/LcY+sZj
QOCcIAixDkUqOct1UDCwsj2GhM9EG/SBiasqZK8ZSvpyna//88iji0WK44OIgxgC+g3AEYZ3trbl
ICCQ02PRcXEFkOw6wdzmhMKRxOPntB9dsnSdrrI7U+NmvOJGYcahfCcmzvO6OKftGaL6cxK+9Pjt
oBb6h2qeaDa8yoIuK/zXI8JpV0Fj1U4UJMCVBVYLyIC+LmXSj9E5iuvHrb3puWFhatKFuxHKhjP6
kvSzg3f20BaA7oQlGhgYFtpG5i1Qg4mFFKNSbNeLQ0rF6R2O4KpoVn/UKl71xrbZMZW81Hg8Z9iy
DQlCyNHRwbjoQKfjkbfid3wrDxEH1Ig27X6zoPmPk9IK+wRLCkx+xsUn6tBNIIm0OmHYIVnHgtZX
G833eoyr+Jzpr4uSYjlIKivrumQLKvk9EnSFOZdLsdf1RqnHSzZ0IHl6Shf1UcTxLAhRSppLVcZH
tYWJFwRp0DlNK6EIUVme203zjX7nOqElW/9vn4GmmitNFUaa3K3n/rqIfnC9y9ayop8ALn1YjL+9
I5xdSX3C8jyF28Mtzxgg10EBCCy1lXKVKB0sto4rRylpbcQcGEgd/ep0G38rJMIeTk+ru7dTVlbC
R+XMkV9WAkfSMpjx82+vbmszcspgVsr1TUoAgeiY7ghAQ1gFVI4f95v2WeYlLl0Kp9wMHg7hguQ2
FWooFb/KSzsKLJa54PxoA4ahwn3Xtrfe2UpABFZ0a6REbrQPg0AY+6Dc8KDcMlKZIQ2rtOabuceu
5tEGZsWMd27UkhfU/alhix3sKukFdHm+DkWo6DGXEB6K9svC9phspEbdSfC/IRqkrANKMxZ7PxSb
CA11GL1GGlJF3+hCzPIfGO0xE9B6CtBb8zRVRDmwZNVG2B44N2GkpThZvkYx73g+u7EEVJdA7xW5
Tf4RFG9m+aeQ6wy295Hbn86meQHZdszNM6Fr1aEuTW9VH7LWWEUODgs/Z4psU5lrSON6YsQ6Ivbg
4jEkHYbET0HkUi/RzJculE3WbQYygk6BBExbTh7HEXLiy9iAgaImBtcLNduHLlgRWS/GSm6fu97g
2t9Htx7gb+2LwBG/5BPDafxTe35APB04jAbkP6r4JYYf6ySu4jGF77WxSNG0J2WI5lfGqwyDzvpB
aKH5AcMa8Po/ZKyyoyI/8DPvOHSDD7M99xTSWuzEBZ+26awz2fMJzmGOhDQrEO+waWaGUre8NILv
dCCpNC9tMKQrmKYuiVyzYYEEshpffKhZrPRNx/LVYa04iHvlAfKc39fiE+xegp0UY7/aEW9ZH+HY
NCvaa/0Rsd3gS46Qox0KMSzF8pnQUw+7mJHVOlgAXBWKZBXsYf3HAUVN0jRLokBlC0pbK6drFzzD
BVzfhCgMYrOkovcKWaj0+UKV2JE/TBNQfvdpU/bZMQ2FN0lo3ykHq+oLfyp0UdjjdkP6fL/e0kSQ
GKJGm3jxpKObQtA+MCgaHrgGtSVXlnJhmqv7z4By+Dh2ZF502HFdFmu9X//5hSbILjqZnfemtZpV
jQC6gfAs1jwqTpoeAvXo14CXOQeio3vjGwuTuHGXbS07oNiSqUkWXcutoTlaovTZQfmMn3zYBN6t
aySYLcOuv8nGL5XHYRpDzWsFgW4kcVPSYp0G9UDJqOlMUM2gScVotiBXKIyJG92WFp3o5E+yh2BQ
pQBe0CyK1m96T/heTys4wUJf6ZN2dVhn1efs9Uxx3xChuPHikErPbu7Xt15w/ozoMw6/qH8uGTgY
zBRMcjLMBxk2ClHTOp7IBmk5Px5OmjHJzG/9DHMS7RDedeH+AXqCpCEKIC4FbLLq1dj301g3WwgB
QnSJenDig2DaW7ZJfOcK5aR1L7NYdLNN5TtXC+7O0G3Eh03ijCnZf2Gke+bwjxPz5owwpgA19xMw
48mvyrJ80/8I9XCv5XrDZ1csnqzJwGoxUEQzGPkyIUwDGoVgF8saE9O37MYkLDLEmTlXsddUTzxm
kXvrDB9aSgIW14k1JQqYOb3sV5phfJp6fza84vMvIts3+yUtHjdSHMPOkcwAMIjptOOtGlV1TgvV
yGixFq8xVi5yvJhjz5kP535dveojiZZ9pQ/iIcy4QP5U5VazRtcXO+6tvf0DcndBcfpIiQXqomt0
XtSzc2xBKoE/t3qoi/Oep7UqMgRFsJxDGRPZobZZS6i5YlaFWfAXC8t+xReWujP1FAHuvpUtgV8d
K3LCpCaOtI6EWnxlk1KVresXlBD3JkyfysrcM8UVMFq7tOJ0qLQmGYr9jdT2E+U7QW08GQml1IhS
LTjU2hpnhwzsbC+e8Fa1xh9pJUrNsNXkWCORXemiEgllB60l51MX5XLh4ngur/ZVHaHXdN1LfHXj
RLoO6/GloyAQl3vKKld3IDsLqsx4MS3PnofM9YgX/O7OcXJIwolnOwuLYFgdu47JcB/UkhSQK5Cl
970D52chyIkooYuiluofF7E4s6lXpswCZ6tJ/Jlma971jVVBuMCKtchZDbnRxmFdQxR0Cn/SeIOS
jZkWbVXAYk5qzfBXFoA/VRhes42X2gX0x6yxOu/euYM/9FdtAiUReo8+c06qRJw/8hM8oMy1aZrP
/MhJO0Og2kS46SxU7rFwrzt79d72rvqW2Dru6pIZacKrKOjCfh7rZ/qh02WI+VMoYDGENzQBMH+S
rwBu0aK1SGBfvCYdZF04yWX8MhTYKgz2ez05SPxeknpL9qTBdgURUqlAxtKsuWZXlo8k5/3/6j6K
Z4g7wGfkmXsvKIbASlISn1TzCxTnzOXEaxaozSDn1O9Jdd8JeUJCL5brXi2nVx8TJypI3eGEInvN
cBHmwHD3/dt15IRSi1K5J60IrVvi8hcg6DXnMWvnlmEyAZwUqQWXzMtNlYUQ0b9F05vSGa+yYkig
56gu8Ym9embEBK6TdVt0/7jv6c1KPYob/lN85KDOQyEqgtZ0OQB4kYTZHFHhCu+h6tOGEpDVGkZN
TDkYklH2vQlUkLZ3h4oLzOJnOo4J8tsxf+bv8z2N0gLd1nYIOlaGrM1pcylubmZ13f7v4aov5L8/
IQfxtI+gAE4FaljZAnRlj8DYmzFzcDlVpZulDtGVfNEI8p58CcPx0i0x7fMvM4oy7IoAU4yk9/gJ
ybMg5EdTJ16dcgL61Aobf4dlJNuXdTZGLQtAiF0yNEFAiP5wr6T2lSiVqXoyNwa7PiUKZKKcHNVH
dCbMihQO57g4sNfPb7uVwNGY3bNKS38BAw0LKkYbr+mnSbQA3MBiCJOoGze4eb45UM/IM5xsKPAA
NnSHE7/PAtlVNav5VY2l+CTufU6wRcHZpQgY9P+9/ZjOplZGz73CzqftTxdoeA8miNWKxxn3Ul+W
e7VISZny/BKilLQ9UcDw2svOwfCHa7j/kFuL+X/QnZzVYwuU49Ko5FTZmmaI3WWwSVDcpM6l8ZNb
zlwEeiAhGTM4embWocInN1xt62R89a/v11uP88LsVrjvGaoMSNrEq24XY4+f2TQwIrFLBRVTxc/7
ENconr3tLu7RQNEbCpQ/31w+Urb2Na7rk2cu+W5CArfDxk8M7WKSlyXvM44vAZjSCtLdeaoRDFv+
CO3XCA8Qhnwmqpqlbm6QUy84DdM1+7mXrgdamGI2FLbUgvzBPf9TCls9ScxJSj120wLvy9OhLSGx
LbKEb9MYPsPHEWo+0Qxz1Q2lVvwyIhBEUvi7uqpDASx6qNnZ41p8WPt8OsUfkg4y9qCfSQbA9KJV
4Kkrgo9d2Oc5FVakFH42nYXFynF1EggE6CusaUQc4ybNOhRN5wrwbGFdcrGz0jZkLMaWBsZM0tkA
dMkeklZQ5qpJ7BUsXo1YiYlO4gMUYl/WUzil/KzizUlyWEM+T06MHc6HrCbweObdMevLM7RaBLMD
PwXXubFzUtnWh+qFwYgtUq7yhnEBKa1Ie/EaERJPJjubc734EUkkhJygznnMbhzXXgkd3q75BoVm
5Z2GHnebcpW/QhAOj9WIZyFkjNXi2U38nxH8jl/xZE8vOx67opTmQl3WVon9JWMFgn9iLABMdAiA
ej/BLGjmqXpvdVjNOH0IGcndqZmjnFP1AuFNj5+49BNyb3OQpW7aupMXSc0PFgeQaWb0pdxhfses
k5WYTQxvIGK6RFnnM+FfBowKZrUTXqQ1SxW5Fdo2a3h+tHdxc7sdS0OspvMTfRADxGwcqiOCO5b4
eQKsoJjKZwf9fc3X7MdQ5K9A+rN7qkODZvrvwG8PRR6/o2tD8U3AuafYtlg3luoelxv2sDkXAuQ0
r9Y92woii8HYyDXpMM4Z2r9kwlEJYmY4v3/JY6lJhSIC1i6lxiR602NgamRszgqBQc7vXJQ0fE1i
7QTLNMkFoNj78WhIyRfEnBkP8h2lga/EhQXevslHNEd3JvM781JRfBCZdLIZ1UVkgWo1pbmF9OGN
f5zm5YzYZxnDf6RwO/0WUbe2WyvaONLzMgd/FabPQL34WFEPkDJ8gytSKvWSwfasHyrZreCbQMlc
l8PiXWWyt9b5iD+cL9tbz/OliSyMguOLbW9wJl1v0PZ13ycumJqZadFYzW56c64lb8+0E76jBrCH
j+TZzlxq3fZHwH++mMCOHw5e+ghmNUZlGLGNDfhjVLDqzhTTj8d1EhujMyUyPoR1fWi7xp3zy+Y6
0/ddZGeWNOmDd1R34jsdmrjOvG7mMcaXW1p+nI5/xbSRjhXU2X1S0Yfjr9Pi9T2VWme0/EtcWg+s
o9bej5FYljLBZ91LZI9SWAA3TCdd1RU5WeqlgaCsRelY+B6OinSyyltmrUURZIMJ+yzUYBML8OGj
ozPDS6LNoc0DDbdwChpkrUmsCflSpEd9vnyTD2KU7fxN1V1+of6tp8yGkRe/WH4uN+jBNotOqc5G
l53nQAhmS9lhe49Fc+J0Ltt/1y48ntbaUC8aAxroBHCr1qT10V71XPH2GDuRm156xmPWoTdfRcVa
nG4XtfZnzx63/+dEUcPFNOToCgsz8Ll3gT80/+IXaGvK60i/sjlpgPhGJEqJegf2DjAjReMYUPvu
BWgZaDlKWZ3vMcz/wml/brDP1vSZMhjnDC2SpmAf5DyVNvW8SF1XLgLX/7EI4jjmOHonW3Nb9wk9
PhN3LlgM79NLibeIbPekTzA/oe/2pxXqQDLX7QxtgFIkUbSxnyso9vsr1j6IqfbmAiq1efJeHQXF
UawN+KkionoqbbDKGiYU1Ug4ZsDlyxNJ3Mk43pGYp3diOhWIsIQqtRI9jT7pMz+TJdKHYmKJrkpE
r9n7vohQu+G38QKUaSl5a7nGM/TEEF73ZbPFXz5Wiih6VmguAMLNNUP6vZ0ZDZ3hZfnSMzx4ZRdk
5gQB//5m3SmI+OEnOpeewsP973w4MhpcqahYFMEeLQFTUXEtzjRoNRRI40vGdynFB0HrReXWGP1u
d+ywgRZJCNdEcoyFKqocAb8f58Xz3I4GoanQHwM+bJ85Jc9ztEUaXkfdfzhHdtykBMdiGghQs5DM
iuqvTh5FgZRpJ7OfoCD/XA/xy57/X2aI75Svbq+U2YdUi9hSwmtLX9TWnzDUjYacj3DDrHsqMq8v
ObDSyIBvRDdTbEBdQ1Vnmp3z5ys0gAPM3pa/x+dmwepjp599yCW0t0zvHGkGoMCviFsjc7wOHtve
ZDaTm5Qbx5w6KlVV+EE8/7tPt5XHxgCiwWqlghS03biXgcjDERGae/fZjJXgld0JREIjYY8nvXt+
dRra6+eSgB9Ltmh3a8zQg7Cqrx6tWZcE9BUWyhdmh4+XW32yiPUMcWD4VElaJJK78XN3RQ8CtlGy
RSTaeio/G/lH4jRuiyyyxTyotFvpcTmDm6nWrrd/jYJHejC94fUMtdnCBNJTFoUYDWyhUkpSiRwl
tp/bnB/VTsVl7vu909MoaeV5Jhh+h+NF2ncxwDG7kIoskmsLefdac07WDNsBTl2raja4k63o+O20
XNc/CmUxAZD2wLicg8bAH3TeIgjHu8bXlDiplOHI8Ovm9rGqnIBB3jt6671+Xd7ZGBy4XZUnmAAK
2lWa/M4A50fKFe2WEGwvyshv2g3SULjDica/V/prJJntn1aFaYEbveJZDSKk2F8EnWfmSV7Z8WI0
nsy8Mmy00v3z7ObAeWpN4pP7cLvlLRL0DjbjU7svdqxPcs+EsB4o/OYmL4BUpBbS3F+urxFIPQHp
AtS/wdoPSmkQ36LZN24/N+VaPPiRdtR7PUiLr87bT4QN7IxSh9+pGxcVTf2rWR/bg1QB/6h9WruY
O61EiHigxFnY3dC6T7zcSlzLsC+1XDwQBi6t7fXWj16tgZqH4XPd277yWml5mLjqr8+E9jiJd0+p
l+Bh1zsyHo8i4jzGn7wCV8nCSiIsT+BEd7pYj0B2tuXivEymZueyLeWUDKPje2OdRNJHnpV9P3lA
Jij7+IHY5MAOV8VVDMbiT2OPJWTcfDzDwxSTk4qbDvWnJMcKsJ4+EypaXwJmfkyPRgGZoGPnqTV+
dHzLQ+H3dvD6eD8BcauNBw/BIiQUZ/+pEGTREAbG8DbR0m5G3+FeGfuZTz4TS80J+gnLHUiXTJNl
ZzVx6HPm3JFPTLJiTdX04sH4pl4Ges5BilRyG2iB7L0jvGc5uL4bzzQgOyZDAFlZZ9FOgFzOdNz1
8LDVd1h/r3ZThea6PAbdm5mVUkdzm5SoSOddinN0Sri27t/L/wu1iwaXjiaK/RI2IzNmZviRfDi0
j4O4Jf/coDLfpqSM/cALwJegA3CFv3Chox3zsgxVxx72QuDlTM9uMqrfXOFYXjhKeiUWFjsOGSw0
wEmINxjhdyHFc2SI1Q+FgtIzcNxjVq74kb04kqoGbkyEFCQpABrsl7onC9EqDIWlirgNqbDv/pD8
zR1vY7QOwjBCl3YxAPZpXJ/pCti5earC9M3jq5bDri+sd3XCOzAkGka1J6Tr48zN0NU6i1l2dZ8R
J+1EsFPJvejBumcLT/BteqqWRb4eZ30r/sy8gJhYKvEoKiQFqyi6zUIwIXoG2g6d3NM52xHoMzOT
LEA//+iAlyPOE/5XcwcH0JhicwMsfybEO8QovYWfZGTaxDpZXh/8EaJcmsnEQVe1MyMj3ilzYtK3
rPM7VfQsmaef5fSFQYBdVQoNs5Da1Q8hEvdZrz2n8i+dWTNx2/3Avogk/qnaPzNzcerpvAONh6p2
EXaKIUKwAKkD3QzkkfUINiyPGd6npKc0NVuWn/zY5expEiE66ml17UGnPsZUqwu8z0d9b4fwQYZD
UOexrm+8Ze5t4RXQQh6OctlHy5LL8/UdylEESLJsKpz8ERd4SLlYTDC0BoWgMvNCwkkY+WhDjnu9
j7vzt/PeezSRHOYFosLoj+6YRaegqbros2lUZ4rZqc3ZdQa6FNREdDKfLNaR5sAMDOJBDmdsehm6
KTt1kCFN0MpMkavfP7U6tIujoVYZtAT4TSDdeeNS7cPBeDM3e6zLmJs1LGjQkctIsdNx2735dyN2
ncV4zmX/fSlvmsWflMrouae1XuJJ4folCAjY+7f6i0uc4F7t5az5258w7p02UQn5dq5ZSONTrgum
ET4mvf3NfCuUCv8WKgD6Z/cANiPHOhyEVxXlfO/08+k2y0wHINTH0xwtByf2DKFg2qsCslRAjSQZ
hzJwTl8t/TI+7cJ1Qnr78v+8UD2M30j2YTkmch+JkajmDrOgrISO7z5P+JSzacOmYRIXUJRo1LsE
A9U9HheqUFVC0duOp7o/ydTOvu8+50QUp2c5wqIpLjnT5+TkgWU4Z3l98mUJPK6lyabNienl/CiO
PSzUvJmPWHjefGym5u1mgVDZtk1guwsFX/RQYuFlnmXFzZb3EUbJsB0buFgjbSOP/R8XA812/GS9
MbiTnxijgSyYPIl4u4HwvH5dv8pamLFt0fpDgiZJ63dmOVW9x7vcG41g1OawHKGUEytTghqShyHY
N61Po1Yx5VteSiusxvLXMrUaXPqZs/EEHIVbPItI4lpwrf4pdGONWnxPXioRX6F4GACPErwYjQ/k
YpbbnTOB+SljT4sxA0M3Z5zIR8ajMl7EANsAxv6Z7tDS2Agh27hmEytLUwv+BF4vwYOexnsg7cJ2
iBJHf61Mnw6MVFkm9kAQWVLq5swWDw8TTYaTz6RgOMLM6hAOSf+6UsrVAs2QcuG/eT0TLzWQkvR0
XxPuYR0IQQS34Z8e1bEy4mw8+xfxg2SXIDSGQya3BZcwslgmgxsE5rnipOtPVPo752b42nijFuuJ
HbTA0oFGPNzb2tfG5PhZW+2HK6NKAnYOWw12SgV8xlb8ZvMjMgF2YH1zuslls6kkuL42EN6rm36g
468UVr3VOD8KMXXJ5JFNu1+lpnSXOqGITGOxlJDhyW7uYofUFV7VCGFM+twu+uWkUN6VnfgkcUkz
J8Zo42QDggLzY4qYF2tZDEwa5lz32Lul+XDFTNva2RVVMnjnDOU0PCyB6l212V0SLDpbsmHhT/Zs
pJyYM/oWLBiMyozq7RcHTUO3FIV4/FMUN+7mouHBtUgVOTqlneHVlNatT/ubJGvZRu/hzuEZeZzV
eILtCNn8bh9nb7LwbusC4ro7txj7Mt0hpEMsoivs2yrNzpEnTBk3M75pO6/0BeADrChP8f4Hiqz3
n/FbYN5zKGxHxkjF1MisxZo4NRK6/a9tgLGh8+x3gsW9a1i1DhD7jcKji0amGMPKVgQeMaa5fhBf
vKd1npd9VqlCbr/mvdVekHyE9MrSUarOQtyrXrGofjKkHCNN4oJCM8BuarfaX3JVkq+dU94SWCN9
EHg7Qw+Ul2mby4JVgkoIv9ElS+7x5lK1UjfA5HT9I+YdNQ56At89wGcbN6/zwAT40RYa1jQyqFbN
tksgbMTxD6vqKQi5paQVqfOCtiJaWZqoyhJGEaRFlRol9Z8qf356DqSjd5tmNauJ0qzmdcIoE9Wi
GupTm7or9UUGrTo5omfbJpZo8+MTAAb9iHdLO6LFRASmiHBSAQgBzsiT0uhCXFX+PNsnHR27Jt8Z
/QvyDkulVvOiDDrbsCMBO3Lz6FR17sdvRYukugPS5mdwJ0ftXfr4ETRkfpSX5poEX3YaM1mYi0zZ
Vl96CTud6GYH+tVRm1+/Ss1pyKmtTl5x/8eBsyX7Rpr0aPdyWc8up/Z3V32vTpY4A8v1zs65ikhz
pb9zN323vQzyLtJRq/CRx/z8U2GLkhnfB7NuMS0w0x8sxupHZJUL6JCbJMryVmF3EROs+QQdIH8D
ZVEUGFL/H20QV6hcCv29PTKihIRNrk/Pa1q3HzAcxw1yxirTEc465wkoZhshAli+u3w9NaFxP4dn
jmxTybcCiWxAoaccik/RijXTenJFcYeSjJeAluzlHiYisfuBcpbR/nqkEz9eDOebQnJQAkJ5Uzys
Sae26U4xnuywzp+A98MuCbxG03UiGJc32ymia9CP7gOKn+eC7FsAL/wZdJjEB9Q5Nses+/2td2DN
qTvUpdzjfDX0hrQaHn3aqSFfGyKl+iYNVsIJ6xlP8/nB2B8YY+thYQIDQ3vn60OmcRJcy4ykHjdg
Upt2+5lcSyJBhktgE92vK+ige9QRiKKipfOYMl7Z8on2PV4oA+bp0zxyfcfRUQbyya/2s84k+xIp
+S3eAwcsdZg7Ga7DzIoHep5Ecd+jamqlwtB65G3/1PWnOWgpcYSV4fmjtePwUbckScyVCtP3sgjb
CSLYyTfqNpIuu7DQurCxybbg32GNVJffvAXlSjh5LcyZqcC+LyJ7BZJp1mosqMfVldjQZOn+lMKR
Qg6j9EYxNkGmGBMbpLDlE7cG4UvwG5gq3pE0StxFuKBpkyQRre7ws/F5mNnpeZGHbbDoHAUan1cD
DTzwFT3ULIGhOSSswlKXzb+xQbZhaM8HWgSiook9jkCVPzBwH7rISr+hpy97dA+5NSIi5McKRzmp
sp17IWSXJOnpb8WP7YkvHpGoEr9xhsGq8zZroPHWVhKYZgtQJTpwY/F7Qrnk512GRSkDsOTifqqp
5wTumSU4D57rGjCbauwwJq22uQHOwPrK6Xk9S9oJs4Uj/miA1OIH+04fpYOQb4GPxDyc0us+8cPV
DKxfYKumvZ1vjEzDc+e2MjzIMaHRhpHoVliIuZWc4F0vVoNTrFbgnh/VX3JwF9utfM3LD3jPrJaH
dBF2GJZndpe63P5d2FtCu9AHjVi/twNCUzSN30/bL9/DmcDd2Jy+9lA4xDNQMoEaVKGuRPDaMoJm
wC7vDTnC0FrkK/fA3eQYfe52fOuZrX49JWEqKoeBHWFy8PPZTDTpkGehNsXtbYeA44o8imTxqTbY
r9jXMokaTJrDNkYXddbbgh4XKEHGzBv1VNxChJK6RtuKZiTsNWwK3Vil3KRqR0O3j78kYVx9NtSz
khGvscvuHhWJN4DS0DhHQuRIINioci83vsJas3LIpMHs/GTV6y88Bwn+8ITayX3vT9d+yllZ4l16
ixBj0Psviy+vdFAnVpRzvM6Qi8NAAN8xXocg27C2IKLTY1I8+BSlOagRTfqt8N2dlxy7VGdaGGFC
CXavPzHJUMKykZE46r02raY0/Cz3imaZLIt+Xvrjp8vk0PRUSOwzJ2j4IhZrc1ERdfZ1eB83Lqo8
p4tK+JjTeiqIAoJF8nFPpPBg6hm2XdqPl6eHigry8slnbyWkgy8kDIhcfcDTyJitb+AnwpFWRwtt
EwCtpCiVeHMdHrxivLw+gbxXf43SJj8+gzwwtSLVPemnWbb+u/WoNNLy0iXjnEkaWJj9YR2Oubvz
sNQUe5RVgyBkUoaZ46zzzQaSyZXQAmnQ+WMrqU0/FWV8oXP0AfYtQ048WB+LzGH0xIl0tQQWxsHh
LYqGkEGv2Fc6R5QJGt+9xnP/R0hMy8iTQYYbhnLvN71nkCjItYEhA/ULOS9+z6TxTa5D78TZ6mJO
sBd8aLTIDWaFifEYMmgm90M7MFGKJD61rt89/+A5zDQVTfRBI0bCi+XwSmBvnWeabrLNIM+7XXDO
7hLnlNGpdhZo+j+HGU5Ge9Zshtg2K3r3pACoQ9gTeZR/nNbrhXjjoJqLOz/MhnTnJn2uQJwUKlCa
lPsOi5hfT8AngsyWwdUPnWlS/23X+ez+72R+H8dVbzchvekSV3h0asUIf+p77T0bXOfx6FZjfiJz
MTHscXdDYewRbwantAIfZTTzNjKNRjZO0+ieFXbDNNvve2XfjbvAnHaLGYWRpvExgKVGrw1YomNj
zkFTDyNCc7/odUGxXzitj+KqOSCts8Ef5LN8MQehne0VPSTpbjjhp0cpeObatvdlvRYag58+jgDK
/jij2sY5Wiw7QTNqBzYV0f9Z7jRdGY/wdgG7FpAAuO9lxnj0Vj2nzt5fP95mYIld/aOq2W9wrFuV
frs5b/TpN9nhVV61MDM2cp2W23L+Wn7HJgCo3ZI/bSVM158EtPTVAEuFWhSFb/4Ku3QWcPQHguTY
NscA2R1LqwOHp/8vNNirz5Zvfz527D1Y5Mf4fewCmTC4v+Xk6XGT7rqnFay1y4ZEl3k//0kBnPbh
cjz+v5ugtOdjdlGt3ejMZQ8w7WVi0PxUEIvqX1nxR4/U8HAhKUs/GeAhLeyAQuQYFJzOL3lO6F7J
aqhjPSqpWstnp/k11GrWO/JF6QRjVjOn79CNtz4nX6XIEMjQ+YXd9fLsBFONMEarZxEE0ASih+36
JJ23B78ORpx0AoUim6Y0iZ1MYBg1hJv4ATvwguDQh+tdwFy6/Ll9aJU2EUzgmoIvNBSHyKtUL2Ga
kfDOjVRHED70gxXm+GMFHFPX68jVOLcZJQXRUYYMu28KMsu8gCvqIaRdUMW07VlbzhAYvo7U4Xfj
csrgPQlNhLbn7SkdDhGkKI4XnPBNJIyhT0dvBN4bMDIYqc81XZ3ZThlgVGvC4FRRBZZeKXwikyhl
rmMIr3DwpzD4tPC58SGL4JpH2G1bMIZydd4km7NTez/rJcfv9noEnWTcu2fqQDQebf+JJF4tfZb/
97d9idzvKUssKZJmh8v0m9EBTpRiLvGYz06Dapsi7xRvfY4AYWzruJIV6KPnPwVqw4tnICXpFTqg
m54ABEsrmjk6pkcPEWpWtm6CFkjlArJDfC/RNalEYmkgyIQ6jglpml7v4gyqiATUDOFxTxiaotUp
t0vHrCTGC6OJgAZRjOEasXNKDIZNwP5+0N34HilM4u234LyJbFElWVzvs52m9s6dPzg/xnm9X15e
KJoxuMdoqI3VuoL7wNdNmpc2/lqxgcI56ZuaWyFxDkr64agS8rTepYMYYcZU/Ob01AUbEQVuxSYg
KoH6pKbxyxziJ2gbQwOx5DQPAlozYiciYIRQ+M/DIIrEhRpMAbY5JAV41a7MkXPnpqxwr9l/kn2b
ivJyIXHPa4d+5Fzcf4wXtqjPxTBRI+2ouDy4Gy2S20kus5HbzM6NXTbX0i349X+hg+TNT+++Zwa0
hRpYT4Nu2uWnCNdAVuDK5KdxBojO9469XaJYjQS4aUO6A4r9ft/0sxWGlT9J8PNM7XiZyc3iOhg/
Nf8IxISrPMVcHobhafRaAWGE/WkTcMluNLN0KbRTK19Fq1MOPr1sm0xLbmjt60HVcNyK2Lem6G+c
H7LQEwN3/OF8FiGcOpo4rjzTs2vMXKgqhUMvYFpVOLh13RXu1cLubpsfI6mMFjZSL80VRzl2Tp/J
A+q96CwfbGDCPVLuc9+QjeFUnPluVPaeSZUURKsBCk76TVYdJzqNUPV41nL2vV+WeFIPvJBo1OMg
ugRVcUJWWrlxG4FP+EsDJQn5gVqeGVAKN1bE4EqFO9R/qYJN4bbMdvYoDSaVC0MNAYJSaIrx61u9
AV5Y60ACHpZ3O0dahFk3bbQyjditNkMZrCHHp73Zv/aWW6lKOdejYW85oA6Spn3HMEWVwx2xtYFV
E5AzJoiC4zs8tsig4+H6coH38xhCL0yNjL4tT+WGghI7iQXlVQfsaLiU3Y5+Ja1QUcEvS3MrOOod
qb/kyKuEANiEcTmbst8HSR8wL92bJ2yqUGiqrD3znEWgO+BKDRTreWocMdbiYMYvjYUok3tHmd4L
DpzcOvhKqWAoId9EW8gf32AhbQoWg8t94TlwwHXu87reQZ+OMKcAiKmtP4EqxHeNrwxrJyRKBWBi
YyuMupxeFDgP5uCJdYALbQcMXZk1nvFH4rsf758iB1w/9aIifqR1or6a9lnmmQTybYPq2M7IAM48
MAFbSzCTfsFX7aT0fEW9oiYeDPbRrQbpXJu1FsV2oasIN/kynElImaTiFyckrl83Iu8Get49/USN
gQftUWyfs0Rik2oEpmb2o1zcek+euU+RXipkpzmRDI4cexmLf99QFAYcaYNgZEF7N8kf5Wq/Fdkx
8Kty8dgZjsLwlOi9f5yfzURhMuHfnENSOX8q1bNiO0I5TzFQSqpi4YS83x/60YuN+qKsRTofhOUM
+KMGUqaIJyjLmO8kxGvInwAwULQp0PpR7UiHe921QLw/wLvwxHZSxxUivgwMoo+mjxQE99cYM6Da
Q6ZW+ioTVEszA27dzXq+nzqnpPcyt+YH9f2DRmWKWWeP7ukmLDCmhRAx5tVII7VdE5Y65afloNxm
giil1gNyFJ2WRQr4iX405CVDShdVFVMjJ2lnlQWdiNM3eAlKCEIHg+ZoVsxecr9jnpBy9sBkyPWD
oogujwh0e1WV2C4j/Baef0B4XRmAFk+iAvuLVJIFoRS61qJSYy6kw8RBmi/ks1PQCxF8Obbz4rst
WE7uPc5ce092RYcFWFc+vlWcxOLUgjMNVNU8ZVjR6q7X87WLufa4X0aRrCPEV7RKTKVMYa54w/5u
5dPz2YLUg49/XqwOfx8nfBISNyqm9w14yoWqGbaztsAxmBJnIh4x8w+Lr8b60W8o8LUmr10bRDUD
BnPD9SdUA4s2MoUfTDfWN9jwZ0v2yA4VRHiLTWgB7K9lZf4Hi/OtLsm1IbFUN9AfcX9+D0aZt0x0
lhf6IBy/raq7AnFCxcc3tRoW9uB145NE8542dgwjFMr1sJzbq8b9pAH58q55B7pBqfwh/KqRe4P+
DcoTnktcjDhKV5gijIz2UC7Gz5cqTwgiiKMxZd23gYOeUx9PsLANwo43YVeqIRmxg7rVzeSb0brx
JYPuxnDwX1uXjwvWm0TJpQza5F3WXh7Tav1MuGV2MqOhN4uigymsJYNolbC3GmktfsxidaTly3g+
PPLawnx6UFm0sYaLJ6WG2qWtWdwEw+ew7Hbrci6XG10YNVhJrkAs7zhij5UJCZNWvKr0Uw2SbheD
JcRLUlMYfqlRCoXYadRq1TIwdjbANqy/gvr9BYFiCgPjIlZ7WrJka7eexDiHofN4l+iixkZwP7Of
v0YgGGfr58qxgEt0qoJavZGAvdQX5oNgo+jl8BbjkcMaveaoGEC5E3cV63N2uzuiloPyNegtFMlL
oDcoljECbdBxej3xUaZkjsSI3SMetDzPApuIrbxPaUHPGtakGByLeBkp1fe8E00tgiqO1G1jn1Dc
jYJqdFOD2owCCLsaFtnyZj7HBREhNnHcp0bu+nQevNJta7X/eFsZlQLKZhXF7uPdVchP+0Zu88/I
DYofEmB1vEQM65krkMmuyTnRB2/PdBbcCl9T226uabQVoW+eAVsrpA0hiZyAked0U1yPbDkxWZi/
cS1Z/KfOE3aJwIeBA7LtZNeN+07YOpRJD2ATFD8zCoKjV3t9W8STJnbDZ+9JMHVNfTHj0ORBrCML
zchWNmPDM9U+LdjLvlwqIMGxRiwIX9zqvKyZPhaOoRRwzQJOEFO3sDpArHw6oJa2Bp6Pucyk/bFu
mO9SeP2Hp0cC0LU7hPmXWX8FHdC4/Mze+tKag8dWCUnXS+go6L9P2slngMnXnXi1nQhPN4v/qxad
Ddc7f76RWnaX5i7OEYazrRJeBTDFflNkMa6MejwipWYxiFreTlb7MjurPwDfZEpFZZJQG12LpXhU
1hhycpTqdjSQksViifLEHmZXzWcOcY1Nb0fjzMXFGaN6NLgqU4F8+hkTKW4RMOGzW+x36HVAECRO
XoOHDsgQmJmzqFmJqYt0fShPGNzGTc5vZq5KeIY7DsqfwACeDeJDCKJgs9IsmN34eWO50M2H11Vk
qLIATQaJMk8a9uWFcqBOllqrXWfZE9Dcu19ZrcQvwwQyQl4wKLmfZj2Je6azRxQxACDWSySMmX4J
r8Dq+bpoygiKW6a4GV6roDSvY/n12YeMgq+HHGzi5oAIiMRlWW6CcfPhNGwCK9djrAiOhxGEQ8zc
snCc/DQVAuApkzmtoZjiKeSvCbp2pBeuC8nFIF5JRefKizxrCbZKhnMzdZFcgUk9APdletuZF8cd
EEPIVXQEup6qZVObOo/rpsVxFEsMA6ScJ4J3tiKQnsLXHn9a8dsrNtecHB/Bbe9naF30ijsbpvFS
IE61MFZfZUVYDxUjekTUrWhQ1NO4VOCgy5azqM4q7/Ob0ogjL1ClJsWnd+7C9sFe6Sb3FIlsV0nb
jq5tCSMbEuMG02TL1TQJhNauCLZZ7+173KI7BGpkZz6y4QoUuexskvg7WBei7ihT4CYJPf0XRr9X
CrWwQzsP3UDprBwKYR/RIYAoFe+EcalmQqDcApzV1B0arNBxfa4y05LWVB5AgsaaLW+WMeoOWZcs
sMRvAac1X72taZAEAdP6aCVMzQrPNIPK8xMpCUtpOliO5MxOBqXiGRqI5V6jiTHk6iqzmXixY4On
b6lPN1s0kZbwCKpX/GAvjs5zUiMRaEv1E8ZP4H2K5T+8/Gtl0tr1eyiADkDbbKsGo46FGwVWOzIV
hcKZh3uSaHYjVDRb0k5Ie7G3QHHdbBN/qcDiBRJ9vMix7ODcxEZUMSHcpHyS67Ej4b7yXczlnEM5
9nIqvSvuEF8jvWQSRAaccBOtJJN2OGDnlaOAXdFXvvG8BVDOEFc+EwPO6p1UecK0dz+H6dU+jj1V
7wYHTxm02lnIO3kYYQGRWSEXOuuqL8sDltie46u6kpnl3BUI84tLOUqu8YKnthwoG+Dvf3f5FEQ6
z++kmLh62dLfPoIsaGx8pqYiAryU5SEup7T/yiXHZETLN9dSUSvKb+v1abLw7D/6mQ0saTSsRM6l
exCaoJpkBnoZxN2uoC4ZyqeAGx2ZhJwz6j0G9w1JahNCaZi/qngQ+ksPYdNtGdJmcCxbVFNqEnsL
mOOu0ifBiUhacm2H416ElL+R8UT3aHBoVOMhLSn7iXW9CpiFZMXysFE34VMkk4qtvwxgFdQYVm+o
Il72vHKOOC/voCjBGyLT5d/zMF+77TA9vElaBqGFicEBErGhPaOKRcTWHZ3WT4efwWPIMHLWwYq4
p2yrTQktzQYhBqc6iuF0/f0B8DO+DlqLcfa5IGDVWGveQl1awousqMY9LWNQiZf5P8iFDP2e3Vpw
Rsu9Zk68dJdGyKjdacAsdmJtVrBBkqYVijPwswy/ddk6GpMi5L5bdOxqA9qjoZ6t1esn0p4Ivs+p
0IgeLkcmR8DbD9O4gRB4+uNT0nd7+iVuCrHkh+jIdQJLOhgH/Qb+/CnF0lm/AYbyAaMFHj5pIPZX
4F3cR4FZWcZQAYAblT+liRpFWnxSDD6aJfTvkW4KeAnWreFKJ6tKtYsV51+rri9tAUq8IE+Db9Y9
vdYQ1DChMkjIzRqvuX7lJ4IGwwNzKS1gL0KW6j9WPsAY63QzGcqpNy+osPQJ9qSIdhEeP6M1K1Ta
uHJi3YtipUVTiEAqdCyH6oHhkJEHaTrwNLRJJzLu+luJZN+8W5gGo3hm/lc8lyVjaddQY5l2hMmh
+yw21mchyKmalU2VrGTRcVqIAtB7X3jEjuFGwg2Kq+XJtkAPwYSXip29Cgtsm5jNSbPqGAauoKqh
u3/1NFRJGMgHewVa4wXDg3SZ16PDqUnFCdin2C5/EL2PRtQArTIltZq1wL7gtQmMlr8urYpfeqYG
lLsnXQ63+CaAzc7vv7PYo57KJyOUJiSANQwsZWbDR1e4Sn9bDtnBrtKK18VlImeA9NUbrp8oTw6a
qUNcAU9IvH+JrDkl04BPuLnoeeFyP6kRbzKcZ5lmpLxs5Bl4rd+VEduE7r1+iAPy41WO/zv8G1ya
yj3b9dxVNoNivNrLW7HHm5YpvyBWdTrafPqSldK0ImW819GWz/k44WFxZoqelLer3RuVjt08BjYC
XkYgFMVd8sORGV8bPtalQmNXg13QUvMe2SGei/dw3ps0s2f3mwfZTWffKf/7pcU7muuV3EjdZilf
qe5MIVV8UWFIs2KFG0GMdIk8Lnxl9WaZz6K9nDTE13hBXIcGeIYmrvejWLvPHBaPPTiQml7Eb7bq
n1VBtgkTrT6BUvZ+0O2JzvI8SAU+Osd9wCLBlHkcFblImfoAh0JliZP8WdKrdmEUNVPDZA2DJNy9
JBso3VwzDd2YubxR3R4RZY0eP1IgEGIAZAnvwgI3M2dJp0z9VIGB3M8Wn7eFjhPvRKp9d6PPt4Dk
DjLEbA1HZrSOGMUStstiHRP8118tBGUD1vNvz8oZr1H8Yy5yjomxie3IIqBIcTovYnvG9V+om/k3
wKrtuIwQy5iB9LXoCNR30LMw/kViZIj9e7Q39EyOugkID8ip5b+c4FyXMzjuAr6IdVAd7g7LFf3l
siYYu/zKKIuBPFd5Y80u+hxnZeeyYIFnJ5Y8sU5oEsemkhpOFQPcNGLqCCGMORIIAz2uh106LsYT
iSo22bJ8IBlx1KffPL7pa5T3mSbWr6jYT2bS48SqI5sft7CJN/g/E/UMcCxHGV0AjJ12GFWlheYI
onmaVZU+LUrsBrURb2CKgEQUWkwEtNH+m4R9YD4kkp41kZH23TKhxbJHXQk3RfjtgS1z8haGEzC4
4UIH1b+JAiQAMHU38TfWo+AifwBEoPc8TCR5xKMbw7EtAMuf926j/vyd+sTv1R9S1QLSgnNykl9p
qWUUbXvn1MKay3BrSij5dPJNTcgGFk6BI5b5wkU07tOGKexujrxxyZNoKl0qMgSTCoB2abbdNJbq
k0Vhsq86blTeRoNMAJeDaRxQEby8Exa4qMi4ZkzF7+DNw7aH78ND6BFcegn4EcwsFnBhpz86JZIP
vcs74ItIBGN7TF0xlaeIu4pFmoMuhInhpY5OS1IxsNYrTc/T6mD+uNf+fnm5uHuS9QHtltvyCOg2
UUlABYhN1+biQslM+ottMGCXp9eACkF62jdTXFMTqkbThWeH+cYryE2ZeLuiWXcwcFbfaIheRVP3
6+BcLsG+nqXdEe8okusSUITiSSlBjkKEEaI5qGxFgQ7fQwtTnHCmNGGvArhGpu4oqNC05O/sNZrK
YnCE+boMxG2t/rZiOBgI+aTV4bOBq6UvHO9+umCVB9fVI3CBCGaMGj5Irz5aJtude+E2IU8yQthq
Ijg5nrNqvNzVGIdXs7vUgkFpiQy4gmjp8jQeI1yQXQG6TurLrKlRLifJYeQazWvASaNq7bgcEONB
nipSkwwoMVFZApg/9RRgGYE/ktJOAa+8AIl8IqgMCyXicJ3vC/3ecbTxsjju4VFH2c3I9OCHT5Gs
loG7D7Un8+eZIylMeGNkn4eG2zL0Tpvi4ntyPigJSInRWNTJ5NDMBUFJ7T8kEfkHz6HlZJGdOFl+
3YNuX0HwUUKZ6m9rqNKm+c27vOjNVuGlM+aDz3IbjgfN1YwgAZB1WpxG6Lr8OVlH4izt9fFYXrdA
oGbS0nDaiH9EGbgsF0ymIX6lwAC6+itGF0Yuy1tb0dowOhVmKinGbBQxtCSvsWXD+grz/cuZNwOv
H/CUySCwtyuEUdC6aef9RxprDQiIQhdyE16BTn7X5cNZ9zJg54okmCxBBA7DzBHur4w+6JrqjaKT
lS9fRwTOSxSQbkdjp5xBDuOa77Qy/blW7gBpcmyH+fN3vVXx9jQWDC/jRvQluq3wbWDyiJVrLdow
7iBZHgqJpFFj6ShEvQb9ofOBk9OHRv987iNdELjTPMdBQzmbwMa86NSH3SSCi9v3xeJ0fDxlqC+Y
bb+FmBFYYQSJPGYF+F4B/Gw9aymoTIdir09ZmPDWguv0Vtd4Ul3/7NGxdHzAAqR/AIamp1rtCsNW
BkVTXUCXL+uZRS2sS2X6TyPVxaOTJ4wrjU8t/hqVuMF7ef8h0gqJwrw0tMQon+HNR1GE+6HhAqS1
Ryi40aind8kCUDncLuKW/gFFiY0tBTtK1zob8dwPPp5DkpNR/XYgVgGOsPiuhTAyH+3izY/bJmKc
BZBDATidapnta5AzkfG7BdXTiFV//RnY2i8Fn9JSdconk5JSTTqoE+woDNd8o/51/J7u/MNUqMY5
+IGMbVHW9r4F0i8vDm/t9MOiIIygTjr+Ej0SKfK2R2L5XuGrcjFMvt/uF3ogKKBwmX0RDdo23NzP
ew4CkCrBYvbJMUBfrj8a7t3IU9p57FqBYgbVNKZp106u1Kz4D3XYHe0qwEkFcb9PgD1Y+57JDwcV
nHdSZxoZeRlfN3htx8hAUCSbWFV4wZumgZR9MlWBYQZ0Tb0+mJZrz4mL+N1bB2z70wtJcvsYeVaZ
xyOtdN9z3EQj0WI9hqb13D2A9yL/Oq97gFM/II+4+2esImoKxZa3zqc3IZJrJ0c23cMWn18wE2WR
gFggOzj0bVnVKR/8eT2qF5Gfe/HAmLgPtNXZT9I00x+72miJ6XyY8+h9a1Hv/KRu6LMUih0DEURw
neUdCWWii8Dil/80dfs1fhsmOZHHX2pqw67hPK3KCzEv0HvWP60OrFvM+6nwTSZO9i8i/NQy0jsC
4Y55l8dZEVH0lpM9OwgTLEZlLK3tdUSPj/oZv9KaoEuSBci0KV9Wn2JTC61644O3ZYYUbZ761YCL
KnyWfiFitiHzwe7xPW64FLbINJqnHNz1ZKtOUdImM+qyQAxixq3mMPrNr+32HYMzGCNjjCKA2YDh
8urXpOdfBj7cXXZFoviz460hwCMd4DLZwxFTdcpNyuDjq8a7D1STM/Qf6KgZ6Ro2w2WZZuMxJLEl
C/AtgC/upZw4daICqAqEdxOqQA72g6FfG3zI2GVKBoNlztYyrJx+Vd9Nw9VijGgkRv9QUO/+njVO
t9Cbm8MGKpJA5/aBOutB/o6hFi3J9oN5kSCSCoUO4SiwFcKjHIuQYd0tAHJRS9ToFnzZhXMkaJZ7
zm5OUC54a+uAV/z4IAHCXPVhO1VW2wQgJyBn7H/9JBpc56YCN80xgF3RUDcebyPPj56dciTz00y8
5Vs8AkQXdKBXkUYS4SdNCwxGK2JphDJSoFa4oZP7CPDSIq8ZfHJyNkvw5nfa7PldXTHAYT6VVVhZ
elDc5R80kJfrhrsrsYhTG1009cQtki/dIm75opJ9n3NoVOZ02iSm4nkStYh/zzzk2aqzUTe1JUTU
jIz9VKuiaN0tY91z8KSQU6XzMJejtS6wA+Wkiz+bsKorGd3yRSRteXFDVjXzaLF/RVH6+/Rdg5e1
WHei+JyJQpLl8haEu5CRM/pCDWwdYTfKAcFwkky0uTXjsMD6H8Z24X/Hqdan9Q7rP58CP/mX3F1K
8Iei5F8HWoymDfVITE/NlVyJ114e1TE/9ScSd64p+R3MOfnD7zzoeZxGNNc2bvDZG5QzjYLlq1O4
8I1Tseo/TiQpeCKvk6swtakkjlDsIvli+bV3ONz9Gk72RcQN6ziVdx70VvaKc8AHArDxDE02BEK8
Qqe3P800VrnF9NoxGzWUUy4lunKgKxyLiSuNl1wTHnsTmMQGnbmyZQcNaVkLlL5d+LRox0KrnbRR
jQ4loyoxN1g+kOsV/roWx6t0/wZzl0xvxjAjA+Nq0CZXWuz/nqPAj5VcxMZZ8XxE9cFRfdZrrdAs
YOVT4TJduX47OOoBxBiLOM1jMuaKWqdQpfj9NoSqcXQjZWT2o65TIKQx/GcBmg+rwOavE4WVF5OK
rGjAzLJ0zUiYumHXTxV9CWMIeAkMi3VttliT5u1BNSy4vHtC1Tyf2Gf2zfDGMJWlgfUWUpkSkQEP
MypR7qHqjSTxHQPvjlc6dn4G5Vd84R+zuB7HdHgtYxhHc56ESofWAobT/xokGOd7gKIEgdHVd93l
4qjaJuDcGH1D0uks1PbaGfwMGK3yzdLXVZqM4stVvT2vS/0+C+PNZKKxLBP+7aX7xaMIptn3S0O5
fdBuqN41c9vnN94BfI243jjasDzodiTH5VofU7KWACxT25Bnopi9FWLtE1a9QE7V9h7sXQe1iymk
Tee4EjzFxhnSDFniugMKvYgDuvFyw+YfsMJvkve0oR8nwKKe8wU/ByuyaAEkcf6acXfJSzs/W/9S
fU4XnstDlAgfDOYn8+cBwKQhJ31YMFdBuv3IXzN6wW0gwfydj2g2FdclgF2fQUQoYYCzBF3OwlAN
UiRk3iy95tqehZe88Cq+pOhRHcWMwN5Xz8YizOvuKGXYDQOXFMIhjp8iaV4NCMk1KxQ+44UtnW0P
75kRKfn7jLn5CaMTt+9Cp7mii5p4ipPmImM08csgeYRH8f7U1lPr+cqa3NTsvdU0fJzy4Tqn9iS5
Jx+y5x77H/m9O7Zgt6KCzbEHfnhvXnVtgXa09PnAPkXbE5SG7wIWBkBgceUZlaXvKXOlFSJsaUZ3
deQnfyRU5PUEhBNC/OW4ByQ2VYRuJQFqObPYMf+uFU4eJ5tZ8gd4GX+7IkmvDE7YcY2szq5G6LQ9
hLVz3EXxFnHZWNmoWArsjAHOhx+EnQgP0Vwect9RzTHrjr3nVhjCLjFODd2OqioyqzGGhDlSz/pA
GD02O/Cma/x1vu9m/qTPpfSW9obzwcb0eex61w+t45TkBw+tzhnTfON+lsFivZiwEm3jIFn7RYaJ
z8uV6LlVgkTgR8S/iMGiAeW4mAn2XG/qiUcIC0d/iiwQvjqMFViAxjMz3jxA8ExSXGEYFVHn14nM
1LNAqQbbd3Pqc2gk2iSEaxTaD7/vlbxcnIC/LKGcqRnvS4tFcqOXaPmA2oR9eBxFfFw4h1VGqrk4
cO249SCqyxI3Z9BT5GsLGp2XknCqdDj6m2IWb8EznG8VGZYLaF452R0LCD0oYP9jZE0ukZINlWVz
BuVwo9HiUvYLvL5xzK0Lw41BXogFgAMsOHq1A4cqkwVRkpgKn72/TYwqA+TpJbfGThuEh/GgE+ia
jAhkUTQ6L8/BYgLjJXfknJXWJvCf2+CPFzioOwaPTgGc3b0wtk7JlSNYPTX7UHs2UYLf5nLauxRr
bvBJVQbuHZNZ+wOYcUalPG17Xe4iPxpHlHw/iKdERsbxmDVjEE06ZscksW3bcAo4u+DQnbYuS/E9
QcgDIsA3PkG0Av4wzVopKy4/VkJSVsPJHtjFs+faEx4kbsEPEFbNFo9bvATLbQQB0jxp1TOGmo0s
qnR1nrn58rS6if44STxdWlpjbyssdoXRoG23bdfip1URA/kIvG7MXByCbzftRklITxnj8DzykmVW
nKEvEyKVU0UnICxtoY6yPxblWi5yTzzIWi7ZxBcP+a9DH7if8yIDwsthxT/pLaqLV4q69rDOvBi6
plFQUmkDnOyTjaFRWQeQet0c9wAZBSl4AbGN2wGtfG9jEqtxskJbMTUPFjiE4xV79+FkBUB1DBDu
SpAikMgfFFPKY/XKJS6Hy45fGQrGlQYcroqhuCO6HZEs/nEykta6hKhAE3qpoNCAe1nq1dVJYnm0
ISUX9b8XRUZB/EuDo/ecRgJbM4EQGMIYA+5zuT8HzzRy1vz27g8F361hIjYPkxmjR+eOTAGz+EiJ
GCGyeMXdeLnzwIyCrh5Lw2tQ3N8BC6jQGPkfWrDjc909b61hfI3S2KepOWNca8Nzdox80B6aSyBt
LkE19E3dqPlwB3jrN60zaJsEtvaUToYuP1iH7CYk54DIzaRef4hJ43Uw8OmY4bNTX89diPYHR6pX
PS31N6sjqSGiAgGbq0nc074oGqZNYCyZmbbh5JQ0/F5s9cTSbR0Xf88il3u4BzYavfoIqOSp4M23
579zFUahDjTVsvGrk4BV/Tl1TMBU6NWjslSp8RBxJd7SbAKNMa7yh2ipejZFcuqtnPJP+k1SgNXc
iUr807qfs/GdiipWpbmKYvIWK3pLMhqPiX7QoBBhn/ZU9TQj97xUqCqFqmC0gB10URkDXhydMB3c
CmnKZ8hSauE0flqt9/J3t0W3b+SsClOmaa3LJcW6WrhzlNTNfyp0ENYir9xZek3EeI8e8c/Q5qoh
aYYC8IxTIRki2/xD0h01vNdvxjVGbEQBsaza6i93Csr+V9qGPjwmmqmA3renSIz4fV6CMClpnhTo
33P0pvHfRoThszxP3DdPVzqrq+micmIPSCKTyz81Rkql0UuSa8IBUmjOWcD2yZEeoRiywET95IhD
cO9b88gatcdUBANs8oEN6qCd71zGEwRgVT5nRVDawXmpRfn/t9esqPZnnZhkZLIaS+cEl9iFArBQ
Huh6hMocoiJUXQoJfPPTKBxzpEj7MT8blREY0ckxZE5Jfw+JXCSprGXZtlXEzWiOEpEasXG7HHLR
ySGODeoS2Nw108/eQFwBRQNbU22tNRuy/5XpeyB7glayRqsW8ket49MWzXl/Wff6uG3QvSqzZ142
LMT3k2IolGVEd5P+BXQsvEBWrcTjfCsr1yFFsCGMEjGCr2chuLdz7x6QvuiKQwSeo69PM8UZEnqr
v/ck0vPsS6iQ/81Mg6Me9eCAm8oC/kp8GIULDNQqhKghv+jsm7vfBc9ycSd/2l93SU872XhV6MO3
2/8Z/T95Dtd6r2BOVU1WBOAR/e3EIjI3bO0W36Fchu/cozz0+Ip5ohPE3M/ljdDPd1AMsObB1yfj
ckgbpNjlHLLNG9tn9lYk0mv90W/jzfRlTVSvdPPXIwnem+33aZT/qJfogoH25iPxbQibx8pQzdhU
1v5cscEHHo9Uf70OJy9ZKJwlZ20ypvSueckG7O/GyIy5hI0RwVCw2b8CNbrgvQRGkJ3y5ITqdTzb
7eoGRMlzJaWX4H7mKgTX0R5Y4Q7LyIIFTBYOawHucjPbwIOySFLkS+JbauMmvw0g1JApa4Bl8KqO
jcP1ZmL9Cm372jJsuUEjrlnW3wuv9MkaZcZbs39m2Q7s58Di13oZstLWSS/VdpQU3fcr5+lgkWuv
8j9CbZ2V2zKq1AJxERwO/LQqiT2++e9o4MfTBnwR7hZ0cV5yxPPRc+thPy/G4roi7Ewl45Bw5/Go
Nuj1hBpI3ISi27cEYGiQYibTS2TbphTltouMAcU9VppoCIhFPHqxtML9v4Bt11xdMGmOCMpfzSrS
yn8xLsOB9TFX3EuYcOLVklCDxecLHJ8t3xqr3P2uzPPQhCPN2FFuayc8A33sRfFoIXz+Vvy4VKzN
EIM7iso1f8bPN4PxmTlSi+b3c7/51CL31OaZT/ZYmmWIx0HYQXnwxgwcd7A5Xrku9GQqlPK6nrcb
9IbrtCIGp+Q87k8rJkBw1NQyKUOBW1RY0g8G6dueHqT3spRZb6EHP1xsyVhWlU3xSLnmZmbSXtrW
icrmE4m2YWVLMKrxcYwPz4pzNuqMMLKD00LuNqZl0i0cU0J4j67/Cp0b4fpmXQcXV6WVc12h0QNx
mFEV78M3af+l5vrOPpGjy9puKeGsTs1s+VaoDEQFxbjXNyNteJF2rd+rrXBDwUDSxuNBzHFxkVj+
40ked7rqJ4mYxmkltTwQ2pA4Zy74bhvLbr5V3QrNus0pJkAb8NV1zNQ8xLJ0q5nXbklV5ktsoYM9
z5Yyw5T+iCbNWtkc4HbwXYDYvbgScp0W7haZUdBmm2E/GZR/pKGyXNwbBbXtgzs7LlJRugSp0OU4
9763gAidGQpaHbFDAVjKAlk1XSHdCqawhQGOMTwlS+l3inONFGecbNrxg2/6SfPtdtjfgSV6KBBd
1c5vVN/7FY7lx664OjI6Is2ZC+RBimPv4qDYClDGHUiCHoXirWQ764VfUVZu/Tu89qlF2kcS83h5
4UK5nnkh9NN1QCCQVmoyPEuyZo3KZaSIkKKHouFTgpCgjXKZbdsxWibvdAazkTG0k2MI1AtJzSAy
IJGq0Jz7FQGuqYZW4wH0EWPY23nZFAMqOCgxikkeVglmxY1+TzmrSXGP+3qu5DIzzfKXXgLNRmjm
lpvjlSXHeNqHyQEMWOXG4BgeLtx84wZOm0YyjqOmfFhHGJlFI1c4tXH9lTYZ10955v/K3qut/eSy
gl0L6Y8VEtW6hpeVIhhdEuM16OG360fpoetkzI+DmlzRIU9PmONtpouOyMALQ0F+aYWLFRJigOCg
T9tXwEbrESFcjuxeRbsdYvTXPFQPwrs/35BXVPqqvOOuUFb33NAWn5peTR9KSdYwtmM1Th5Usn2S
ZunAheoJrG3PJrfmae9/XdP3BM6MAbWBjyFI3ZGVDTZmDlPgf33bX/7xa4goYVRlYBIOK/SGPCAf
5iG7O9mpWp1c3+w+SGmvsxLKfiJ6gBeKI/kXQkXnmyTq8Sc59BENwmoa697bTBwBbJUpDrakWMPa
xXfNl5fNTHoZUksMt1cghaxZamGMbqTNdnx9pN2McFewQEW6tvpT+l3FEDoBK2nMQgNgU+gX1e5m
+hMNJmfU1BYgWnHixocPxXQy8cTjJXdSzO4LeDZb4zET8DsRybTOAR3b5kcsQR4bonN/ulUyA7xh
uteAHkId7igkoj2FsV+e793fKs4ad2XvLvmvHdjk+JFkQUVJBG6Rvsa9MtqiJVdfE0vJ2jLnBb5P
yH8lxxvJ1CPDWGTnrzgintjERolEQMeC4OHXbLqHWutP2ffGem4ba/HnEIWkKUOB2lIb5/RudH3s
DU0cFwCyridjyxDI+L7bCKnLWN+p1bCT2q7HUGbHQh1zyxolHMgxI8iKo6T/9d8XJRvDScvfpK8a
FIgbSN/3Il9n/Sa7PTtxR4Cg21gDACQn2/8UZx5JcN6Xm4aLhlKQcpRM+onO6+EgEkFYLnNcluKx
0ZZP/+/I2wwucoMAKH1VN33dZk92U6z/Y7ivrXaB0233cr9AKbPjYjbHG55NLqkesceiAI3lcr9B
L9cZRFqLnKdjegq3lkOA8eoUaAm/W3qCsRqy4cyisNDGyQaC9VGyiYv65tLzvCdfIHIlWTNdTKLU
GOPFws804H4Q0nFkhG9jM57oQsUsoMMEgybVSKyHlPwCUcPmi8QI1jyp5jpA0lvwFOXc3lNT7mf2
gAMGOwFfy13aJizNN56h0PNghZLAbEf8fAQ08QRCrbYWIMMtbEZeXBhnml8vjdXb8lqQ9AXH4vf3
hLsna9/CdC4mo4n8i39SzE1ji9HQsFKAagdLjK4VUHNbRc8EWS/1kMiwT140i+yJdaTd0itxsYJZ
mRURLHX0D3gQTP73/GbncMR4JbJ6Iw0FMx2ZqGN1M0kxsfurBKkll1Kox6ISI3U/PRps7sZPFuUP
3jrFzOFicuJPZVlM1bHB0ey8Dzjw8Dbl8b1l/3pqRqYZhufIIU6QDxAHWZw4/SuZjsE8OwHRRM7H
o2JGpUZyzDKQumk64faLM1IJDdG/6E0kilvN8iJZ6uupPB58x92IFPUOfbN2U2p6i5w5wByE2/zL
PWAb+9yoZqI5NWIzSE1THg3TlRTQNERbZaTO2dBzIt8ILYtICTvAB2dqSONFrxX3YpwA8j+A+/Vp
QquneR33AU4eLxkPOmxB8bdsf8wtfsrc8hrCAiU4/E692pi318ieTG1+DhQGUqyM/ijuymtxHPe6
nCRQYHv7u3VXH9onyMkeEew1K+rElxxAMsyzWXwghPJ2jz7HgEUhA+IhSFiJbCb89Nk+cf2x63eM
z2KAyZ1UCHOBjXws3vRFZ/GPxyH4GDYlZdjy+G6F8xSD/oBjgYIs0fq/TsnoUPrwKMiqFiwUFUyO
RRKi15LVxhE7ryB/3R9RqTz6VVQPhjAtxWXv78V/5JkHfj9Cvp2vpvqVyxt0YQ+gxmSUiI1Mp/nl
b2IEcQ2m+9bQEu52lOZsx/XX///iJvSthxbqtJoQ1OFIoni4onRrU6+s+wi8OXUdfcmr9EkSiJCs
jacLgx5EE8AJ9Lcd9GeP5YD27+7PZnKDahI7gTxY3pW4rLMmLFzA+cSGEc8RnDVY02qC+mpsHnJb
Crl+riSjwBFuhqPyk+lI3B9gd6t7PU3U0T1EV6akDPtFzCqZNhw5eKnW4tgm37gTw7WfM2Z6pLYI
YTHWPoetw1ovJrsDHTm4WunClFLn5K+avxdVYUChawjlv8zqNAAyKH/dvD3jusOqqEYDdoz43LF6
Yo6bY86bbaiStQgI3vtQFn7G7Xiemy3VMSZU2bG4dKd8mfwlAFcxjNX9uxGoDm78ilrQ++gQJF6q
opAnf1tjcvO2Et5/f8KxDJjQehsQXm3H4BN3a1fXkZ+LFPNx9CZqAC3NuVbs4HI6xazRcCSWWaGp
+HfPXf0JTPTl67dyfRBonFQeRrztuq0FQ4U1UlCq4vIbuzuM6s6La0A0fID0xEK8IzS5HLL58QGl
0YHYHsrRJK4rc0IjBiN93ZpyOqbD03u6WlbOJiDWlibGK22RJKAxttxT8rE/WS4Fjpun7+IkpY/4
EdygcUhpqLnVp/38kw7WisYAmnyO/FoiXRXI5osYyz0hXtUHHzLRGPhFslIPj+mNoU8xJfA1lUJ8
GzoVJ+lpRpo0Nla5yHM3Pk6/MbnksNlGrESDf1OhFk3JYl6vzrHtF4SEu5nJ9GJiyFhEvGNNKMTX
NwUBHU8CbOhmhl6+d1LHb1uO9TKqyC7gYYS/uIeZCicTP1mxyqVkg2gr6ZlN7u2SAE4w2IiBtx3V
/Cu3ph/tWM8+Snl967dAZJ2VfB+3Uaeo8s/WaesuBqUuG/bfi8roo+8DLH7/z0jbmXnwuoomvGEt
o6t7AAoPH0SHRCJSLQQW5BfXxyzl0Q1teg86ZOFf9+dyNffax3H7PAWp2P5/AL95rXhwvxkzC92M
UJQf8vkXprOOq86bpd/lknyth+Ebd02KAjaH8q00ER/PCp37W72v9kNbTwn8iBDKHSx8owqoQ4an
lBwsWe/e7fkY/+m6fAUUmiurjPleqgvLiN/mAmCF21fxqNgk8IL6R0YH/6F5jbtOt7siXU4cGOwu
WU9bD+n1Lh0t0lw+/+dpccOGMuxbpYeVEULW3DokTbTI4WJZxq+3H00e1G+az2WeoLB4Hq0r2/Yx
WzsqlhLp29sb3FpJbIHjjUKt0YNuu2K4Nn0LVK8Te46E2FTPgy8dFO96jo2f7N/wOfGaL66W+TfZ
9D/IEeS7N86B37kMfCH/VbcAt7ic+DBqkXsH0ehSReh/JpNYYYTkz6POS7xZYKqCN+3Lslnlt3UT
8S9jqC+Gyb+sjDiU2/FhPD4LyFonL9Qz2bc8LE8LCp7BuyZMD7PPM8yz46YhGoIyO6cCDRojdiLW
6htEX2O8fFrSKqOFziKSD2SJ1qHzUfO7JjrW1X0y8pFsu8QISSlrPRT/aHBHpVUYkOsZGwLTdb2e
GP/CR3b0klTnTvA9ZCk8OwvYyzaOQ5AyGsMuNUX4fwQjyY2dG/KDyDOVLH351cTT1CYYd5RbwtMj
+4sBb2Bg6IJE4LnoPUEgH00eW9RfspVPatQXKZCjOUHaGElFO9+r2fYXO7QR4qW5B7ajGKy6uGcK
zGepSfKdVvuDSjbncOXoIGqwOg02VTcxr7pzYuHMoMGbnrqvcylMMhQEmNmFF+9tLktpdSJyeJRC
aOmwV07DoYvAWo0pGh27oUPsahx+PADV57Ox82znpk7VN6c17uuLMaUiaQvERD7DPQlLoVf30ctX
lDv+UD8hUJw6sZwrKKZNlywpcEIl1eMTe+70JprsEoBxcIXhB0mbu13pAcy47riEjRQAfGaAIAEd
FYzl9qkIXzuZAi6uckPhrIoUCry+zLsL9HJJ45rW1TnujLsMHQqTdwNYika/y2+qJJcuCXhMzFyp
F9DmX1sI+Pgh6OZNVdtr93u3Szpkc2eWTU09kphCfIvhtP8fB0dht0KpTxykoEUOaI3u7g7GTcID
xfsFzi4DQtVX/9eLaTwyVyFCVH9fMSwbVD4KzaLmt+na6ATEK8KZj0rh4D/EBk/1ZAAlIRweokXv
bbX3LbSOlYxgc9RUSvwA9OLrOPWZOd7VVjyiF5QxeV0+QkxP+bodPys/S7wiRdDjrtCTKpy++jFQ
YMimt49Oq3/jjr+bQa4e7akM6G/BQKcJtv9l6vfySbCHETPlpSLKnv5G1vDGmGqUz7fpqPhy0ghU
qboWN9fE7ASs/WFDKKW6YWDqh7snzK0HYPMSX/gWP4HIZ3RFn9+Sd9ONz9HAVjLh/msIvStg+Unh
6/V972BejCgIrelLNI14laR/GWx5lf954Lcb1sRWlWi9M/gSNzyDo8t45X3+QdyiFyve3pGuPmRb
buAWQQUTovD9xjiEWQqafqpBkdeOpfsxrjbwalsz2yVJzj4/NiPw0HXwrNpI2itFGVnJCga9cWza
M5XvtegfCrzvgrrmdr0+CIb3XGrjl+w5UvV1rpYQ71Blx9JKinRynp8a7OT6Rwg90Ll50Fp1WMt6
YFGLY5bKR6NGbrgz46SoOaGtoN315nRVBTezdpMBsCvA+R4/4cT36A3S+e6E4k5Reblrj/DgAB1+
OmBsMS9h+AW5PISvkbgkNqylKvkXDqIcL3cJuzPu0SlNY/AlbOqj544VdKsrEztRoDGMXkRMPKg4
73u4P8IJdj4zyinhZCGK8fHVxomb1p3tnRAGKaZQ6Rg6NXFfskX4BPIW+tbL9KqCL3+LvbIg9woi
qWHnCrnqcq2cePDchHw7qwz5aGRaHY/ASLJJoYui1EF5MkThCxr9weBjaXaI0UdSyZKIyiNlUOQo
noZIjFIHv9sbrD2JoOA9RaeN+tmKSfHocxgubTVCzl2N27sbogOF/e3MyUkkf16cvG6MOdMggPzj
iNM8k9eIyK9scTjnjAoChPE5jTmF8ekeni/lGFa1y5knnKI5hvW1Zd9y9tn/+OXGjD97w8BDEADh
cOgmidJGAw1V0c7gc1woiscwqKkPQL8VeQfYQOr23uKkq3Mv7JyfBNlTb2IzZy+b7ik9HgMYHaqV
GkkxF4rggv4xG5SPwUjSy2gDAXfNcXLxHQKxxbVY1pYsIHX4gspz8MtrXIhyh1Q4/kT97alnzfsH
JFsjDzob6rSjmo7KL3kjQUe8gA11zTLZzvNhk9Y3XArHXQeutBCx4fNSWHTya3iVks6r86yV92k5
t1Gi3D9+8l4ZKg1m8ZhkiNuueCdqLXhE7LyLBb/RdtO4WfHcsDfqhicDUrQMIEpwMSsFdj+y7DMt
wJ82unNY1lYNsCJRYzgcy4owrHOUfU2pOLO7PjYT74jb96sYkWz1w4lSokZoiv2iAO/2oxMxLA0S
GSi45v97227yPuOu5oVThaqKoAk1EcGxcFrkL+KzdHV27f0gwdw6wvxEWLYSfBEtnTcjLo5qpa6f
UquE3TrRiYTmGYTWQdys9dD0KPK5/ORFboLFDJfcsYKS1pzRAjfs3QwiKcRCrKh+RlvfE07i+q7o
F4YmuG3gjE4KcGCcXXIXMN2kSAy5tw3ZZzsQQ20kezd3uXOLBCtOZf8UDWZ/oK+W4nESxQtN8XSQ
BMDRwOpl/nVBpWK+w9bPFSwjjc254nnKgSAYHYcz02zuxB8826qmk5710NJfAoXAW9JloBnBKHYa
Y4D4G3MBj72E42a6zkZNDq6omfSqhBzagobWUiG9W0+6DO6fJf+DjXLAA/WVqSctsnpvj2UpoEye
qao8m0CGsbgDmV/58Ft67HKsimHdF5g5E9Bx1PxyKBmVoUOOoQiSD0ifWPpXRQY8dVLPMP91Tw0w
+Iai0wTDAgzn7KTSSD9OBGKqolD3N1AIAPbXauMLYmCRoJAsqR3UELElkwEQLG3EBElz93FEkEKu
gIOs0VhfgUloYoMoOBrAHAqHHBhCIqQudP+C0iJid+MFZfRhF6LtlAPYcoS+6a5pnqbD4Ruqo3UT
+5W7HzsaVl5iT2Oe6MSblYV84Jn9pvYuQ6xodiSt62xyPwOmzV/ezn804QUfMp4nvl/tOfawFk9u
Ppgg9CKlByvhaf5/k3feI1AiiB/UhkxyQwXH/EOUymXmHvl0T5KQl/+Nc+PbJz5FfvH0zZcz01/j
RQwXor8m4iWGsdsoME/Pt1twV4cktjQZG5LJNFLarpb3A1KKYjGFIyHWCZkVQuzyBpz02BlR0LOX
oUXX+LxyTXZO0sruA3ezO7tm+kbvE/VeuAoNXVXVDdoyOAKOgr3cjUjTkPRP6plrCN/A8vT6j6Dq
X4zjkwr5D745HEQYCBGCNyEQ179zge9zlK83asebsuobp6u0Jvy5MiWWBR1Ix91K2D7b1lhy0Gzl
bcUO4KMvtiOPLkFBjhaJnjL48H1ybnrCowznxlwa83MU4q222q46GoNTd2cu6dDEmTBQ5d5rf9Q3
YgbFYJKSkEPMLHKdk0RCucRUw5gO3HNbQ9soc7obc5/jykzdwl2h+pgAA4OGVV4KPEcBe8Y0vJf1
ZHCB+3OJfliwPng46PR4iaSY7NQ2QERwMZ1m2QBMOqIkX/TeRnDAOe5wTwBFUgkkFPyg76zNKlFL
TpGALNu26HoX1b3ix+zEm3LE1LR1VHqojurDnTNh7FKcMm6Pd28Llgv6bbMwE1XeJzZw/em1F+XZ
F8sMhEhqfZOL9WYlYbXd+x49EKJooOoSEKaE223yao4gBRnCHXk+WKik5PIrPjygdja++8aVcfa0
5u8VktrxWL5xn8HWGr/WMY92415Q7ENMbGynSFeXwnG6Dn3T4mXMMI+2NCgYBinZZf7nbnfSIj8g
isxZhWjFLUyfBCDDFvUriuebtoqhqxvtkPLojtABnnyc+pK5Xa+WRFU0HUEB04lyP4xkazBsbTKN
yttciQTKAFs/VUQqHDu8AAc4ARqM2axiN9v3RcPWmLTNmG8g8VLQcTTR+ey9PPEdpfK8VhoBdhtB
lYAV+3bIvZ6ekCb6c9Fr7LVQfxIawMPE0DEPcwzHs9YOWcjeg3edoWOH6iIy7T84B9FswRixEsOG
LzkORsMqkJOzBwNzdlFaW+F5+lnC394T1Iqf4QwH7LAoxDYRNYcl9YqlYcnRljQFQ4AIMmfoO1C7
E7aylVxQZi44pwnO/IkGNi9gmLAYrXdxH5GlUeciJ1iy6sqONqHPkPdHlNqgu3iPQdUsmPyQTgdN
n9cXIpBT8vXBRtlINoJuVQZN53ZerwErWAdtylB1QQ+uyd5ER5MLwH1K/v9zr8/dd4whqkKxuSjG
wfZcU41cBcPeq1qH524xWZiVw4BhJ5+A/wdjcP2J5SyEW0+die88O8hlpdZf30dGDogIizfr7tzl
5sWbpYOH2Aw7JYtMBqDsQ1mBMphoydMPBWWECmblTsmNSIfvGC8wmZB891cYYkoDI8wWU0IYFY6n
J1N94oxya19Er8lYCcDqNdt92AfrFE655xgrUpJCbak7ZF7e/B5BrbmvmrsJBQvBaZoclLy0CcnN
IhT/QDTswYudUbFNPvn+Ch9Nl0tehWJyMMjo+QVMTjtQ4AQt5pjg5S9DfhBGQOkZJD/GseBvxfWG
dYysIpu1CKmm2F330VL1EjJEHQp5Xd6aQjCfZX7jU0xGx9zHXgQG8zWZ0pTgAa06ot4NLnY6QuBv
ehtYlvNjqE/7zSRv+zal7KqeZeaDsMN5WI27Zwm9MOnJ/xsLTuliCbXpJHod1ScB9WcBTvJkPzAm
TsSjItBnKEjpjJp5R+HnjTcIb8lYJ1f0/FFMX4bN+VaTpAbxiDD4zJfuHJ4Tw7JeuVgfdIk2GxJg
j2uyrrlp91U0MJ43drCJMFLktvgRtVrdWJPQPj1s8z2V3uFu+Bz2d0cIjV4gMINVk0bI7IA7wmXc
Ev6r9h6vYCa0oLTGCb5MxqoGv0LDYgNtn8zDmNF+LSewm2lwINULdwbEB5qt39GvqB/XCNlkKFH3
FtAclcssp9Wia/HykBS90RzYHBZDSANmntiICv1mzD87Ibom37oZhXnRc/VIL6Ea1BiZakG/Ssim
HJyb0cHFGqsLb31n1BZP/sGKCFifGs1Z9y0fks35lN8uEvbpspXf/ohzzhRBC7xqiZwOvjuVR2Xb
mLvHI6X/Zfui/EsZwWd/nq4RkZfmoGeeqSxMEAnQksQylVK1ejKw7brMLI9R9YOzt9kP1x5x6err
q9MC5rUBKre8tvGZe0+/FN7XAOCCtLrNRMHw9DoG2LKWYZz1yuFZQ22BjfJV8qHasbvrYgud+n2o
JRCzMdyIpaO2/iwVDS47gIme1JYiJ7P+NkO2SwcDGF14dJSKGSI/AOxnS3RScYtg2Ffaj3Ydnhjg
jLnXRpBaQWC6Y1UN8V7SXutRdU5dD4QpvkFhwoMLZH3yDkFfqiHjPN0lLis/4uggcJ1D+JwvQi2i
J6iOEQpQJgD03LLlChenEWngrHsgNvIWZUcwsaQDzLY8xnrts473b92YTBL0MTJmp3/t9oLFqqh8
9IAUuKOHNavbc0bC+74/usQ6xJ5IYKKl6xFpmdYhCcWwdPiWZGOwVOYFiXcn0XIRBGC11XwvxP5O
4UoZNmNXWo0QYSZCIdmo8lc3VZyZvwgn6l7Ir+qiX3jEFCsxbxNmi+971sXr2D9az3uH1+IMXhFp
h5FstRDKB90UPgUZVh5BEysLnniHHSdGvIst80tWigiAnkz5i2PJ0r/wdIZHEulMGAZuBouKbRqo
0spNho5jVUcAr/8/Yln91cR5z0Klfz0PmviuTwjZ5RyeEMaAetiMwa8JlwMc601EDK3mhZEfLXdv
CotmTOnU3iJ0kAv1Inp39cdQdkiXrmUvqz61YBKtFhd4cy0TtiYjQrIKNGBS4XD586z2HRlzFK54
0b/FgGzjcS0EFq9b69KgFpcnhv5EzTn1dLudwDZ4uquvVZmf/GUtFkDlCKDhe28WsCb18XrjEMOE
m/bXNSQq6eK8bXJqDUJhsaZGNHpxSNGE5J+je1z1MeqMk5wjsb1vgsCQrz9vCzcxfxmpRKXkAesF
kReRYsiYgHX0z95PX6BPXxiA2sMSEN2ja1YGL5V5Mc/6oUI4uMoBO9TvNW4dlH4NOwosJY8AhnSz
n2Pi3wFt5HctvaH/YcpmT/357s4Eb8YDCTTiD7kx6UwN90GgFgiy6IUTESWkAuN/Wz1PWTy2ZlBJ
7z/U0+Hamf+G8gbe8GRMdh7ZS1W2AyPcR7hjV2JXdOj0bUX7QRHhbXDea160V7tVHGtojUG46HgY
W7dSMCtbvWDVexLfq8EjI/IaVCeOkpAReZ1ILRL5w6C/H5yj+eIpD6qLerEzs9gDhGK1ON3c4VHH
/L5yz4fQVwB3qLJ80Zc/GjSKjuMVYY4pTz3F+YyZ8PFVrreSP3w7e+WhvZDvw1hfB/aWnQZLegSz
UB00MK6OHh4dCbOO5VcENFrvvrk3+2vj1IQ5GeWvyvzB+58+z/ovmw7z6oyzgJ6w2sMDvPXWuClW
QOfUE5L8XsyS0U1iWFwgjwMWr7m1AnPsqlotl7UJKgkuZMi82QCuAkIOI2sfNP4OznhC+xgz71Dg
+F7Scgq11eixWGdlIw7ieZuBM3Vae75JmwhFIe4lUZ3ivrzGDnARgy554D8bpnrDvDmzmZCb9ldV
43k9zv+1HfeH0JVE19gGuPO1X64S4T2/TB1HWW0srRp+7sEQh8UKrl4DtPRcZNiaNr3+C5n2qXQx
heXow1ORgKZ9rcSCPQIGHXJG1ezfguN9w0+AqkEyTTmRrf9dUE3qDXctwwWaFxVa3kKp5js+lOmg
/uk1kkpSLLdLkjV1etZlOcog8SNGd1Q1XyCJ7FtMeigMq9JFgaOMc6BnUAy4wKxxQZrr5HdHeRfQ
uf3AVjJ3eo266UTFvOYfV+X5COwDjuEoUac/gUSMH1/ugjE3Edh2lvFlUdC9fnJhM3Z5HSzUVA+j
R+Bi3dpTrKmaPRLnBqKZm2LXmbgtIVueMwGryWSBVoZsfwKgpTlqW5gtCvPoejVKckIX6g4iIEkM
GlgBgBAnMcJlxy/v3C0o1quSnh2kwRF1wyvFNxUxA/wvkoz/5j5ImPrE3LyENy32AwF/yrppMy/e
Ac7DLhzp4xdGdZC3pQhU3268HoF18tM2yDI+RqaZCrAzZNM0fnRfDkQlbNbe5KBCQKVgH1eZvy8s
fV7G1yuMsby9os/Ne/6PQcv127uq3/VcB6DHsmCFA7+pufvQfVOpE/LvJL/SLxXHGWNUt6tXAUy/
aEJ0GgOAXUE7JbyRGKut+hOoEu2bf7NM7qaiz9cgqwBFIoxJy/WMevEJtwgC4J+0BiNwy4HR2AjU
fmtZsxZ4k4IMRpIWT3b0pOO1oX97/jm2Uy99e7v2ZegZLaQqr3inCAp6BmQNXx9Y2JInMWk/h6nn
AJizmggEbnpXe8RiyKT/RWPbpUU8pTZ2R94wP7Jcq0S/9Ls+4hrP7lfzrNsGYp+McnMBtdnnKVQr
LIelp38/VLqGKlph+MK3bHjkz95Bi1rgkQ2CUMSuAmOq+KJ5DlXEzYFL4vOQmx2sNZL2pMG3dYln
e3G+UQD27EmYHowlF4+owf7t2MGdXEO2YHgnLbncky7435dj6IjIM+i84+LxoY659579RcC6OdV4
HsQl6WEpsE5SyeMwKzSbBRFCJDIrFBNJS4mxFvXvakm5thahu58GBSTPrug2qBs6m59NEQR3CGzE
bsav6w58bxrwvOlKVZS9b8nKthj8UmoyBfxc2YKL+HW6TwpGWjFWNGIynQvKBHWMgkJy1SyVaSsH
f0LPI65CTzGw9crL3FE6JNhRk2LKC30MqIkAM1kP3mugWx3x9E4Oa1VeujQKUct7GJipYW6NgoRf
yAg3RjXVCmzC6HE0FZScFPppt/bV8cfjJ3FQSkBSn1vAxiD/CUCcaadS6A2BV2AUj522oGEpcTwn
0dGgBJACJZQe1VgJBN9SZWte0huZBGZgmeJoS48TXPyW24kvXQRbBjLYPG1BxCgvDWpbQ0yFUwI7
Y1D/438flGbZ3Nr4Stcob66RYwUQ5mDpJDk/LD/JF63MNnTb36QN1F0UELBRMahaJ7GHnk+n1Ryo
Xg0RH00j/E3cnNZDwYElLudW0teqEMB7tIwek2n8wLR1Q6gj0R5qcT/apO9Z7zGljxvid6gIoXJ0
djwhwfXOQkJ7+Cis+vrTVhimJeTNE37CTPN+yxOrTi/KnBeQTdzzk2k71xP2uxO+nIIObSHWi1EL
vQNxOrKF+xBVMz1v3UuK2ALK4QdRGBfARtipzn5dkptaGTGgp5doPlOhgkTL0ZFCfM72b4aRFZbM
BgrM21Iumw0R+pq8/rJ+62JBLSDpJrI3Ec8/kbcTL3lQeBHscLfDB/QNMuZHVDsm/IHJZYYgI8NA
sRgX0leavBE27liMUFYim1WPfqhOUn/8j5N0vtPsFtbh/wpMS/e6SW9x5rgUTQCsTxlALrDH96aF
4HGAiAHBGgEekAdE2Dlkhqs7SMkD8UrA5s4UyOCPm+dpWqdm6GumSD47lXypyn6Fdn8gDLnfpLr2
xV3DrOJHX6gICIb9Fdb/dniMxHOfVpSnddMVzoOBWz3KOF7q9+y4ghMYcCC+4YDgsr3KvKRpNVkE
4uARPXVNptnYGBnLFjl2yUqSpK9suRqkin5sbxNG5jpfk0LYh6huIWo7T/sDtQIcFG6PuowdAorW
nVtJUGw1x10P59wFXWLCb9q+ofsyvvvr6P2JbtFvL5HqU8vArkyo49lBkev+XVCLfIdD9LNHxYXm
tGPqkVG8pDBRxvUO4N/SojCT2Zp0j9YrLTy8ngJACCMP1TtCWllIncFcTH/OtH9ReRiJH35KbIda
OlJeZG3a3Cc5JyoziavZxyNVcqNMMJ8uAGvCa7EuVMHuBwUfy507ZDETT2hzvIW0EdNicmrMtYKL
H4g+9Gtqx0XAeRQaGtushgS1DGBlLbaeH1mqubvUH7D0T+ZHkAobCP5oPnXPCLu4XF3/924IjiHm
5bAnWHVnoQKxvcuEcbC5++nWGZnjhc9uu3rALwqVWj+JhXfQvEPvg1A5GKHvzZKQ/fLbP8US0JH9
yhwFql2pJSUFGfFy8XmAHK56GFap5jEbVi8fXG89GUXauoIk1SS/VITYfCWQkz7caGpVDUZS66kJ
oBiLM4JTCMXlTdV74mcv5GLli/ONm7rHKKZb6AKCT2rjYyE6GnTdkhXcWOZessc8OQ3ZskA/Ks7q
fq9i0VjiSErUXeEkizUAQJL+BsY7iLDp0xD0xOcFCNPxlE5nrSyxd4TjtXGZPB6POaAV/79jvZpp
9bsD5XWHdmz//FQVvObHFVY0W26tIfoMG3LqwBwxYrOzdmkbWwMv5jyOTuZjs4aJWBDHaZrc+kkT
dBo2qwxPajwGuHVfnp8K9O2XAGk+v51+diJrqrkfUgKkULWpS+qcszCmuBYfK6Tn8TUJ4Bv1G6nh
rMRrIsTWCtkE2nTCewUEMjJFQTu74FvOMHMl3neFJGeqfesjuTuD/Yb79fLACjHG3F0crPhgjd6u
S+WVXsJMaLaGiKoDAojrwEH3aCQ0TYjLvHacEhRcZ7v07Khwcteqf9pfPsvgrmbXajKolgdGjrMi
sjZ+IJBZ68+h3OIPg5RBEb8+I5gm4gUaBQ1JVYfdWyj97ytLa403HOp/m474Ck17f+FFQuYpL8R7
mKoGOv0nJDMDwfDxQsvcqQyy+rpQbhSoujfAcX2CYSfb0UYywz2di2vEP4agBExZiWNFGykUo+fE
F+Wo1j/S91YddkANKfCxsUYUMadY0KWbewIyeL+PgiKIh34D/dTC2O+s20JLsnw+LTbhJQF0VOrX
CTZJbeCfCeDvQknHdPVBFEuuqDto6BrDOuHgVwlI/xOIJTz0rO9boiy5O+kT4Iufb50kSymehncC
7NbTBEnhxlZGWywImIpUubkrfg2jiTaCIRGl4kHwITbFJczpSP/IYchKhFR9XlpzbL65X5FR1+RE
AzXhd349QvKGeHv7H1fBzUdwAjx+l4gvJ5x2UgqYEJtX3/qaVH7rjqdaLGa6AWjlB27t949pm0y2
EYK9Z5QCs1lnfE3D35coFrH0+caZCqk9lj0B9Ibl0absCFAjItIITApaDw2w4qEbdu61jW5KO421
jc4tipw95KF09tsABTtTwcqwX2oj04GTfAX03fGPMVxzmfrQbhoH3got6XZ3/9/IMn/babNDWZYc
9xNj4eteZLqAmJULR/YaNk+m1Z2mp8XQtExjvEQC4QCbh5Qv1H1wcUVbsG56rvgtvGoKSm1O+2DT
UXBKvGicpgzHrRtidL93WEN+PRsXBjE+xWrlt1qYN/eBowkDobSP9lbnvXF4988bnPBjFC16KXOH
ZCLy3nm22pB6MJu87ZxOpn5ppRZR8kMHVN+sjVg2HqsamI3QS+VrwsyeEB4S5XUAh0Te9iqLkURn
s6ivYSE2H5+zp3otJORflH63S3ArrqpZCSOkF5rj3joX2X6zcU1QuhKgUzN0FCRgOwl0txs9SrVK
yyrYKjXX5a1naejdpMM9AZaa51u2xBZhZW+R9O8xM0cvHTXL8cVxn02J9IBtzSBu/6W/mRBQCBCX
oeEJamPJtt3WZukKKQ3NZw41JgpDbgh8rz/woOm5LAyEs/LZI/vlCCXqqGmEAoSZ2sn95h/nWQcD
vXrHxCjrjthd6EKZ80oi8cUUHvxoKKLWNBi4EitUXzNtG8CkJlyYoSmB1iwRX9U9Cq3UF4VgyDns
CfT+rTzK02XtHNSQhCLKgQWlKlq0Ce2nWG6GVsb1qxLjZNvf/EA9Yk2eZ067lyjcswX824F3DcrQ
YPk+VYIAQfbi4NPoheE9P98dJT6H+v5T4/kVBShf7pTeWwcQ53zXskVObQ8iHMP1xva44P6ySw4Y
VkfGi4tsplzeAozxNwAOGLsPHpC1lhHSqEXR2qxn/86tMTukecafWyPwM4+vnwHh6ViIgJVwJ0Os
xTI7h1YBDkRvpwn0eGQGNRixupoPMgzMyRa4knJukQCMOMVzdj8w9qRKevzMAR9e75PmftPC+sRI
6W1lKxuGp3zb4I+RqZOmJOVb8gM+DLYjsWD3EIdbnNfzjsIVoCwn6ZldjrHTwbYuESyHcalm8bj/
+/XuzGP8B/Y/cXegSAaIq21uRHm/Lgf2L25yvSWzlj2N8diTxfZ2PJpu8oEXp1LPI32NPk3ewWpw
XOYg+PBD4/6fXYhoI7wVNtABHRJB7YlHbX0Q+p2/cuZLQxD8fPGhJ8iQdMoP6lR3KEmjSgdgKOZb
W3WWDmcz8NiSkr8AbRGirJ2vEm3gRr9XkQO0Lai6hvjlYBWdjUJrtd5H1TYBYwDoeTM+z1eL6dki
aWPkY9lq6PCfX2USNWKGoWi34g9v61XkllkEH2GEb1ARTKmxwhgTqr0FvuSRkIPLla6u9sYn7ItT
DJMgP2yiigNKYvn1jYUF+yTGEidkRCGM/s209xMRRXobD1dQLMGpd0/LUrCMLCfzBly4+fIjlLLA
Squwan7+nSTKtDkWZWMNUI1cWKt7NO3GPh8Wa5ZxAklsao+qj7N/knYfTw9EQdcJdAx8zR+LbnZc
ZBd27KwStZ22VYb36YUbA4x5zrcc7LjsYi8MPDudTmCiqlrvyAo34QzLJiVroXE+MvxqhcD8pF+E
IQMhRKPNHzSnFjdfI6s7nImFQ1T8SLA4cDSQbHKDNcyLsLAmD8xRtP34iDsObvgoK+echic9974x
wEtBEj0w7rIF7XwCJ1IFdtdtx6Dt70J0O0u7pEur3+wJ8zL0MGs58rswburDJP/WdLoGd+kPL6Td
WqGvLOlnIDRgkCy+86kUT0WqY0J+gn108lzT1iZYjnuZx1eNf95RjhU623U547qXQ3146cA/qTiZ
aG7tHHN2c4fHFlDI6gX8wxijke8YH5L8uLqZuqYJ51iFP5raAoOq/zhRJIrWbynyWzQuDBHUBZjx
+F9OxM79oM+xRLGwFa1UG8+vIW62OYzfFIFtnDOEy0+4PUceQBOhINoU+qboFgjFBjGGTmPdZ6/K
lijJ42+YYcR8SDi5b8eZ8S9DBSXkkMlLRV9Gr+DlVZlHOAgJlk6xjCURr9mc7o3Wo/URBnv0fBZ6
IecnwTo9V9HfBwCMyXVPlNlVfyhBtiNn5yRVnSHyGHpL/Z27b6AV3tsbRKZZQeoR6rMaeD2CGKeX
TNkSNVYHa2fMEIxm47QJEUL1WEO0iwtOSlLhWax3h6z1SOgb7VfNL76xraf9/5aAk91jVOW6aNj1
O++MHEPrVO79HGiMuZS2XRJ7+oWAQpS1DQvdUz5yYV0f7XSFSCG+bmyYFgNE+lHoHH7holPQS6iu
GqFCotWVQJVMTM9Ikr6nAVMXX3ndbE5YDlz8ruqQ05UHVNxhc4pqmbLM1RQsZrChY46C1QNPXBFH
CVFQXrY6sNLNO2RImCWgdqkzevvNetKLiabbVHkqpd5wUkgD9CfCbFVZ7nB+DKUmS4bufAUytHJc
l/3OYZGdD2yZL9lAK5fSb/TgfVySblivXOQMnPPquU2FA65yM+aitCPw4gJsb1PqtTwb8cpb9rFp
AcWekvVMW2epoB+8HcHe7sTl5MylzNPfOloy1U+tqj6CPAK8zrTK/k/KXKa07sGPfLcfUA+FQgpn
QY5aDWdIpD36O0imV3XyTmgNz/nSpgl0Qkx4b7C6+mHYQwoYoJxmEe1DfgHHvdiLvMur0KhqPI+S
F/1q7AIX/szWNsVHqUs8+nM2yiP5P+Fu8jZ0vRZ91yQB8sekvaWmkl/kzPcVY4apuU73tJb+c2pd
O/cCLr0S4JYpaf8+Lcu1qpCRhvuqtJJHJ4JpYd8Buv4YalmD1YSgJh434b0rRMBFhyX296zAIM2W
IPfcg4EocQOMJVsfWO2K0ZSLCDy8oaDmx5dtMq2ruUW4NQVqvcKSb5Nbz+hNx97cuuMUU06nJBUw
Ox7ut2Zd4UPkFjwhcw+ifjgCBiDt4U+BYYJOCZc9qf9E972ihbYCp8deoKQi+6o+hGu3NFlNxxkg
Fp6684cr17nrMKCaHzOZnhtlWygk2Rp61SdRJMMZgkN00+Tx9uJUW76iQVHhIp/GziA2dgy1DH5W
geHuiBbSX5EmbUHch0IYy9/y+guJZRee46TKhVvKfLqm+qcNi6p1aJSoIDiDvMRKqTL5XycMZbJg
HaJBIEwQSTBK+CSCKHB6eKnFSP0qpdTeGwLCQ5VyNGNc9za5QVMJAtonQZfAsJW9bajiklmrZAkt
u7VuLA1+aTogBkK+e3oUBLbKQ3LwyZiTbdL6RDGqZ+1n1eFtxnHIcu5Xae/s/+jO0B+pyKEQ7tVY
lBVLDlBSlMWXiJ7j3TbbT58yjJNT9i/NRhz0RuodvPC3yPenmo+o5XTT9tjQJqbY0ef1viW0EuSL
x7+1m5vSfvAcND6wQcSwwCxNbufCi+aG00+I4qvKWkUON2iMOK5soEFcD4YpTZ5MVtc5Gh0Nj2i2
KwCV0Ql9jhGzYLVFqIeMKZPq49OEOle+33miIMXNKBewwTWduwyhtLtK3Yb4nsWNhawCz5wj+vzV
YS4DQxDqNbSWYNahh+UjDaeCVxIGq9iFLzI+tT83hQVSAlvOu/T/aOZmEV2AmWzk4qiakHq29jXS
/OFJFJplLrnM6GzHbJh+EkW+62+U5qWXk0KuaIXoyO6IBpB0NQAeTSHDsB+upWkhpaCbznirDB+b
SGYuTxRXraVHzcog6h+P7kD6bVdFFwKBaW6ciRTHhElhXfvO3wc726qTzv2mBcKWnwTBvb/MD7OP
KVNhE1bu40eGJ2o40E30eRWVkHp7cpS122HRaGJ1Ytv7KZuG2/kyOxW5gJ044Q5orxjB3GNN5zIF
NazvY7eZui/yOzgGa0CG8p23nUAiskAXwsV+3aoxDrGjrQBgHIzGpv2ABHwthcCrBXudU24fMxcG
BKLBQNVXOiORT2ElrhWdqT75SU5zCFGF6qwjF27jVLJKYZ19GSUtO5M1rGCehsaei8HrGnnZTTK8
VkT7bpc0G1yYxtvIvO1tyuEErPH3maiNdzY69BmvD/r2OczEM5boJ8YsRkTHEoyRWo/efO+ArI+T
pBMYqJpEsqWo7wAHjJ3cpDhL02BVN2o5D3SPsF9s8qWApKQIo/rxv9pFrDMDNA8YKuhdvkcdZtEF
KYfMYX8GnhUTu3KSgaNsTMzN8X9HsQqXGvlTwlN4MSgKCdY/axFa8JWAHFK+ygBsgJTi2QlW5jaV
K5nonzN/HyGTufY/M+IG1W8tcvUEBupyfEW44T/gnM3rmAnlZV39e+wF0fzx6Gq98fqcqhe1WMyB
JEkW7B82+/7tb30Pm/HzokWkUTUaAEyHSryfBPNhqxPWTbfeQ6Fqii/KmoNCH1TrewZ4OmmDPWdS
70fePfm8HVjB980Ek/u+oPPjthI0wLPWSO6RcoJZwIgF0Af4h8HL2LCgdu9DYPwyjWlHZM4qQ+xt
6Tdmnf3SL6KFDYNG0j8ZS+63NlNK10OPvp5y8xhY7JR61tJh2zjPr4kZ0oXDE7MjFPI4t9/tIJas
O+fLyrgabQF+s6iyVm3VyOPngxYVS/V/pfU4egx8jywtg3XPBIMPIT/8ZjskLZXiz46f1HBK1uwH
EOqeTtEzOWEL7VVWWTCHALmUceXQxdG7TgXZ50jFEQPFWnmnwRsgIMOsCbld4LPDSV5x9JPCx9qP
9x1w9GaBxdfTklk3CXARxocG8uzutqbzhdRuoXDElGAUNlsp7fq/P8v9uhnEUvQJaxwdCtna3Zu8
huDvipcrEHaP7RNYsQUZSbex1nfzlIUEwVnvl4YwFF2ufyCUnK3YOyg4il7z1gebiHcWWAp5J+Ie
UW1BSCieMWCbnep0OkEeP682zOegf7zvbq8VHfpXS0NhqsQNIudJzJsf1qHSd+Q8jZ384jTb8bSp
YMdT5ivCN8hSL5M1iU5eUWFro8ha7hv26GPNi05uJSRsus2UVskDrOPrmnqPxOx2cw+Ajn3prdha
BJgbEQKbf1ahPId9DyBDHxF8x/hr4opqWFjCMaA57br5giIPPupcIN6QgMfPh/HiiO6mYJO11meX
bgQSVa4gndkv72YCuN46t6plbONqZF19F87oTfr1G3LokpgJP1E6U7+6+aWZOKDT0KBW+daHCwcq
fbowG/9tsavQUUvzTWmK2lZjexzs1GgXoyIht8zCXxT8twAg0mpJ1rI5hku00xOTy8ns7wrYQpFV
63i3tk+3KEMSHnT04tnedun/F9bTN5etUx0LIvzoEEOpgbotU73XMSYaG15KWX5+x9tzH5xC9eRR
obSsKjT4E+MoOBM+IK/H871m79d9FZlJ17S2b9KIW7Vgr7QnOUA3ON8MlSOPEOxjtV5HLDYrEsNR
MI5ZBDdQzyIh+h+ACGQXMQJKNQLPcedfwOR+yZ2fDVznXxVdc4+TeGe/vJduW2r93AQbDiV6WG3L
Su7q44tywZGWqCippTwKHlLAfVPy7xbyo3Ig8fYbVDDXOhKo42KiO175Oq/Vtc+WkwAPYjbS6J6Y
osQs1krhAehEbPnMZALlUIRJsolViiCyLaFrZWa+8NaFgFHP0QqW+UjMoBS49lEUrMmRFoo41nA2
2ptsB8XjZSIxxGwn1iJGEWsgra4IiH2PIc0XPDW86KQZVVVLvF94Hx8H0kdQRa7UN96FxtE3w1rG
6WFKb/wEXF/j1Gl71ml3gQ0vQEws9nefTN6q9tLixCzJBSkOQq92VJs68ANdtuB93pf8MY1g1k32
nu4/7lU7ULQ9wwY6R1UF8EhGbJ6Xd/JlXYePI32l8yi3nwh0kBBvjT5KlBG65qNOaMxH2CKUntTG
nkkg144cMe+zQIWXcBvYD5fZXTAmQFXIqJfPONyY1oFUQz0l+rYTggGdEVwY+Dp+aDMDKFC6SqjJ
XQvEv2fvzK1uF8p+q3kb4dP84KSiZ/K7eD5NmWiHUenH8PboHdyEzsBqC52ww7ViTBlSC/6u78Hd
gaOWe+Z//0UY8q9K7zKAYWJV7apYlL1W+YorEI/6l/pHSJKqt5wU7aS6yOv3TKikfv2t+YhMVVfD
7xyuOz1fhAjsiuc04LFVrRuqyJUSoJYhBvwJkzgliPT9gjq3uDYbAqZ+wUnKP8sTyyheFVVwfgmR
7hIl3wQ28/w/8EMF7+EnWzYXXLP/mj+bcICfPKa/ckakdvVT+4WU/gvhqLRDmMZPM9mTWIEXLGYl
KrWAgN37Cj1zCK4v/g9qE+YSqR8TfOjRzXpKDLuTYtwFpkx/14nsl69qsA5/0urg05GRj4TcpAIt
FRByDyJDj5H/A/S/Nul853cvrWoYK6kDTCSYb1kJF9R4N4j3vEtTrXMm4P/sCdgRSc/MK2ebnAhw
9lXZr8Ul1BkUlR7lDEv0NQT6RVbJuH8tfW7t+fQmVqITSTqc4+fsSy4H0Aq4atOANXfETO79nDqp
AMrlGsY5uKKawxNQ7F++yVXnni9wWF3GuKJieWI3gfRoKSuix+738CJsbu6ObALLaKL3gTVo9Ndf
x77X3RNCHaMER0JAyALU8yLAa151diWtiL8pwSkE29nN+WXkdXYOYaHgva076EkXSyaO7zyAOZgo
lro0z6Hu7Tr+zxcEuANHgQXl1dpCOqkPpC4CT+Zvhm3RFPrNSU5fRzW3/GMjYLPW2Fi4qfMr2/Dy
fM5dU7G8VfYHmI6UrU+wBLYLzyeYIeqIO077PU9ymy8Metl+vxQRoTIIy0+QWB+CLuG+1i+x/2lX
bIYyIV9s/HV72E07gQInW4ryuc2S0dgNwRI0nivIfxtWZzixELTIIwCrUewoLNiicBpkDTCdaRDQ
hraXqQ+eKAOszq4yBDRLQDXQ6fScx/X27eF7u1yw6CXyZo6k7wuMJ8/epO8AHpE19aA3qb8Qw4De
J7njG1hzZK7bIDlvrRPjSWrl0+3BgvjFgQ/xQSNeJgiLtJ8uXGMelKIlJOVmksqk25TU5CEOfsEV
kvhOYaMLQoP9yrO07YxZM/ZHWpmV9jDipwNpCv2nuwRzU4vcSiChD0vN4SPaYkWNG/Yoz6jKD3+W
JjfF1ghMgtcMVdI8IDVLgAcFS/p1qbgea4+2qtdjySdjmuQxfIONQEG6k+hh9+xgzJZUTZjRwiSu
Yac4IrlPdfexTOe4N1WQ4guQNm/YFF+r/oDQkB+S5eBnN6PaZNgyd2FMQ2WJF+7XWBsfpnf+aYHJ
O06QQyJdlJ/+GOBmc5m0gZH7+RzJu7a9msaHFhbVKq2rqvteJuMMe8MC+/VFLSx80/z2bNoesQbX
OJjrwRZk/iDR9oZXArYiAdZqE1neKH02Sb27JySq3vODzWB4cAfJZ3srJnH+chwg1D0LTm61j9ou
Sd8XE3TS+ueWwf3rI78MgybPzb+8az09zffP3Jl0AYmaebNh7qr9A8oddEsOGkBYPH2JnmP6Ng7/
oqjteUFVgn8FP4pXWImv6Lq6kdLzyFR82yH0qau0caCg9WmP+uXe9vd3S2MQS15tEqQTxyOhau5Y
JlcClASTR7dx9d1yidWr2p/ArA8+8j1sSAYrsIEfshi29atphMYedVJwQxQFusolHoca4e0g6kJA
+I+5yjqkhRLHxd71ARm2a9K1fo6xHYn6g37ji5RvqGBH/mmb2MNZIqq6IzdtCqYvxRcivhE6wlrt
QDjpi5z+UIqUY/WGfv/ObzZnNzfMG0e43uhd/a0S5ujZERCfYD4xkq13odoVVlQAvvKHVNlAM62i
AE7kDkgL2glN0EgZPLkIsuQYB/3rOPoDnqe62nddVlzACCy1ZzSBgXSJbklhGNESpYmVCzb2/x3c
3ZIauK50SLIF4DIw4PF91TW58iz5oLG+JlvyVyzwVISv0KliOP9lT1S5GWg+CohkIP/LeeFGd1nB
KKU6bdLL9cctIeAhs0KZw4n8HtLwIVJw+y8oXQU/FL0YJaC7H5ZYqktIyTF2abTkGi7bM28SNrGZ
4zBGhqIMlxdFeWZ5o+mRirOtSwEuPtTJcoeNO4YtS5dfGE95YaIIQQJlZsJ1m5rrtJhLWLoxggyb
4cla5XHFTegCByIJ5U3KClR0ZCR/oIo3t1pQpZRgO28aBwJ/omNLrvK4AtXsQkoFgGU1LB7rff3R
nvnd1ODYeegy+l4I2SUV0kdfo3Vr4s8LgOKWuvgveEWP/nrhujs39LFsZZgkW/bLJZD7NtoCddwY
zR72wHxQ4tpKcvtfoArPFqJi30OJQnKN6ypvicKg2IYzy/PelgKmYnlw3bAYMQ0/WhBJPxyR5GkP
uEo593VNWJ0WTMKYPbvSh9bS7BEnRzjuDQj2ec/btmbRdK1yNd7KHELXQAAWKwWvNwUylIB2uOIR
cPgJWUZ/LGVXpPfnZaxgxutprmi3Ouqi7YGptPsP1r+kNaEWjUTxKFpmEoefyml0o3jEp5wdd1PQ
Ro5zvV+aSHvX/Pht/bDIXWYIQtwW72U/0Tf4l76VKIoHtoPkAHPKIqHk2HJbtk1/V3drJ3BTObNU
G8T0zEkGiHuQ9EmJE/fev3rse8G33SGFooKz+GkzhlkNJnglG6sJXG3glx2akS2RJIWGN6eJ+Rn0
M1JMf8EJXqXPerhPdA5vZMv6pszHkVsBblh7bYBE9GeUPLVfYEVfT4kaIjzK0gbVEB/iR4GqunAM
ragZjt4Im+gpdBcVlLBnPqXJAahtK58Kj4ZOMHvSKAOUMdV6sEs0MfAD6oITdIWwQkpPKwY3hOUr
DSCTESZrewhKT0ugIIhbr+JxcJZum9mlRwSnZ9fPof3zemZNNYIaqW+qQ6AcBJTH6wLpslXDC3Ue
78FpAR41arb6kbg/pQ7+NxkJsUVf+HAM8b79d3XRnUk79iFBFz6ENH7/PtVpeeCDJ97o6cknJlg/
DViKUTp4iHEoHGN9pqz1zVYHqZOsQDtl0QOmluG0iO+uBav0w8Dk9ax5T6kXxFnMNRc/rjKQwpQG
olQ+Z/WVsw1xjYIuJsFEmIOBJnMXmwLXfNUMimT75nFgL0wo377yC166ahlI9WFSiG6hvH3X8FJ/
WLtQ43fBdx0DsleAeZg0ohH0NJEOnlzPslC3y9AdlORSnpaEy2Py0kJCiQze7jxQ/TT06seXgMWe
dqFlZXfelA8h+psujFx5Ku6qGGs/naCrpuBam5mIHzl1BfsNMzttNL6mSw8FDnIJLKFuSrl9X4II
hJRof9b9Xv1AuuV61kHbAoWEZn41pPkkD6BZQkh8xzJHZRGk4VFZg/8zPrPhgQcmzEuCryyRXimh
K1ypoNE6bPXzKSGWx3cRzFfb7a1zRLudY1dLU7+vkyd0x0zV/FlrtMA9n9XXG4SBLHBD4JXwnz9x
rNYANrtjtPPQXRZ9dOiQAVW87RJYfzmgvenoJP6EsJurARhhH9mhlhR3QUyJ9/RdlUEAxZc7Qukg
ce7kFAorUQSXCXngOqYY4fF0RgTIH/iAmnMfGZyVxpMqLgHtt0yjXEJB0rp7Zn0kvB1cUBIeD1r7
c09dBAtgPymWreJzvqyFVONxJdzL7NanJx0k36SmVVhA6R5quzZXQFW7mfU9fyqd/JONdgGvm/up
ISVuWenB6FOvFL5hvIsYPwFNTXRMHAfu+J4u0V2lvejbtML/uZpMKWG6KAY098B8nNKcXhil5pmR
SaEK7JERzS37uWtuacDAA0wFpcP5B1Xm8u+XYpxzXYccvUpQ33By2qfCOxaeiVBSGLbBrpGn5XVF
hEpMLrHn5ZZz6wG3YYvuAhZ7g/uY0sJtEkoeiTgD+vW4ZZ9IlA+mzd64IThQkNw5UhQS2zfu4c6Y
DCrDfvn/h1QaYBYxth1B+Ni9T96J9zPPrPNSMxbSl6y5XT8J7ApjLzqQUq5G83SGpHZqNQclwRM6
36DlV1fex4AEpx1Evrka5K4sdLgdcsPwnU5v5Tx7GdchSnPqtYTmXXV7ti4XEzDu681Bt/uAmpU7
IL/JK2IXqUJiRucxeCBpoh9HHL3veoXtfTHQnRnmPb46ubzVyk3mNW0PqIfDAicH2ztHbn0pb/ti
/Oa7VQZydRyNhjqVb5dF1WqA2GrgUzrfLuxBZbOZOUvPZhZhj0UUcEwctkF5rLryhTXYx8wqTCu0
iT43P371IkTJNW+OdiWFv9pPmexsJn+mKsqq1quPrnMqW37rmvqrR0yPghPGMESBT9vdM+4JTrEl
h+VsazYsJRnNuetksonoqT3jb+bcBUUDTiYlp22esB5IHdaNDOIAc0uSv8+ydIWMm36ZUpiT2QOf
TQT1VGK8iq2VcHvxt+Jd5YVzTAPRtgub1M6JkdBjhvY5PIc8KjJ67Fe61HVD8uCDe/bqwBKozPL9
IZI2UQ5m7ZQ8LqsG9rNoyJj452mV6ClvQBsnpI6LHK8hURF3AnkaNP6y0yYN02ApK2PIuqi9/hWy
n3R3Xznei6y9BJojI1UAatY4ySh0OQbng0CXTKxJoGYAOA8THhS1KdVrlxIvIdlMdi6PMmIZfRl1
t6WEjOt3H8ci0X0XBWOt29oPHmv6fgTnD4799qtn9PtHRfig4RlZAzZZe4VcHXkta3aIAWu+N4sA
8Bm13qx1OqhuchHiizAJL/Psv2OV0Q7+puS4EkDNjdK4dnwNH0n6TQNb7NgKxsBq0QO4U8YO6mWV
e8SH7+qZ/OR2Tspg8OUSLBwAsg0B2b7OcEwK20iGeapf7t/qWD8aUrVF5aClAqZZzPc7PxFfqk+8
G8Fl+UcicTLWj7jDb3N41ut4Kfe8MbUJ7j9YXn4FBZFxkgD9dpZCPQBWumKyARIwoTpraU/8p/VX
gNppG337iUazMlVpSc+H04Tysw7H0HzFjtl/E0GPMrBcms8lMSPiVBRlr0lwzNLF3HFcrxTOYJTr
N/kXLLly0279Jj2JBT+Lb/AA8Las3QR/jJ3hdw9pVRqpAszs1q1/1lZlBb5HxZ+8L2VwpqCHhKjg
IADGm2aVevATHk3azbNwSSpZUqHFw1yyBPjlxNWXa46d+s2C34JYSmkM+1Rjwe5p2v9Zjtl9Wd5D
iCRyNOT1T/GCTFLCPpbA5z9gR3I2d/mOeq65D/PoNYzTAZ6Mrnsd0q7AkSiwyoaiA6ygzQjN/HWV
MoyYgs8+5q97gyjNgdx9i6CL7n/6WhreGy/Qfm/EAjg3P/VSAdLtkwy+hFRskPKazIIILgHSvRLC
a27m/iMdnm8YrC98wJ8XNkXtP431M4c97wj9f3CYVvesZLRzVYUyJoq2z+QjpkRTlYrP+74ahP6l
pL1f2JtPIepUddnm9hw9R84nwCPltHayuaiX69qu+Ubbr2YV3sIqrb8tmcIhHkTrTIRiGNQFsx/4
yIs1UPvK0tuWsUI+GnDaWJTam6PVeQrM43oOEQj9px+ZCZuiWgCLRRK9CS10Pr4AHCYLRBlIkOkD
j9weabAL1Tp9pwNr+oI0/MfdvNZmZ/nBiv6otkEzYUc0l9PUEIkYRmR+tRVWXQuw33azWhM9jp/y
Bo1QMZAjGxQ99HF6VOFAlt6JDVEun5gamJNJmDwiD/HleBho62n3hNSyIo9LJdrPPz8h6CDGXOBT
ivWJ+ShYmdzBNQKSBakREs3NgteckL7dObT1NB/lg10bY3ng6KbPeB6NQ6hohq3w59PB8bLbg+TZ
V5JFMRGwl+L2SYlHGroqbB6dOAPUwQ85XLi1kpl73QdPTc7T3EgFjXS2+1P47yH3S5ryT2llC6GU
okm/D89sdHje68U/nwQgND3plXiD3i+XjVCtucpNsqHQAtgUg+og4UY5l7SGhN02HW+CLV6uHGjk
J8v9O8UCZ8s/EZ+3xpDF48V9LR0jN7qyAnpYcPFRvpdaLDVrDyq8hqC+MyS9XdpvVYUBLdtHw6hk
GWaHuUs1rxKs92h6b2wCsUwQ/2NCVtZwRHYlyp6ptVqxQn9BHXsMiaVF9MMn2rr9jHCE67JWmF58
wp+0KHhT+Ycf09wCQLPQLZk6kJNjNiM6jSOobMJj0ICOnPbTKvgeP2TupPKeSbb7DMErm32ndIS4
BOGw1xNJcI9Itq0EyX5WH6CEKph1yj6BRd/zZE40BeJbJ8LiKhTDqi6YJcICGfV93qr1nWDPVfRR
Ug7Hh+Wz7gdCx2wd0qLYeT5yWyjlh/xzz0fu3+Ek3BgiHS5tsoeT8GyLPBSTeXN3ZkPF00dW907D
oJonCX9uc9hJj7+/bOQaa0chaIeXu2FjXZkdiV5Adi6ZNcnmmVIA+SLT65tFnzmfAhpArF1Ebb0H
MOUhh3ewBgxu+nVKosWdBAc8LItzk5zvH6jNhXpLRmhRotMt1ZX5Hi9qSTfBiQjmK5FHlaNyvPhj
rDinVoFQfE8E6d+VrVe0uTF7GiFrH9WToTFDHAUEJR4EZqocFW8zX64jkTAYQ5tL3r0entlotnaL
dK22FzOPAEz2FVI8gf+m2jU2rdH7Wzb2oyVTnFbRu1+5DuU0teYxnn9Em/KVGRI6dtdrmh2J3xEd
XYfNOXpbWdUt+mVVuyQ1zBqlUJYiTni08E17SxC1W6FX1kLsVpFjCmbsYHI+LbA1OsRDnModSA9W
xERrRmb+75XJzxw3ttkEc0fuLlBK+r/HQN/5Ly1Ux2LDHplgTauC6P+UFaWQL29da/iiYmVme5eW
Bh50aQuZmLPxLgq4XnBq6JVP6oaQss1cJkz6yaglWcrI58nLPuFcQ69itAEBdN91mezi+VsBBv4E
cKMVfLlifmUsBGpgw+cfjPGANg9iE1DFQ5U9un/BFeSMvxRnVl3fyvyRog+E4H+FwzejLqKUsvlp
pRd3lD/qKV45klCwqv68KDXvKPkm55t/S6WDcfO2UskaHR3VK3uD0vHNz1h3uvSVTCJIInj4Pu6l
sXNMKk0YOmQx3oDaicWe4BRpdEv3xl5j6DzUZRKad6P6sHhFPGzF05k/pISMLRJZCTTieBdwJwTL
TBHwyBXoFWvBbU01MopdrJS84yzT+giAVfVeM1WLydZKnizNKTpFWpIu3GnzS10hnGZQXJ09oV+A
taTwEdW7KaokRskOJLLnKiEtaZVUBeHRuZjzZRuguqqI9K2YjWRxSMi5WyKW2BTAgg0A3yYpTtGk
K3bBmrCg/j0QWWdexLdLV5cwgBYPeQWqt0jMYGIGQ+BC4DBrIPA6mX1EWZSWGIvVCy1SvE85qW6N
lCCfcbQrMOSvrJtyaRnFT8AwjbLHSMPdFaT1PxiiUXsQk9wMyfHL3U0rCMOGkIP+BJFd/683ocvg
xpeW777YpZZ+xpZK6YLMHlYbdoj1HancQCiJI+5cwiaTsFnneaY5uS7HoNkfgO6AeV3AWSSuvFs7
81uUGmDhBOdv5t9pPgW4J8x7YNP+oB4G4PCQKUiytrhVUpMEFEHlr3m42AvH+Xounp0eyKFH5GgC
pb6qHHunJD42wkxQoMS6bpg/30XCtFV1DJ3jrpg5e0pOrHXEfHMLi/IiKsIk8OvqV9jHDTQZY4v6
aD/w2hCZmlqY/vuDtVlO9AnhttgjHnOCravFTKTCbvZGyEst42PyDLmv22TP7C+hl9wqzYRp460g
VfgrgNd7ib2U3V50KlXpt5GespuNRXRugeS002nC1LCQFPc0QFlaV1Z7OCRiAhSwB2f6D7zGpIMn
j4VlB8TpgGRLrmlzbni6V9Sa3tHvhOvNIiznXPe5PxobAfiorYvJI0ffG5wmD70/zDcy5kscDi1v
HSv6BsNQfiWBJE4hwA9S7yvq+QHWcGFXu0Lm+bSSfbc2zok9JKMpcXQP2pDv5cuYlamv5rwztF+9
u64idQuNv1WozfE/ePeL7UjdMKMx9GzjsDE9gUXNdIiZQp2W0FJ8kE+TXEbztG+F5uv5gojs4YTL
oR2ROEopn1xKbKswTIZWeEmeFRW9EWJ25BFjiUzMjVCZgJ1Q2kUTlSYt8WHNtBIGbWqQ5l9jMfDo
Ow+NS5Oml2S7HgRjzBR3PMFvyVuSZaSJ9fLXI5Vz7fjsylhxkc9sb/HzxG0Yz1yxjHsaxxc8enLL
qHml/0lmHiuFf9AQl3vcCxO05PcOGufljiBTUmQw1GWMfW3B41jtIYq6mGwtmx1JWBwPtRJXuBKM
I0X+hDTworfNm1ELFuwlw51Yd+UiVwC5JmoFqb/c6L99douj68eGnnGLyT486N6QL65eiyM2bTcN
A+x2FfRj45xNiqArsq0dAPdvLQz7N4lhXpcaL7JBFedqW5HI8IM2fRKjP2kxjk8Pj18MylyRONet
Pllm7q6qg2njGcErp6Yo9r8COkuMTjDa6E0v/QrPaCt6TptAxgalxZFq48uo0pi/NWhwM7/1bA/f
DS6jS3UfY8zYxb4ouF8dt3NOmg0nVnu8v2iSHm6Nu/7gZzQk5Uxi84D3rKkAg1Rq20YzxJqlz1H1
uAZLGuboVrchJQE62Dc2nRHbJWY2Os7extAL9918DrF79dWjrCFtavi1LohgBY9EmJkFXAPBoP6w
tkFXBHVn/E7CM/zwuCD39DUtGe9nzJLrMPbdzhHe4Asfd9iSbZx7RQSHg0nJGwFNg5GERgyfUGc8
F/1yVoj046mZMGEwzsb9kRi3Jj+FUAShzyAPugPXpkpacFseQcdprJbTc+aRpuHcgDOzNQbPgpkS
ukGdBM1F/HoRNnuZvyVrW6Ux0BnKVE15lyqokkoltgUZuqb+Y1c494mqQuvkUOQ/pyDumkXpUSW0
EplK3IszVxtvzRNszH+QZ74h9gT9wiayDfjb2I20A6ezcWKyil1pf5i9ej5Nk1LMipHPCqFI2guD
Y39A0o3Ls86tAEqQXFPsoFvRJAPPU+C/YyGVarxhBJvqjrDlgQRNooRCWf3Et9W0UgCrzpFkcJyJ
+4G3UM04kUn/GXC69Xtc6cr5wYWZrjeJmrOrGL732Xi/Jeztwrioih7gIdN372cKQ64LB4lagqqP
QxXiIOvpt/ntRPP8wyItQu69MzoQdIdualDayY6QvuiQ4Yf4XhkmTLRSMjxhQXmzPGqhs/FZEOII
88raruB+5Cc40OriJEEHFJO2nUwSI7YE0vfOemuSS3X7+bnhK8Eu3V+Qya/uQ54WpT8bUbuX8bG7
sYPT3zsLB2Or1eSo1d/U2MAPEL7HdE+JShH+A6wH56QYHJrTwjH+lc/QR22/79E5ga35UYOiNwkk
GYwGTRlpAxkD/bvVL4WZm/A0Izf4B0pdTUzddoQGUiiSxQqqKU0lOqNWkMOPW1zhnIlaF1UQ/Fzl
ol7cXUHEleiqpC/SR9DmZ3qp/TcKHMC5OWmJ66eex6aeqXzvE30qnZ1NoM49hvieQrdKwdE9DG7s
Iz+sW9CHCgPyK3SNMoTvo6tCrVbPEScBFm/pGhjUOKoguDkQjHLNngYyK39mR/bLv77bpWAoN6D6
MHdXQnfAfbKLbNiyZZW7H+xw/a7dtu0SEbiSOR6ZNrqzeYDSykxs8tp+3x/Wu43kdToe57I3SnYM
gqOxy6siXNZfvItu/KRuVoj2ZwKpHTwN+OHZpE9xxojZu7dqR7CN4V04h2KNKbwXUi0vF14pMA9J
Zrx53ZVjnkDgQGN98eZaaSMZyq8sBOCdfWiVOwg3cbFXMjVOw+Rm4qIERz0oqWTlqqZsc7dsJCTN
bV0lgGJCTt9mPTcysUvukKMeCwITqIFEOKNriGYBc/nCBCPfOCzWZPbdTlYgKyO7KjbQLjCHy3iU
+WhQeHrkSa6MnyWtmOztElmOgvLHUUU/xNBOR3z7BdtXhyRlvC8+Q0utkWM7G1KyWOjkrRZTI21z
9F7/DyZK+8Ecn6XJqsRSVIXE661KHxxZy2BEhchKRsBk1qnYwwCPOK13jj6JEkN57YGENxL99ZxO
gnW0CqRbf+KzLOw3UUhh0KPhPVYU71BMiYYERWPKsG6CPjz3LK2oi9sjUcD0XU828UPGNecywa/r
3hLCJeWlbKNfjHwqhMJczb6kdFq34YZ86gOI9zuuaZVqlYFaFm1mWdfyPsf3zleODaRbiTwAx+9c
fGo+6xUnXN+Q/HruyWC8Swi4ewpuIyCRGqSmdrMx6ZGFXFdTTQ8gtEz0Xgi4U3YTddFWbxnGPRc/
JofVWJEcBA1v+WBcNkaLBxBExAoTvHZPXrKNc4UMTKAm1I1ZOqxJij0KSiQetbSKlXF2Ae4DTHLW
4xHYzsA22ozFVockfa8ym3b92zPN0NwPZahRoJ+Cp1uctpH2fmhRf8iVTENAYx5dLw/7TOFUHRNq
BaD+JTR/0df03hTTbnEPMk/SBUMGsV+awUPpAUPwPHwaQ0v64ttF1IPGKKOhNRTL5Ujx6CoSVAGJ
rTaYJCz6iVRVWcjnlSvP3sV1XhVrnhOafwwmX/qTQv2upAulcQdVIwLZt2kG2hidN+i7l74XufQK
2d89+qHkRqqmr6Jik1+eYfjW9fsLBWywTTOUteULtRl5+2y0ZSp3C+TfTTMdUDACwAgzy2otze0P
Q5IfStJ7G62fDpbufXC0V8nUrE+3x3SoDMLoT8GbvqKp7CL2O3/CkW3vytbKefQtL5AUTD12Eopt
Q+ZynOJHtAD039IvmlT/QR4d9oCVjpsA4Ird+KlLkb5MWpXvDIQTZIGg71ftEW8F8odrGeqzHhxs
jEgCtwsye0QHlotisL/Ut/26vwkATJKBuG0DEMGEW9JR7sHExFlIjXNC69IjnmcUwrBqarMKZ1yu
r2JeiJ7/hEkdkD39zIeKi4QaGX8Cbi/lyUZv/7t98a9BxWOVE2+gn03qahC+N5Qqr/NU6NoIyjYY
dSgDM4vZcHCFVK9Js9EoPC/WukMN17I6c8UDFGbJfoqOy1xZomDMu9MvN1VZZttnVSnH9kBhW0Hi
XxfePpMaerPtbUil/o0e4o4bPgFpXlAc9B0mfX6bzmr9fRBImMtauBMUkRT88ZJDnVNbE+2kZFRe
Np9vXxJ3fj+xv/cavkOUkycDGWuJHH/olV1NyXL3ZEJIHPg4MWfzoALb9V4zpJl/9wV3H5TN1QyL
dJARSiI9pYj8+2GTspDHfD23obevsbgb2jzDVYYSBRzBVchCy3jPI00nEd353qwG9VIzTeB2WGTz
ain4Trpz8YWtnwsKizWbUIERznCOHgQJsR1IsDyAcJZqD855FE9N+z8o3k7EP3x5IMcEGxSD8mjK
u/FoHtAmzZSq9Ml+bXYnsWwy+7XrQ7zs2LXJ+kucbEsN5PAfRddxYZ+XE7BkxhFkXvxO96VcpwSf
HuSkWJlZyw7FLQaFyyPkz2xIDj6VDoKARAc+J5BarNAjlnDDbZrX+bSKs+vhmRLPSDVrhATpX313
vZM2+X36trUwhlh/oSAkX1FU9XwkJ0T7SusS7WUkuPk4ORPmHub1O9bfAzNv/M4XsAkh4SOB2l6l
Dhp5apodEU2V+ISkj3D7EvBrYslFr5GPOBOD4N3HEdfC+Y15woXdU7dc7RF6IXl1wrSySXIgUlY5
nxdnKC4SKMo0fBU+aQ3Axerqc+Z9NBLKWqLa8wysIvaGDhuujVWNUVm2yBM/7CmjLKXi+TrLg05D
EWq0VI/6/MAM8ICFtAjuau+jSHgEgqowMWL56I2fvcls4hAxv+DyT7uUbTYsfPKTwA0HUonNXNEn
Vi9fZgZ6sFIuvZJugjCGh9+p3y/ouRy6HTiI0qvnDbcoKUCjGPZo26HglgYIy4XF2w7uLRBt7OQv
q5eIAKaE3LhG1LhTG5IyIltm0IT4ahUKjULRiWxv9o6jueK4bbBLNX3VQX8PpKRMcGFcopNuKFoo
XGFCRzT34fvRtp9eMUE3bVqRGno4Sx76VH4uIj7JOq2R+03w/556asHDJ2eKjaj2DEAj7eg4aA+c
nVg5SchblJARhNnh3MuFOpGQxi45UyAFuvj10ohVIXL4Tv+due+xd9jvg9Gn9ArdIqDTgcyt5oI0
oB/MTZ1xih9hqBB/BRYyLXncqkbBqYuXHVHwYlOULF46BA/3me/eAlYMN+VgJNhWa4B0/9TT9EHX
ZUht8FAb+zTfl+19xRGjBJKrCcgDNHhDEEJGouCdJEKRH5ARNPAsY2Kl+No94vRwEQ4kRF5QSOUb
j3aCzdYqG++biYBKDoA8ymcr9cAdTb5TCo9s1Oi9P+xmLFtAmGDzkO+YOEFV9EgmqhGNdlhf1FTs
3uOiH1k0N39P/8VmY0oIQ1N/AovnBfMogkRd093h7bO78L6xpUP5uwsjkQgFvME9YGgusbTwFvYv
WP2asPzCb44ab8h1ZJG0K/QE8bhh1t7a6eh9QncTOR99hd+fCS5Mtkew132bhZ1rFijq2VsxIMOU
qGaa+NZx2o8BhYvGHUd7Q8KyN/lKlny6h3VmvRcDbC5aeiuKPDLHiVDQSiwNXEY9XHhActxb8o5o
zM/YVIMmx8gtgBofVSnCIj/biRua8Yu6uOI2RtcwqO9Ki0lYkMw9CPG+AFnTBGuA4ynFMK9E37bW
kUAZKtW1jw5J0wW3XBquWHqpxIdzIBVIvF1uElSoUdfACPyi1EQU5dH3HsWjxKI59OkM2oc+y55k
JRSST+PY/2oEDGG4NJsOW9PHp/qsuGYuENF0Sz0eQFlRuHYKqPYhXVHhGNk6vtAH1EOwAQ3ETLJ5
ak1GrFrdHl2vu2klH2B3N7cKrGDP9bRunKLks1C+ewhvRA0IqgUkYVqMDK/Uo0mLY9bCxZvZFaZz
WRIbJQe4HxQg4SBdK7rxvisUDT1nl2OHDl0zsny6WfbRE0+dULJ8RMS916tvZhTdGWNqD3KWf3Ye
lIsfcUoucQr4sCPh3NG5EiNudu/48XvVmue59uZgNZ32lQIE92+gBsGdzE+leH9763+aKlw41jeb
mQVFKiAVflhYw94uxKnryUQagqHhalQ+rR5j1QdslfRGyaWHFXtS/6bgYbp1SCaxSv6xwBzXmc3y
ncWanuEGVipF6i7zZeCX4mnRhaBYmAN/Ur3piMS0z0ANg3mUzRVReR20OsvBEwOPIzGnQwGPveQB
XwWAlgTE1qMig18OVsmvQWJDunxZTnP1TuHXdDRg6vZxqjiTm7TN8ATBDoylIToZSU1rFyXgwm9u
k+edWkajtf8KejlZRueMkissHL7xZBqSU3F9qo45Nb67OGPGvVBbimXdS9PBH71jZQ+8yybcgP+s
YXgXAgsbFscpwc4M/m7oxt6FIeTvdBF5IsJIq9sc0sLhQi5SLt4qSjqqyL5bcLF2SHopJa2X1EAL
jHH+OoN/usHEGxpCJFqbW4+6zWczzWBRgOWHbwvaerl8hnGTWYN88ZLqfD6DjhQPmIlpDoMnpr+L
SEGnJr9iMGx9RiI4oIHaP3b2stL79U/vtkDMKdHHU6b+KOyqmmXrfmdk8pgvaa6av6lAn0XDZLqk
5JYvWNAw+ScUmQ541LlY9Hwx//e1ReK4s/j7qvttMuTbEmyVvPHZ7LIU0HWTdUP4mSknkAGtdqYj
3ujeSAiVPDELiL8j6vT++uwXK5khXT+U9RVjeIpWyvIjKEoFkXIalonjhdcF32uD7mmlnCZ6MBsS
19iBxypimJEWWKUEk9WyC8e/1dEOxiZ4Uc4msewMKATjdl1XuVHYZPNf9CzWBneF3YIQCLfGA33i
zBahzifEHeMh8Q88cC/UXiHE2In6blPsiZbZprOyhk9O+xrE2tEhCpS1a8dRnx5gLNiLRwdTzBt4
kKXyWuhPtBfWnz+bwSkMXjf29AgSk0sBLjUEOlpuRqLVLP12EbcgD8G5NB7NVFjEqk3vyIhaRQ0N
jjENXVYHyTsOlATE4hW8rYLUfHlCQ2AIJR+RbSQcJSw3u6Y5QZdafu3qUDTLLkAuzpDrsdbDbnoa
FtoVFWuGdy0akYa9YFbjclag76oGQ7jdRmROprml4wayNXJ8B+q9aFuSv/ngpg5K18MfVNTvGoK8
EOvMTA4mPVrfzMiRBGJNkymN6kEhRGWmhZkxb2FISXyq64QW5qfQMJWTvv5nniGO4eDP+KYuuncL
ouyrmGhrh9Pib0yY1dXqWvzoKbvCYCIj5yaab5b6pzhDCpeO5dbuBC5n4fC3hhGKnpUaGu3ZYhN2
Rt2wrPpfDEQZMLnCKaeCrNEFSeHhCGhZ+PoGinx2ks7E4Vh3/8n0uTTNgirzAhv438vvwFDLB7Ij
gMi7dS09wBUaETq8PRO2ZN7ENT1ri5PQkGup1ibK6Q/ZSVMgM/tBVEPKChkyW90uA5+3djmLccg1
7bXEfXaT2MeeRl2jcv4TerRniiwsJtq+BzgFfBrBYlyboriyG8CJq0at1y8QY07qBJLKy5CVqIdq
PzCnBxEx0CtRIrf/6FqWNbfkG5aw6P+OArnLQ/CkmTu2Y7pjx371ZHEyMe2WfNR8/4TrRU73sT2O
s5m2MWVN/+5IRZk5GUFFARrl3dPdVK07hg8lf0+nESkQxDKSXiE9O9LBHxasAEbV7EBubhd5XyU5
TfhiF9SujRT9L+sg2P5RfO56oQSNJL4NEpjMdCOVearRqPeeW20Au9O6t3S0wKTtjj39sLDKwg6W
ilOciEi87goNyDLr69DvS082Rm97HpvQIf6YDJflHmsSZSEHDdmjMUOtESSe/qx8XyIWTBo+/BYi
qXMWsE/4dfFuqDgwrlm+RYqWj/WKMbXGIz8R99EyVwsZ9DP+UtoysAZ3Ec6dhoybFJdMl92urgO9
2byChQjQ5yEI2iWnrI70z3cDUzoGk6W/SzYH0Y36sgHieQ2+WG2qQn8QFxNw/p/ukyhSQmyGSAXz
bTmYZ6iac51M2h5FilioZTzF+RjBWuBv8fFTIHQ4/UbHv2Rgnb1i9Y14PudxaERun7kMfscYOYkx
sfJGBcLj1o4DbUFsivxVdD5fo+K5z03uktKjgQK74WA2mP52GIAYfWuo5WAyJqcKiz97s745YaqI
HBO+2ieOstdA3hYw/bfIyrUSY8+Fv4LnggzOLBq8OVBguf/x2yUKpbkaiEQvYiL+IchdFRpye12K
n8QHzGAIbtz0lEnxpOnZgHehHgZzCegb7NM5qg34EkwqHbpUcLdl2EyO5d1EBsOFPBmbhto3H5lX
VukEwzvxmdPhPzBcgWYViPVs0O4+Q8zYIjnhmocESR0h2XCSAkCIuy3KG5g6oaF9RNrqrDQzz8DL
rOAL2GEkJMgbEk6tXrM2fi9aqTw3camfwuhz8RwdW9cQzhvgHNN//IX2xT7eyjq3QjkDeiWUhHYG
npm68MGhmFON9hdbBwCQm2Lajo0jVFrKwloFnJCz++O/xkZRhvW9hFqSD4QSKzxDDxAeeBfW0+2M
zdLARccoAo2vCwobrTHDhApWYqqqskXPujefhRADM5WywHUoTL9JcTx9aNi1FXlveQGI8UcYrrGz
J5iYihM3yfUCZ7IvVWo+GCZXe54aOACB+v9W5KMyZyw99EqDkg9jacYU02nC02uG8hLrBL6ifqpG
2XAJG9TwKQ0LMArteO2EIyR9QOMwkMrlNS5aSoNJD12nGbpucybhmL21O6LBzCum40AH+tqri6z5
/GungegpYlmYD5nG0Q7RiJ5YMqvu7MQKQCAbuPLEybmQjy+2NetoMbvGewrTR/0SR7oZX7Z7SVeL
q7MIAnlxb8Y3T8IydER2LyVt1gD+zWVPqVk8CfFTGwv2jlXkLnqwc+8Vx439IcwV6rGoJJVFbDBp
0ylL1Izr43x+J/UV1GHNX8lwF7/MqkXVoSxdyDrZSVnejVBdLvdH+rik5hRXIlU06hIuWJI5Upts
HBwo1Y5uelQRAPZkQT++DR5PH6WrFz434dPcCe2sw5bSUltzPw8qWVTMHVPA+T62mnt03omNuilH
um6XX849AG9JfDljO0lywRtL17J1a6LWcrgtdzDmKs39G3UtLoD+FCwn0dJ5tkx0DyXjx/YwTWpC
iRaPVcZfmi8s/oCO98fcvhfCjtkrpYEq3k2VwQRX8+ag0OGCIlI00ku0epISMHs27tIPKDImql9f
r2/dD81CayjpXe91hmzszCWsKyLYoL1u5waGK4/BkBKH+qEgj2Gge501YQXnQ9icGik8yKs23ikT
c5L9pAM9qlVfU/HTgcxa8q/p7H3RzEMbUm3F6Bstk0GnKUo/6zRnOZVFCM+UQH5rNMLwx7jl18WC
i0X+t2h9g7cv4zp5pBhRZ7U8rcfPlygtGFg0dTQ98T2R8XzZmaCHUrHcBSOOAtUvOnVd7lFzKJ4F
w1JGZejErf4eB8BYCAsuGSaY566ZnMqZUm/aWc3hcT/liw0OO0nhGiN5ruGvt3DTGF5vNVeuM78Q
nhs95rU/VeRQyRUrZaL0k28MSFbfY1PZE5D6msnC1FA3lou9GWSq47LlBeIYxJYIhe+dGNiakmCA
Frleg+ImUa1Y8vvyr4UdFiecGpVQlfTv0+3l309nxv7HB2E2sVJ960SHpNF8rdOUGXl5G6jgUktE
p1V83UGIPboON9eEbBmZ/yxOuax8hKacFKZSjELTzLh9Xs7qmIuokdl4GUqOZpxlLpYpiStdVGG0
UDCZfBN70NhNAmfhS6tOGZQjUY4tM0oBxw2PuKTjPu8kB7/ejKDNN3esrvgPX9hQHdE7nVcit1FP
+1CNVyM+IJ6ILtbqfM1+hZb4AqkQRQjA6itj6b/NDx7VfL7kwSr95kaaNQxI9y+kauCvctqeO6DB
zZVRPhIE9I32LB/Jg5Bh7C0pGkrfLuU/DdT+wI6HloDqdFAsme03HqAVApnBLhEUhaXXpCeFhSPt
Nc2Y5+nWqKG+vbV9TAKMvcxjqR/5vL2ecaJHTAS6BW10gYGHNwrmgqm1HVgMfVXLj0ugDTAJoeRV
6VuNzJe7ll42O4CEuO17DTuR8aHwDoooS88nJCjKx7n59IoThpzixtrXdvhrWK/M63DV5Yf/ETVN
d94oSuNdKFM1V3z96yvougoZ5nVD7fwmP1LhWFbPqwvvpwvvZG7VL7IfWcIU6xXalTbFcQSLz+bD
erEJY++3JLqSXli2Wfqoe8xtuU333ttXsL7SJ4mGNb1bRuzCJ1h55/+QRXxMIyoXGmP3a2Bxd9t5
LohV2b8vIVmw21WiKQzfJk2vH5LIlPugXwjuVdUSOPCOYUcX90KMYe7PLMtbnZtkss2M3dQqSi/f
NegMskvhwIyAYcxzBPxXUS7M8HGpLMFogU8BTINrwwKGhTs3AAhmuRrRi1+FKCWWWrFx4FFMlQMC
JEgX6h2TH90a1tmisI7CYf+ZP9i6+GUErDxMURvFMFus3dF1QT+G3E4qgj4OkOn3RlfLBz9iCXUw
i0fdaO1x+EOsrNXyyD8r1IHxIwZCIs+FLxDbTHSXqKqBR4WG4etJddqAzT1rgVccD6HGGnfuDEYO
H0MNFJU1fjsr9SswkcYeSNVrJLTCEMYTSMsglj5n4TYiWk4S8pbbAwZD7KB+X4OBYqBEjAUUO4wS
XsP5s/qcr3mdxAavkjzeGYwbYiPuxcJNhvlHApcQD6NkV7/dkIDmzmk5KVjPLB7Muu07XmZwETmP
j2ivG6KCtNGdiWj9rnAXTh2u9QBy/tu5qDCCnGs9zpPFX3E2mc1i4XY6NrvJWmKfnJ47tePp8rqB
G9PIMU8RsDrRMGiHpKQMjtSJ7XY5LGd7ozIFnPP90nQvGiLXfnddgYVx5SSpOZgM4MO2SxV0G+07
bNWx9YainGo9rArDFiQ87pX+HTElib0TpMxoYcw4xiLyV66Ftw3XzNZm23hW7j6uZIkzRnvEEs66
83MI3se7Tj6xBrk5cVEj2m7Wehr13Tg/oW22C8WcrmBJF2pWkUwd739kMH7BIH3lh0vj3ZZWspai
s0EJCBnTHmAz0iRJSLK4hTk3r1lm33LpYBotlqUFZuLFO7xnXAoaq9sih4WyiBBckgQ65M+0MrCh
2nTeYmlm6bnqX3dIJnctzkUwb93ssvR8z33zA+V8woTFGRdcsq6jLvEtISe53On1aWQzWaX8DN4o
EtWpum3VF0VtTkSuyfSL0Zsc6jfcLmEvPPSQ/20KwoB3pxPLpPlHOePxRnTPK05JW6IG2HSzwr4R
oC0N8flXWyLdkUiBC5/mLIbIin8xsagwozj9Lfw5KLK9R2xR3OoD7YcaYFfOCx2DN/g8TrN8H3XL
KgC0SlXh6XtMNN3XMMN43IopRu028o+1BovpxiVI3CLJ6Vutb2IWVT8bdTqJswkhOORzsQ5xG9/6
6/8oHfEza7TPAMpYD1grYbpgE5b2w1yfMtcakaPNVRzoSZ0cNmn/GyeN25Kh2/6fWhXA4YzCyTzw
AMk8RFkv/ri+v+twZgLHVbhmUq4g/Kx0au7Zp6mvxOUuDD9l0go7XXHQ4PPudoV45LBOy9gJDtKI
xLl95YSoNUjludxInVDQLZIY5LxBaToVQxLuWl21kNRs0JYthu2/go1c09eV0HVDvySJfKclMLse
TVDdW530f0i5BYmyJfgu8ZCxfH9zEiW7E9MTSGzEp7zOB04rExnAfBttBvRo1mrTH4D3d8rbI9VJ
v9aOMSzUtGFlh2jad7Ma4THo+a76Xb3L+cQZBrBYyPnU6sYE6QZtx1AlVWgxRvC4g+XrbLuMtTCn
fnGGZjo0Wyj3Z0QKewfqD8W2xF3JYW+2Vq1ty4YEL8AVOin5iBVPBSMBsgtwaHdOQemPHdcQe7dK
oybtewRDaBGh0S9g+yZRKYhU2NiXXpHhNZ+nuXjHKcP+tFDdoxInsatNeztuLb7aqVGkVAS1oZph
KJ+/UNB28Dr5RhxhihNOaxz8cWlHQa8hOWAJno2txdhQ4dMHCGQ6xllLI1tphU2P1g22TFvGk0/0
JtWIFVxaLEZy/JxoQ+2p7HXNwkeud+VQ9/aqiygjGWv4w5NaQq1mdI1Kl3PWX4uInvifPbOtmoSW
do0jtEAiE/gC5hurCfpbaNDlEUVk0xX0FBVEm1sjn7HVAz+cRXG/CTstOn/9gTqErvLtcHAnXtsn
3cPGisS850wcPXCW2wTPjzQ5bYlNTurItbxyZEBeDGZq+W8XiGVubmU9yxVz98BUhWboT2H3mf2Y
IVey5CFgP3u5w2/J8YKcuaKkb1W/W/ZFhzNOny8kUqoRaxupiuX1Y7ipRXn83e8Ty92mLEcg9B14
G7do9ku5VUznRH5CjaQSL1S6cLFvdFXq5gYIZakzLH0KsgIzC7kwuVvkSthsS46v67kNoVX0b2XZ
sNqPi3LLFp5L+/NgAEbADS8vJv1eQOpfGrC+N7fFPB+pqBDatR0s7E7hmvAlOHrqjqPMkDeF+Uxv
50YNw/feM0LxLSygdQvcbaAndcn5KPm+lrBMNZk6v76X1B9k0UddlHY4yg+95u3tuNuUh/Ly0msO
CCayHZ60oiTWT8O6VyGZH848TkQO9UXVmx50DvHqcAKzvNNlxCGCFn4M2pHauvp7eoh5PVf1G141
SWMRwjNxYpvznZAuTjPi7lyjEtPu3/Fp2AleEjw9mtK7OCdfpkpwMXhNQMtGn6c30kSdE+g1wqiw
yJDv/QIYuYq3cvL5v1RSnBNBglYzIpNBRkmxK8DhxpogM3dF4b5ORCZaIywpsAlMowONH7cZMfB1
bdd85wdhNULz5WCrwZnAVySGQ2ynSybadn0GRy3Smz+05Mw3spvzZDveUUg1uAxs6LFxBG1lRRKO
WRUijLt8X+ZpYaNR1LakIFVi9K3Nwr6UDo6WyAwCPlz0yXs4Gc3+gvSEDJUq6EUlj8uA9X5edXv9
X+HGi8gijDgYeuE1vN0S8o17EpQdGg7POlTMB7uYFskgUTwHLBRi1/ffFiyPwWrAl82I+gJzYlcO
ZC4GJ9j+uoCzYHwGt2Uf+HIzg9InZxreI78HvQe/E5JU4tTSnu/TFTympnVYQ7bXEPdmPuOTyofw
gXx+HOnPzXFE1fHtJsyPfn8D1ZqNOjK8cfO04Sa1jwc2NzuNvHVN8CfOp9e06y6FlLzIKaxFy5O5
0CLGHbJ4Q3lqZU3P13MJSDhCt+jASvTIpTELtMuvDgY8QAm4vTn8BaRZtnhFBQASX2QYhnzzvcRc
VsTyiAkHIaXE2lFg4xCBFzxLJ2xAjAezX+re9B5CvfHqWpggcH0h0/aRSvPIZOkO6wB6367H6oXc
kGlkvVzvlJOJRa/8LZOuWu1mICshwq8K8p7LeOci7ZK5DeViFmm2Aw5uvshuZusSBB2jIieBTFG0
9aY2zcp3i0y+Ah2wPSVBTNKAGTjrq+WmdTOi1VWixw32RxtTy2YoUx2auPFvw7OKhsmZ57UDmWO/
Hfk5bti/ECyHJlkDp1EX42vFw/nEn5K4vOr69E6ko1KqMAuUdH2NNO8H6kYJ5s3TbnSuA4Bzzov3
iVhlj44zND2GE0iOOaoIvwvH2RL2YKPAMuwHadqRPRmQsC9JFsPfudJEHFDRwArOl++BSpevGrWy
hQX7vP+ww5ynnyhE2ZvS3SA99TwTed3jVj5oTl1/M29MiIg0JJfFG45slz/l91l81yq/IX8eYOQO
yYrH7vEizk7L4mvyK9cHE8x8Yh8/smcfDZuCRkJbHHLaAqcn/4MHw1fZQO/8fLy7lbtrYCWDA+lg
BHNJ8340yJtKdRlbAsfeLAPLTpIF+MHb2YZzZ1NvKqFSIdLzWSXe/RCXCmc8ZCRIw21eCcBzj/Y/
18nRjaGk7dytJP0PzfNIyhAaOdov19MQx/nk1zIHvgVhmgBMOALnAKHFaa6hdAmM17YB/9r2tAyu
L9ymVGaTEe+LyVgzzKE67z82MYW5gKrc/lw78yPkE6t70JQd9SqQCoF30qJBCDJxfenAE6j034Qw
zkPFnWSONFDi39J5keQhTJ7EmMDtYBxpmzZboWep91MC0W/zHMBEgoxXF9/cIcTUEdrqMyFop9vF
jvP41vquk6sWX5ZYy+O0Je3+xEHcjY2lpXonkQ6tloNgSv2k0Ja8otCbdHSOvnRxIZjSCkcBCZpY
kJnBM8daNwrl8ISVh5EX8gaLrZq6kyvmF0iNKlKrb1xGDyjRgG+yioYeXkdBzNIKfi28UsTBxZjv
0CEmkV8kv/Fi4tvMaXAu/Aj3718YOxYpgarIO6X/9hSWUGsrdOS4GuqiPjO7aEetMYOSYWL8U5EO
XGDuv6LmdNqDYKBZrx4dphZ0ZDkY5+WCMZRHMDnFNrT1aec2i4n/FutqnJeWs8lfLxkt3zmAQffS
ap0xYpqp5W0v6ZHivgzjhnLL04/aQUAtLw/n1SqDhmKpyLmTmIsdMx+P/mw9rRhAt2LOtHQOqbPN
kZYd7t7Otn5S+ayoNMYHNg8FEel5TCQIJkw/rfQswvtDtQOHA35d+p8oxi7bTwQrSf+AK7+2Yp+0
N7tHzRrxcmn2KtoGSUgd3ctMvk440rB62yEmCpwgmU0P/MGCrIs/N8m/IqSUQ4b1fw1tDHG4RQCU
K2oth/Iok5wiD6LBagZdDFY2YPoiCk550FBgXXxCUTW6S01hoOFtrG8Zr0UvKw7Ehg9yHl0ge6/C
NHQ4yx3Xq0lCys8PPRrZl7qLSrkMIOZrEjfthomKo7MesgsADhNQ0u/rThmDmYpMFmsI3LBtLsxZ
cOMqiTKGOdgwp9xDJG0MjFyMYvoylwN8rvMqPKqOFP8QquaAuQ0A4clSdyj/z878N6+Au6IaDizd
jYW2QsO+MUcAajR+D5C+mk5mT8Gng2GnY55P7pC6FZ7MXPnqmn3j1O4GS6fvR1LyGm9KxTtPoLc8
8/XYkBV28qwxpGiPjqouaN/ep0jV7U1xoliemZwo8/T2CpAoUPLswhQJdA9Wo63Zp1LwhC0sKeWy
CG7jQFwAMQ3jlgvfFAR3mQAQ7NFu6BDmC0T+dBmIbhErf5RWUm0lX+XmyjvoNFd4CCThxqtA6gzW
lm2abELKn+cRKXCQDtdDtv5Rc5KXfaJz1u7FDCZtl6/wDXRQEKKm1WM18DWeKukfrBkS5VML/KY4
4aht0ZickgRgNvwNj4bqEF3WMyE2W50pK1QLd2mrniXwJxPJYd0FuZO3c6pXhcwvPvYy+OkzbljP
n8GfFzoQVoG1oxpA4ZcB75LK97l+aYwAffi1NR4Tp0wv5cBXX4IBLBf1GY3khY+4AvFaXoCW5cuR
DpGjnxkY8EOp6gqReQ9LCjqBBOdAzzDhUi3qdp331ryV7Q/Q/hiv1WRPh1jX8R9dYvIP4tN0a/yh
PgusSzaphDxazVHY92XnRJlG68Wg+luVOGutXJw9zF+rYTReVuFQxRYVFHD9bhhPL6VS3aojqpup
7iYw/lGMOYztp/CEw97mch+14PrrwUkkjYa7bp3VMg8gwaWNFypAAvQWlcT7ZQ9sZ2/DQgEEGRWo
i0MoAZTEGTmrpDg4kZP4XJPTY26XrpIWHvjw0S7IszhHzE7t3BGSeFB0hY4qEuDu4EO9PAXPHz+3
OTk7xzeU0wnl5ajhHCecAa/fvovdNir0dszBB+mJNm36lQGr6pdNKxOw3RO3D124fPmPaq/9z4uT
DQjjee1JxR8wy/RB0acLBCKin6oVZ55kHOWnrEDoM+8UQ/9LRaDjjh/ffbN8yggqImPtHepkKyuJ
KcT6FLnKenOoGAWsMIBkktajFN8sIMad42/19kJJQVrSoFhj46gFTyN+t83pHChhNwLHvL5CAaGN
IMB7zPoMUBDfJHFllJe5suLUJiSzmhaJAjOvE5mAnEDnKicc98P9R/N2MJgSBPqcQB0HljXJyfFb
9p1tzrKrQDL4V1tJy6d+TrWm3hSU4vcy8ZM+E9b4WcMh9Qd2hpTKE7hUpwIzh5hopnUM4lx+rTvA
n7939IN10e+h9+rVzfzqG7hH1cA1ek+AB4VxC06+a2aIWoLT7NZVe62hoEFPCNaNXVVHNAd+0h6w
deomJbAKspF7vDDbWayQQWMpMCWbJ8skrt8pdXlxdiIBpWRCuV7WKiSJ4tzs7Uy3cdGCM0h2YnCW
l/W5rYd8PjmYcUqFEOg8ivyd0wVIMvdArmpZjR+Os4TrC+SbDqm1bFhISBjEjPMvwS8jEMhzaOWL
vgUJx862W+fD/X/MW5vNLf1i9hJswONwE7Jeby3zcOnN7Q9imFmphqiGEofBHdWDairl+dFowKIE
RQpqzbnGu0fQXXkjoHBpQG5hiV2VFkR1A0h+RUtIxj2WKJleFUHjWPr8Dt7Zbg0Gc3MWVoG3WPQW
TsFdwwk9QCBxHV/Dw1Ve80iNFZQRGN+rtYMPo0YPbLv0CE3PkEitAeDUDQuj1ZvszIgLBNJ0+m7h
e/sKaFcv0N8tbKA25f044sOJROKeb9IO61VCk5rStANY2Mwm7tguUSVdquRBQOgRAkqz5+IlmikK
l6OcEcePX70YfGwmRTGZ0yJOojAJ2MCyBjZbWiBpS0TTFwwebYHqXGb3teGnyL2D7UQb6zQLSnck
bDbHQnt4Qg4BOzAq2S3+OzXKe+H9APoTlMLI51eceiw88zWXT4S2Mk5oU9bbqV6fhy0ac/NnRGdA
WUyVeuZK/LZGlCRb7sqoMOQu7du0ypFkPRUAL94uG7l2UCuCm58+SSe1sG6kvakR1xMX28NZ7jQd
WZL+RluY6m0f9UzXM473PD7UceA7VPvgEH6JxMH7L73RCbsblDiHA+7+jeSK51AQb3KxArHDzOti
wH/syfGP4Jr2LVWyY9l/CZiKtUPAPi2pEgCz01xAB/ITOCvqu1a913vYBZhgoxFLIHVZwOQ7Eu9B
kWDXr8IN5jmfkSRcMXoK+sSV4iItHAvmIXw55gpClMr+jum+5TGD2wjnyRkH1IUL3j6x5nnfXnhG
CVCIVydMGhTuT0VQLVI7CF9bsQ1eNXX2JrxQGPVN4kbBMV03XGSNMRujL6RRrGyatpjDixQQap1g
XIgfWhAOKKIV2HAjli0uTIN4Od7I0+IpOyEhtLjVUUnEZwsYEe4bVsQ2GQIP1shDvV3uJ0g0TkQh
p6KaH8gfde+slrSpAzDMtcADZ78BMKgIGO4zbaVl9n12O/xfgi3qvAYvnzIMCu+ICq+sUwvr8SLI
ZSU4SpqHavL7ay+nptUE8tTkydTdmag0wiua4IF66f/JSUlRhBZg6MnQL7mNaAzB8ldIifQ/N7M1
P8vzl7ggmi2hsxoA4U/mUsD4oV89SKTgPbQkDj4Kezw/DTA0Nlc3pALAvY/QjA12h6ML1+BKLsv6
sjM0SSAd6B/pmcvNre0G/u6ZH8O6OjAgNsSGNqwz+NhBLBLqobgguZB6RqPHchgT1yj5I/HqlwU2
XhJcIitmXeGMJOiJ/UHayubOHgwEeDDyr41MdLBwgBUZgo5Q7kU1A3U51VAm9E0qy1PwEWFZxZv0
xpU6XkhkXSenbJ0kCPSJyQCFqvbwmk8XbeX7rYsacW0NVmOCFC2Ro7q6eIe2vSY1tyzD5OzXNhVi
O7K+9Fmc0cyCBj4QEtkVX/9U1WLTGvZGjJ1qIk0vQ+oaZTxAus5pyTwjfAczOy0z1GFYO+m0wdDp
rDO/w6DP6iS5VkjSEy+wG2fJjdiJQTWAMUp8PNQ4M1qJ6I02MikGGm8Sd8KlJGiTwtCVnjhrvNB0
9Qdgg1AJQxtsZTIQab1zQwzK74KQeKe6oEoPHAc0JLV9+XQAxvffapQZVZdB+DNLhbqVY+TFQSQv
OnYoURVVY5Vfr6mpBs2Yvx0WGZpTXuCdXs8+V60CM3mkXhJQ+gjQUGBMPd0vsSnzVAfThc7GyhrL
1UX57eIbRnqNWCCnp34GFjzUklsBIiJf5t7LmXhzIspRgzT32wOmL+ggX+5XSIX4p+WALRhsS7Tz
0H4nIMoxISRYJmhZiUDLlhVZtTTE5qPBnl+D14mdKIP8Xfmwh0XO6+JW4NTK0R2mFv0gksDKbsio
mDnE2Sfsbe7601fgVV9TIbvnwDXz9+QrtX4NM/Hrl8ZHbVV24bHdbUU4pgqJCdckd7bC61757PtF
h9DpKMR0DrUtfPNe8Q1a7bRTbrTBZOjxqkV/JbbCP40KlzNp/7baeLXhYUl8zEWee1NjuoXTF2Sf
Xyohq4aqiy/9avkXE/TBR5HNufBaJ/u/n2m7TQvb2rePBLoSxScZpMUPaqrIRbpgJqJgxqFiTgMd
f4AVOiTEgE8CZqd9F/JxzGRcht2c0yAxDpiqnf/maIB74exr4z4BcuevvynYBKLUAQrR+KwFcFQZ
IQUXImn/6qtPPcaSd2yxiFk+nuNy+w5ZOv9S++gPB1ChdRcppSplBrnr9dj/tWOa83D1DC7anRZO
Hwf0nwYa/YPODbUq9KPqyri00FEGaR9A1f728nCgNVPuNeJh+yQFTsuSndAtRHHeYsZiJYnpO1K/
R3tXOmEOl9thiCkIoBk0XGKy+RmFzW8dCi6yK8tJiGULbM+bWDTAsHJ2aND+LWhKzshizWbBMns0
1622eTs1cR+G20WFYgr9aPJvUUAf5heHAgbKeUa93SE6VaOtzJ7mIhRwQYbGuUeaX8wBIZPhtCIR
V7mYS0/J52626Sf+ayHT6cWeA7uhVDH2B9u1pkYefp+kdSqbRxzu16qgCCqdVTNIeL52Hc5kWgXD
pcYVvOEq8KOklojudwhvaZjMUF0/A1CYIeoWohq+yN/sozIAAtQ5Hr2fQPjIwJJDnZxtcUVKWbpP
Lnl3P/Oyoav5o25ftbxZrg2qvvYHtx+ph1DFbNuoDFvHqnqoCPHRKXooodySKsC/cFgDEveBuQKf
E0Qmmc1e7H7lkEr71XPQ9ww2xq45EQ8QzdVtzgOwrKbKrCpNEW4KKbuUPQXJ03N/Hy0+da4fcacZ
OxcF/sT49tK/FZMiA89Lp66Hw5D0N1fjPgXO4nQGin3M4fPagOFJTcATsz2IKt+IomHB4p1EL4FC
Nup/Dgq4AbSRep+b3PDuROxuw0bwKPilIia4EsFwGY9t2nY4i0+5ccpqUsg7kToU7jQhm/dNZ5cI
4sHuh8toA6l4rwfymDs2veZ0iVX9OD41sODZpvTdT2S16kgUJDDNcr2/TAHybseHHJzu/cjWq3yN
5CxJQ6TuZJW7IblAMejl9gtoOqaLOrehvEa6/yxlaBWdvvr7XS7g12gjYEoOh0c7B22BtObYAycS
9ouOUnFGoEJpfDM7G3xQgcm92KOLQKt4tQ4im3Zz/i71Qk/cXpwB+iTyTxRovojUGkAbGT0C0/SK
1sbfO5RjAfPb5VG9ZAPpHsXJ6YQzXG1z+skSI7LsRdg57EloHsXwrNmV/CR8lwYf87dC39/62iQp
/REnkCyBQyZ4pgKKPQXs3iML7BIKvdtVBMIf91x0MV78xjBd4COqoiVGE50FTiuVsRrk1WekhDhI
0s9fOG1B42tg2oeO33TfhWsG5/TsryEG99Qn6gLch8Rt+mZjTT7XTmg+lp+ipFgulSC8WxiRaRT4
Z6nkz4ukuwZp8wntthFCBn61fkumdG6hbAQpX28FbV2+ZKkbXBrWgNUX6svJTslbLR/I762iezK5
y0qZV6Umlfs99yLuIrN+p4J3IxnmlnD3/eYd2H9kyuE5F1uQ8syqNXm5KVoIZFf5vjiao/F8R21j
QOXQpKEtt/7MhjuZET5FDu0BVgyE0NHgBHJAkxa5pphSHwaLvZoz56H9Xs254WM2ULerr3hr2+v+
kLKgYGPO9YYQCx81z6PayLq6dS3Owp5mhycENx+8oFY9mlgVgvGUtHU7SroT9JmS9KWebSBk37pq
+Jngp3Tk0zGT63Mdyl8xD02tc2K0Kb0kVTDhw1tfXVAAP/jAHuL7KZH00Jkl8ItAuK1R+ewy2uRJ
Bq2IOCHY9W3kJ4yPLGPPhxZEINQd8OmPO9hYK1vTb9QeimDYlrU7j/Jg/5i9KyJsSZ6fojm/2IwX
SJAVBujL2PE8Cz3IsE5CQmkqUZZfJ5vai5X3njk9NbHGeuy+RFGoRH7mtpAJ6IoIRHXjS8HAjC3a
T9LAEsndnaYA14nt324fbBo31TQTn5xonJsH3p+F2L4/fXT37QeGj/rmyfDHiT0VB8p34bcJlr/u
EOz31HBQfwvYLkJo2JfeiWcBRujt+wRbtYsqQY7HUrcmzg64igXJE49cECLgAmd+dd9Ng5R9Pad4
w9m4uQV1DKZjoT/NZprbPYZ+Xs2le4VC6nPxrSXF+MPsrdsv/c2yoQpTfFZjUCrG9tYhRBZ7M3GT
stBFQRPCkBb8sClVlHvqbSSfW3l16/yu9/VQkdQ9GIT9nhRFR+NitxKlp8OmCt5LWC2R5NoaNdyn
VJ/gTMKLvYlr6kz1VtFZmMdgbrmHEt8mBUdVKGFpv+dEECyUnvxjpdWuHcsAvafHDJ3EXa0i+03e
IQZ1JPTF8KQewfB6I698XwMm7EoddwRKGw7CGSt+RVfEaReTnrswiR2+u4Qst8DRE77GYTUKPJuS
I4HqgqFghzuR4fMFyRUkkENqRD3dELovRqXetN3m4Uyk7Ythw4rirb2vO2o1ioiE8Gqd6Sh69EDP
qimsuRONF6c3t9uL0DNbL9Fhicd7+0PShmkVCUWjCibIxfB3M7egfyCKhMQtz+uJn6yXm618sJ6Z
KTEhjnX3Pnxi9I7ScYpxHHMT8+lh3c9zIUrrzWBRhHyeZnx3SBpQbA4JwQJt8aZRw0PXayoAH19F
RrUhhx8SVS9fgHf5xUAyZ5ysJK+ApmHjVsVuxdFQtuOjjMbUdZaU1geonthkPTB+lrJCsZt/ewgE
2BpJFgc+UEp1jpsm5djtwtcLsPFmrfzJIqTW5KeF2PP035FJZP8lMtz5CsEa2AICsS7Kp9GjxA2+
9SWxlZnLLk2cCnahdVnIOwXn5PGS+D24DlYVMcoRyzasJOeHUkKKuXuVH5oCjQaU5C3cIPhPgr2L
fkI+nz2sOz4osRH0gswQ5xA1sd7rNeRGBpw0dXwLKgwJLnwlPe00jJY9eLa0oZJIyQU2jEHRJvG+
Gv54i12y7vqT4uA6erUI9esRP8idCZkBjsqjqnS4iqUSdE3KppbooKpMYk9B4GrUUFoYCG7MfSbo
xTq5+p/EA5uKKHG/V14gjUGLXh8PuVkfSS6cPmRvDr1vMHtgrFQvs5LSjpQAwAxCLbxvk2VX/bsB
eSWkESXe/yBVx74SkXPrgq1vZSw3lUqbNX86SsRqkuCdBwIlw3/hMy1uYQYDnr5pkFl8Y84GH9xE
jue1grhVxoYlfUJE/aPElOsxkwy0uxz54WnsKU92ddQlGQKU/cR74ux8rUEdXZsorjBrmCwa8do9
944eYY2Bs9YouZ6GQWlsuZDnWZdFK7LUlJr9OCpiSFYTrzfbiSuZJQNFKPjqWEXyFwhLtAZUeF5U
pcoFsMGMzpx1dpSDBtkzNgp8EmC0wAHxzNjoHsgw6D6WASWAc38DpC7iWERfjhia6fG1Kyfehj3i
hc5nM9YihjuXUdudcHrA9du/Do+9cgRLds+YXNcunH4IZBakEs0loX9fGp9h8QfvVO7uczkvNvvm
G7DhrDQXiY+qIsh+wCciX/1nD3jnO0P01jXB5rPlxYCUXZlDPGvOTrEHZteiqxWb9zswBip8fJcP
zSNhxQBZlm7WTJb5Lg5rzZS7wZMj0+cNXFPRaOMG+AOhUzLMF3RLW/ubdUmfQ4DLSG2o6eA7S/SJ
YslnJ4f9WxyoePl38EPxJ4cH0AaBUfkmSsBIyiRTvZRISUGfwj/HJGiRylnQRlRMS70kUMQsNIBZ
TGNwk+98PNxlWNljC3a9h9gdlDuuYhixTmWwI16+3Tj+jrwGarUcKC/fzlvX3VeLsR4PuS3fvK3I
GB0hG+G8/WJlaAfziChimLVL6/vxhHjyzmeo30JvEYqZs5gpprB150f3s3MesGa813fK2gfjL42P
EmsXwtI0XyzvjlPivKNdM48Lo3+6cqpxdr/Fx0b7T5v2S1Y6RWwshn6uqYv6zeG+XquVUmKefW6r
fslvc8Sg9ZbaKRx7KZPI1LntENaTmEVnsw69e0Jw/F1WXv2CEZVI4HefpPr0nlaoKUhSUpUoOEnO
tQg8s6lIsjBtRfs8oqYprrbDJLQ4KkCbRHQCY+oH0HL+jv/kKJaW3uu0rfhyAMMLULXmR6Mx2W5l
htE4/XGB9p4hHeMDs6QZ0s83II3Nil5Lb4Y/VgkAMnn+i3PqwIVVqE5/sUpaHasFm+VxDXY4EN/Z
bgGRTnn2zgygHKXFttdlkcItsg7P1DzZ/Lqge5P5Sba9ClptO7bF8HByw6Vw7dvc8IWmEmGs0FwZ
BSVkn9yfIPXXEbSsOlV67kzI+UIerbtxEvzsioI2w9iYqf0QS+IIvtnGjehneydP9fAz0ggZOsOO
DTCZCkigw9JUJqwsZAJdq6qBdXPtCL6Q0goN6e0E9cmTiO3KkeX+8Bf3OkyX709KPD1XaCfo4amP
aZWhTbUbkYp0ccxaNdcHJEy+G2bhEDn9sc7vyNfXKAHqXPZQ/VslVROxaEfqCnnyXT1ZZL1iZln2
Nt377tte7riQYSSGlPB15PvOMr1dAwudQMicl0YfNEV39YBfzz5KOdNlmhW8uOIlLXYHrGQfJLBB
NrfyWgkx6MZryKgQYHJ+9X/MvLWQOBsSmF/l+atwHLNvz72XEgDE9ZMdSdKm4afYEoHBewryjhUP
mQimqdPU7IH6X/EmIpdBnBEu8wc5gapaG99yptYb/JWYyZHG1MGNPr8cHingw36XnZN/iT6qQ1oK
ulcOf91jUGk/5YY1lIfaUMax8EpO64VqaC1G+b1mKZEN50kwoCVFWPB2QzD+2Y2JqaIYePEaRDx5
OSLWXZzeet7Ho/LuzcDUg9nNth3wcwGDeqDNwFmYHzv+YZ7NkdXf6XVP8aETb+/53GpsxMM4Duzj
Y75BSHSI3GEg1fwwg+hh8zCbChKNrLhKG4UDT/1swhWL9xHdMMr8NMMwxhZdDlksUiwF+iMPOdoj
i9j7XCJLacP0n+TzGVFY8LFo9auw9X7kLl4+NXChYIaRBAe56UyZEkGDZLYZ2ahG7NVRVwLuGfxp
QxvtrwN4l6DNaajCAtazuGyACc526Em/f3bPV13Au9T+z/YsVTntvtf5epFYyALj6elLa0fJyBRQ
x92pjlc24FiI7F6fN2NqntLoEYhqqskw3O9XWVB2wZjhqAyHzZdM/l+SGlEYYBdY+XWb4/6PQAvd
WmuPE2HfP7RSOiDGSzXVAh+xFm43HQAbSTeAfhp7xh0pi57ULdhCynJw7a8DWgz8RA7vMTTxiKQO
DIFhQ4QHMvs/w404MEcM3xPAjHQRLCV2Y36M8PPv0/r60NtgG7OyocVZep6UsHQA0JrI9jVb76EF
0RKo4V04q1PDoFqeX5hiXndR2xEbmJv06oGcZXD3iWAlIBR/cVSeytEHRdnFXgzd0OCveXYYFrmx
JM1rddtSg5pfQi/27oEoHzduP6I/YO9Rn/LoJSLhL+d146HuehOcI/7AcyRM/SR+omX/eEn+Y0yN
vk0DzeruIVt6fNGs5hw0jaFSbE28YYMQjJtiZhtCEfryt6w+R8+UQEI1K68uBECZitRGagCTArEp
2xiYzJVH9poJ0uQhAy2WAOyMmFhkOpk43nmfDCIVxohs5QnGtNYNsvEZvRBIdc64Tm57UjP4Xhgs
SExRDEbiH14wQt3CHwLpTAyixDIbqMyXhfreebLOyStlqgcCnU7ACvMjqfQOU/V1jpHl68IiutTB
NZA92ZvZF+amHFngU4v/jE103hb7egqrnWaggMgUb7Ci0J8RtcEU+giRL4OVIh/njMNKvv+eq0Yy
RMpFUaAtLpRn9KQoFqOt93+LRpoa6wv/q/RcLDSF/REzQIzrZO/laTAZuoOsFinpZFxizAr/29Re
AGfccxn66RHUyEUR3cr4pphn0bQruB132BB/Iv34LfJO6s47eLQ3DTmiC74GXpGhFG4bVdNrdV/T
mbkH49mHHc/VAbA1wiVAvaLo/IpXZd2ra38uZNMeImOBQ1TMi4SpFc3n640m+Ps2IEB5yulH0mW/
7p0BUfTfKZCwEZgviZUL9Zz+Bf4KR/a6rgJR0oOqTEz44xwHELGyxRSRYnyeftJ8oh3PlTs12bws
Li5pmIt/uOi6bpqP5IPri5RnWqJiqMVMIBJwLLz+li9YKklm26Ln/I99HluYmU1f+VsVJ9ss7j7P
bfwPkZtMy81NGEQcH1eL2RJvCmnV53PHi5+rpPzM8aDcDLTY6Lt6stfWnVlF+wDTuXSk7ynPtcdD
U5ePESAIDoV/eeO1WNvfqjSKDS3iWdwKcZ5+0OWSHzZj7nX4gnIFleLC6CLm4p7LnmQwd2D8w6MB
u06BnM41X+TllYoscjqPFLWH8jPDXjzt+8G5zijKk2lBSTWpYiVs8cehwcpERxLe0M+1DKwpev7I
el/06B6ai+XnXCQbLCeFckGVNkhVVs+mjNCtUcs0rb636QwxJrme6d2hFo5EDCwAIzUri8XS9PRJ
hMMNmpIO9FQLb6QdgtcpM0T7oyte7TPMwIreT4I/Ba9Vildm5S8Og4M4oOBeIeWIjzerUBjsmbZP
w9V5fYQnKaVjYNJ/CNm0v8epBVe3ZIXyvzhunsiRpz9ZNig8vK/g4hQRoeKXGXLo/DLIKZOlOkwI
1mF9/INhrpICSpZeDV1aHoL3LCkk0LVIQ9nTdXVXQU5Ypb8pCA1anK6jrl9A2nQkVq3fFL0ODEVr
jquXtJHNV3tcHcromD0oW0/aWtv87+77ZxgLgUiyqDjclkQJzkksWFQn6rrdMofU+ktcJAQv402B
tdrjxkRq4RcgLY8IOdq1bjSkV390q2sEEkD1w8DwwT141rvw0N83zCHJFuuZFb2qCNSEMOoB0oAF
lLs8rreXb7VsGhp8NTEd3jjsBIIcxpvfzZNq/VXTkZwuKWG575PKVWgGbb0W2YTKKBevzpckhe8p
oR6KpSXYU6Bc87jf5lOLZl6PyC7zsiFhwNXMIO8P3mJJ5G882pe2Wt21R8CNBjSZ7jb7EMbGOcCc
JhFCaLCuzseZ7jP0BujBsGBQ5h8vlBNYWN37c+SASJj27X6Kg5/oMd5LFwYnuI/wCo7aJiJxYT3r
/c+azC6pR39vlEIhma3xYrYBSPG61npWmd1XCk1izMYSEA0faofg4/9wM5srCJtEejGHQC1cV7rO
FwIW15/3wlmZn2XLvra8DhirqcolAArjScZYHmA7kHBdDfM4fvSVKmsKM001D2tj4l8yQvMYajRU
S7qe0hfORnhD87ByGvxEWTZDt4FqPj2FhxjgqivuT4Erel2U5wF2yG0bAMDFKQhyVAzRbtBfoMLJ
mQUTuvqDlrFiquTMr83C/VEZDUY7k+MFu1InH+A+pc5Gmd/QiVQxJjDJxH7tsb54qKEEYVR10MWj
t782ws3tPk7sIeldXIoNf4qldrMuVi8fSUtouXyFU8Udj9eEKcckVYHqL3VvXepIQ8ZeBYZFCMXf
KFnogdhjzA5Q1vMYdiLoFgURKc522yDkNYi6bx0ydbBLdJ8ts+MDPVm6wSB6UElFG1izQf24KRgA
Vwk3cC2jYDV2GOMx/JBBTlL+qh3NNlKhNv0FqH9uwOsPaZmcVl4NTpAZny38ZBCB2Qbpd0qEKEoB
bAXUR3inuFKWieymW/xrC8rzzulJ0wMlAsgOlNK7HRpnTD+KwFieFFmdecMyT1HBtoaJbjPv9/Qd
V2RTLKu/7+8LEp5TIXT96acWGsRUIaG+0BJuV0FDG9cYfFSmedCTsnpb1YgpyOkL6PbnRR0YG6Br
++zpy+KYf03B3Ff67EhvrQkX1c6MuciYxAP0J7F2wbtZps1QKQbmJ3bs4CpwTfWNvQKsZw/3VIy4
s1stKxhlFZdXzT6ksOH2jDBiyY5lqfebaCA7UR1aWpzHmlGRczSdL0WI+T0ZD5UFcFudBYp+zZLc
o1y476lCtx5aTJ8zy+YKwvFedlKEgV//psIsJE4QXg4BCkTpNMdBBmJegamkthXi2k4UHwkx49Hz
QZigokzZ/8gn0Ef+W03nTU+cFGuwX8/uz5+ziZYfzgKcV9YFFk7wWqdRcduf26hbzqJ5mUF7zDzm
Iih04J9d6icXrT0ok5NX/s4bD0qM1aEyld8sZNcqsjO8Rz4YD/wX9Htpk85f6t1rfQsp5Tuby359
h8ajqYO5/woBTVws7UPwZSv0tXCAh1TZsGjcfE+9AGwIftMKLC9shV9rF/S9uyexnuMZEVBqvPzp
sbaYsJRby/+LqmECvuR0makF0RXqYnghmIKp/NwgzI50qc9VDZMaDUuqejU7PoDUWRY2775MkXdf
eEhp1phrvBaLvrGT1DLpt2YHK3nLzeTf+rLncyDEp+M4pEkalxeRliFxEKO0VOIeAQc6eeLhdoh6
EqQuWwjxrd/92AJtn9KAHbDFoQFn7+CXUi/AY0LsYM3iNuOOoTyRU4VzgNc24GqO7ElLby157buh
c4eXqw+c3NxrCJ7TOdQ/+lvdhwY2u5EL1fs04RTaWX91hXoNy2Fa2qBOKF5mQUFdj+xfywR0hE8M
rHahVtEbFlP0kVf9JZMBXVVNDGrltyPP5jhfDrlJfcK00UxZL8jLKIndT2G4whx3F8iqUdkACWTn
HDJkdWthJVzM/rP5NeuqeA224Sqxkxom7opkyrd8fvfHOI3PboZQzS3Wp7isr0gBRHCFhRPBoK8x
woX6WoAvCHHUG3g1cTEaVAFav+ecScDjg5IACa7/+5HlKzLs6XSm5UPod3tC9jZwjTdypASYjdZV
5wLR2HOKP+31mT7MKFc53e2oQaq8DyBvJmcqgetoo2keIHwQhv91hbEGnQJyZDWUfo2ZnfrnSB4G
dBqODO3E1RtK/Zlo3Klmn/zoLwwfPK2Q1mS6LitfWill7pbLXegrihSChWUzQm2m9F9CwyWZc6vf
YEi6VSBRmJG30QiEMnyO9n4ZCO/eHJLmv28O5g6xjbbgtl7tIltWxKJiKvvUmAPEJTE6+xo/jdFp
OcRv8agJh+FcOW0CESu5oGlAcZp+hAeiPH9xVSrPtw9lO1J6IVorgbfIPlxVLfg0wcCvsU3zz6Bt
nbbwwb0kIPLb+rVJLvnHF/MrCs/H0kDeTBupzqdhg8wVx8FOhfaTIXhoe/HYTUtOH0KMMCCAxb6n
3D4fajl4XVBwMNJpyuMPRDkw6RF4zJoWckp4W05UHCYeHfYMCfs0c3SolEwW4lJ+jiyo2OIdtThk
OKEsJQgPx71Bc1Xc4gH4fob74szAVOAF3WvCVa5YYiSuRwi2lYYCZtn1+5AfN123DbQib6Bpm/iv
FUM7Cix9VZNqUfkhJXbNdKJ1kNwSuVmO+2ZXWmxSQkdgWM8eTUJEqhH0uFdqs4CQ5tiZQY5NMu0h
hHXeKlckdSzwP81KV70vaFFWvcXVDHXrRQZL3p6WPkKafzg5URxv+UuhfbIDTRdXx22Q6990zC/H
lqrAZBkrrnCBzjCPN63MkCp5zrRneVeAZ/229/mRMH5stJA4D9GM0bRdc30+dZxsyaGjifveYmTC
PyOfkvU2po/6B2gmHpDq4jCYPNu0OKqUiaLK9UeRf0HCmJlnQc0f8/SjF/4158AoqeP34URfsFH7
KyMYbnppjZHGzcG8RP3Sl7GJNDEe6sS77mKvJqaUYnU0RBUPkjcJVt2ajLdk+QQzFcbKQqSYesbN
Lpvd87K25aT60SITlVqtURjloOi9zd6Q/cObZV0j8qM4Z+NcMTnEGjZrOfzFv/wS2/S6kP+FedDp
gfvsqAsE0a/B6fqyDE3tXzoeP2VP+PNN3QSq2VXuIWmu/RuMDpcsYq0SCsLccOM7qybG5G2ooL7Z
BIdC+mdGbExPt/XFmUbyYVsppVoZAaWW+SotAruYzUtehQEi8cDgdr+QBwUHxKIlpcC+8tZBPosL
js82pUYbnyQ9xsH35go7zb/qQeJQrjGWVvGP4+2iCyDH89tyHvvl/h7loiKvA17E1Fg/VDh9oI7x
I4SbfY9r8w9Jksk3JCzPDV+9gbQ0I0Nrpzr1khUDWWmjCNDGE9mmtStI5El5SgUaSG+W7p1swbzp
qiXDvWXeBKk2AuB6LHbcF+Vn89qZv/rvCqLvai3Jxi854IRE5LQtihWv4D4c7k8do4fNrUcRSWp5
UOkcqY1CjxE7tx+cAGBhFiwrzdfVfzKENAQMwOAr1HJWDVPlQyhZVAM61F/W7Z9dysjk1ZRzE9YE
yu86R/WhxZ+mCjn5cM4R4oaZZF0IwQC4gNe9NO0oLV/NYyh/vxj8gQGFPGeQ6IDKfISkqe1ezn+N
ztk16B23ql1ydfVsrAyO6eITpoqXXlfDXvGDU00GhTAQFKeEajKwpTO136+HDizhTAKbIjrij3Qs
fRZQnKnwOlZmm2XTcudWuhQTXrRVTTvjRlCZIPYDg3uoIb2cLFEEUJm805HB9++hSepqff1OLTaz
MKN8CBzr5n8+c/NjXXaAqwM8h/txrMaJrY4u41whVH6QbMn65F9u+WPAgyspDOS5vLQ1+5HqOzNg
GHHUqzLouLbjilMAaXjHC87R0u9Ziv0hlNbKkDu473RJBCs4sSnVWBWfhHyU0MLXJIeU88OEQ4BP
P4hSPm3jWzHNboaIqV48jQD1psxWdMJizqM5lr33/cPtfpQPfID7JlU5wLo7GaBDax2Smi6jT1+2
dNwg8oaSYzmnGQyYAHnzlB6vYDW9+kjPGi7EcJNt+CFv3SQ1hUHupZpVLFDRrpbl6O/oC/dh7uIp
/TbniXncdIOlyCObhs8+zw58ky/OgdhLnaCrO3wdQBtX03LrkxigJr5rOHti3j4yWLYFj9a5w0Y0
mmgT/QIYGQC8ZVqy2SHxTxdg9Z2gu/5yKjfZT5b3EZ97RvDkZDdV3kBwBau/kEvub0esLl+rFuVr
Ff3Yy7AAqpQEpFuaXgc5IsQyNMtmJ7K+EYcAYPmNlP02csPnBTv9y6qVHSvdLU4+gTKRkIBfB5IA
XApha7RyyczguRLUVJ5HQxaLEIqDwCSTxOesE3b5zyxxbQKYRzJWTl0JBi7SYwFAiFFgiSPLFaRC
NzNW5TEj0ocQDHcBo3XzbL2Ia4oHRMSxk7xC5jVOMBEKd712A87nVjpygE6NjJqHaEIiSBHeQoPL
w5dlbrKj/S1ReO3XrexWoMzLVfRqW5c80idKgZZe3AVgwjdfosvcCaV/Ud0GiHN9MP3YzEfeBCrA
f1i1KxpoJParnjh7G7C8P5UcLSQEriK5cjErob52FA6og4sj4coQ9QPpdYBPXuKMpYSslvbJ2WT9
m/9VQXmH+7Yb+IPun5pXIrJx+EmDXO2resNSqy7M1YVqHkAiJ3W1OZP4cx4rzdEOK16nyYGRZgyi
c+jcOy8D+kq4y1V00Z8kR+mTgahq5cgte6fEsIsgdxuF+Zc3RwqSfpXSyijAvwwKxio74iG2ECnt
aJK2mBYSBdV6jYVE8WmyaHkPR5X+aQSEsAgvcW/Vv69kMr07ofcgeFwSa/pejuWNvOz9G2IfC41W
dLlKOO0w+yAfZV8+ZiIx8F8dKM4T65FUmOEUWVMZ9/EKFifpbwFYKqeu4wImkJKbq9PdEA91kZYx
Ebl2bLD5cUCd6zU8M7gKqqnk/pjOCnnwqXo5C2wI7GKlbm8vc6z21IaXoikFUTQZ//T7VH+Rjr8O
GB7Bpwcw/37SFvjOnCGJdzdG3luzKsduexfRp66qESz0JJwVzmXKJJh+dhI5fWYYk3Hnk2Vy2iPB
FCpdMpURE5C5gWbMdN4p56ElZy/UmCn4HBr6faLMs8/h2xrcgWcKS0AeN9nDodmA5Lo8kBaYHkpT
lWr8PH5Q6Eax6zlBQNhFHI1REQtWFq5/+YyAUSeMNDOzfxEXVnBW5tZNdfAgoMDrwGJj3qqj2pMx
NKqBS98Y6tpXKttdKsW6rzsUE1uNn3QXo4OSrMms3jKJIv3OLZr35eNlkGAV3ePqi3liwUC+EXRH
uXnwzBWlREjsGsPq/FKOuuHCSs61xQimj23IJv007sDe8yGnB8qY0rq7+nnDGZL5lNARpUi22Cci
DnG7nWOLPgumHFEvvKMOt9kSjfCDWw8jMHWZfEv4+Z5nG2sXWt6m1RK1QVt8nhmbV0j0dwf6wiuW
W6MA9RCoPm02fZOU1iJCEzBoFz6bbtCC/F2LB9GM2TjFQh88ag7dTS5RW7iUDyU7XUlQa0dzzx2e
h8WizlsFex1xtWXD2AAhYfYnZ04f+HcEJUFTDUT7hkMwjcvGRE7EdReIgTF4F1BfBx17QD5KcBHy
SaytF1hMdmpJap2ZShdAVLFS3GM1DiLwPxuDaDQGBy0iUYNsJcHL3w1ZFKzNA7QPdEzpLy0ZVAjw
KNqJOWDww4kyu0YGv+F9FIPbokeXDrbHbu53tlnJj9rQDWuscNoUpK+UCoLeySMtuovNWemwpcHE
ofhTj3PM7ds/wwq6K/cp6GjnabTFFGhL2cUs+q+/JURc+OYum67DXr61kQSinP97FgFiKp1g47Wh
AA5yPWqBxzRnlGWL9Qv9UPEN97J+zkbcX/sSoj79ebJbSowVYsxKyJTEHJCCWPHE7ZHmYmscfj1W
txUlccEyHRvEtTi4dwuzcjISm8m0WSqfuGhBbHjOe+gQfPCr2OaE0mdtzd8OtqyCx3oseKNfJLVT
h1VlP7s5b+RQXGOqPgMXu0POfs9u/pQQIotpb7etXLQJa3DJkhiZqbSiLKFWhMmQKtaDf2jY2jvN
K90wK7zmUn39ocyICMX7o3JVQOgOqMykjda4gWKiwmxRZ/aYsE6wq0AdoUHNXCxx6pCPx98zu9ZC
g5AeBYhbddlVfEnMiMuhoONjE+vFFkWxymBOvn1/D0MwTish1u82cTp9dJIAPXssxLTR/I3wnP/C
aTOtpIcqD8BCwOBECI9F+lxR7I3ELlpREQ76ulHunEIc30gEpCINYl8NTvCbAkI7XL/4OSxU9IKo
+Qf2mmlb+UHgBFk/ZftD4yk/fRIpAn9r3NASP6AK5vTmtuuJ7tzSZxaXgPRTn49MUfu7gzDviARk
77a9YmJJC/F6ZvXptFwUxWL0yzNZQ0JE9Frcu1VQczIq7RPm5XIZ07FEXnyuJsVe2Q65EIe9bBBK
XCZgqX86af3GG3BWtuVrxvsZuDOfLz6rBHZs7WuL7ok9Amfum66/d26ad4/L99rgEf22AEZi/g9n
2VxyZUOZmD7EQ4x15YDVmtoJI531YW2gIZvfvB5KGQzjjIAZs4av15R9Tz5m5FqEF+BxFLZq/lO1
OuDjunnNSBnsp0vW/OsOUuKFhrS86z/6RrDlDmszF9ggjqZ7rC4k2hvVkkPso5ZNb9P3ZEn4f00L
wUFCWxRG+slrdbp8Fs+OOcYFtJn0VQjQDsmgrSHOig6qrQ9i3Yy6nP+RO8feBnZTbI5Qf+Zunipw
NH5bgoBDGOc7Wyr9+57/xg3eYhWJb/D9z3k8fRQC/bwnOa4R1Pk/N1a+axaVSjxBTXaUvRQV568Z
puBz1PxS1strS1iG5gwFfYIThipejCTLVm5SAkQfDu2S5mUcxHwl5PyBmoSJV65I67RZr/FWr0In
RnpSauPKT7vUrcK9VOgLBJUP9m+7mFrRTPphWPHVqYDS5R60fMNxwFcORexTvQSxEutBhAu3MMuX
Pyb/j5FoP5wEHTDFiYvlxS0NP6jzFaDE78sb1DdFFB+8s7sO0r/t3VC0pEaMlaAA8S031O9kXuqk
Za/6pXUGN6hGcSGkVne/XjMbjYGkLFXmvc3AN+omuVcklH8/LMWwArOohiw/jOm0fYRPXOLiFPj4
tN04ABHif88ZZH0Z9l5k1pCL/cdNPFSDE/L6MP6pTgpQUxZhgSQoislt1h8Buh/hdJfH77U8C3GR
xcotIK/8AczXnisK9iaGmkQX1uuVBY0NNiuJ1K0ANlA2GaMGqZcI37ntIfJGshnjiqL8C2aLwCcY
90Z7DWKq3rEorUq83ezvBzBE1UVcD15v2gXhDReP7RmIu/2EwN2aRZcUMD1xlYBs6Ui/WwB2Lz8J
Z+oOeidzkE2OQ1HqUoIZOIBp0mCUZvk2ROk5wZgqctWjfoTfDrZMWOYyHfYoQGv7VmX2iRZjlG/B
d3rVGzcqlnhvnWi64tgye11q0NXYbWh6rd/3I3zKDp2j+R0a8M0EGxMA9b9jfma91VTVtdJr/vzr
RJMR+aEj5ai6dio0RPOaiyZS7ojSt4nDxj7QvwulTAVtY9iyHSxt2acjqf17rWaS6ye5IZf9+T3W
Cc2ke8BwwOZ5QUXSbP6vp2Sg5Zlo6kDBiQ/sIMEm+dTbPIzNVp1StJx1A/slFqSlhxrCbp6Y5EdC
jl+rdAfXc6pbu/g7VfV+a4wbu0pR32FwA3ZLrxBcg2k9w+lCUYQ7pAlbBbAnC3YyYaF1TTLD8Fl6
vx9+btyloSQ+heF1YcPd9Cvzt1WYiPwRPMUm8xVqMqmQs/EtzNLUPgmUQB6pqkDoclxK88V5dp1z
r6UBrGf84fHMnL8DZ2+/N8DEw1Mp/On6AVrvOzxUxhl7ioF50snMycJjw3OUK2OCl+bM5EeLV0EX
htDBiWJ64D8oKiXB1JPJZo+tAv6apPN9fD4nwF/1Wv9XW8zF00mlAf+cnOzO7KRFz5uhk+8g6mUX
MP57bubSVBBwyH8DTmfxmyU5oPb5JbmNluQF+gj/6aTYCK92nyROh6kPSwmLL51BTw7IZdC9vCan
Tg3INuuIhTotcaYhUUKx3oURKYrl/RIzS2tjOa3rmDJkWv8mnLNOmCTDVGQyapeXmS0SUJz0ZSXl
iP8hDyK67oSRi9tCHL0/VzjqZNLpBqVhgxnW53nWTFDrZtz34pQatUCCu90ZpbEqfGR0p//UZf68
+Hp0m1XXrdhU0Iq+kuHyX2ZIfSMoD2GARwCUKNqVpsrq5Tnd73c9PuIqhbSyHP5qFgHBPCBlYt0S
lr3Yjb+kEfTvlnybloRMMYeG1ohw11wD2ZpUO8GLEkVT2gle2drlH/qGsW9Od/RTp35P+vZ60GsH
HyIZXwhiE+/jvq9E/bGDr6MP9qiglS6eBU9Sg7Swve8xNRTSsBXmMt1GZrNH51C1V2X6DmyelI9V
EkzLXZYqbk7WP3t8q1PO0yBZwnRXiYBz8ulsYapX6HM7OIvoarkXqzEWw2uaOT2sirjk+N+YFJ4D
QMqQcWy624S5a3yQ24XQqk+YyqHb2lTmCMEqOUPweTfvDuSm78GWQEBwY65yfCqghLmGYZWUTF76
CAXg9uOdQCBAEFDHcvFhf4M6B7Ju97qhu7sVPZGpfBZlp2yG9XBzBpyUL7yqrEi4AGMPNC1zX8d6
/LEZjunEfwOiLiK9/5FHujNGf8AG52j6xIQBZOEI2ghxcNf2U8G4G4nHrrtVHKKWTba2cYM2XQ9m
8qccQKEnki203TOpOiTY3jegyG11x7Zs6ahu4aa+c28c74JsAo0eF/m9MlCCfdjUZVL4N3/SlWTc
dyGF7G5CkQK1Y7QaLghWECNLaKr6Tec5P33MNm0KQvVpnpFfi4orJIYyQF9dxbIKvjXjlITbhCMh
fZW6jeCuiQNIgd/tGnGSOpPRelyY9A745dV9zdu8z42CMvqr0O5fbhoR4pwxCfGdQfXWvtyzstU+
xNqT12+iwH6rMv6de9Hi3EmU0YhZEDjtmPAALDxFLj8phs0HwFNKe7cKWm5g5LbriY//c6aX5x0a
gRedHlShGYFclcEBTwygDPUVALiNJKpWC4ITYuezJyEYgQVc431xaBWmHATO7NUENdbPBucoqmXh
PIe8VsqFiO+WXZVYlvqpr08OGnBKOXlMw3n6xXdyz+OL8GJSrIGYk2DK4ZOC0OEIKaNW01nthNte
WwoRy+efOHWmr3ZXKmNNihHZSaAWhfWb8H08V2NRZ0RKrXAywmvmiYgfFpATtTwVynTI5YRkGIlP
5PP9wlv7WgMK6kAnQVvZcnJtZN61ZQEQvnkHpHHPH/bAjp2QmQ8Fq27avYn0IYtM++EUoCwDSbjC
SmXOsfHnE4bCCMGvbvGItecpPKOrb+oBTKxEPTqetwwH7t4QqGYwqT05a4CTnsBQqAqIuvOuXA1T
whRdygElgiY89PLqxnZsZf9ARDbT7nnfjbd42WYMQO1TmiFQyOBMH0Cn+VVuVjciXgG7al+SdU4K
X8SkGt1LCdHOcMFcH0D3GY0Q3PYwtKaN1e8At4xZhAv8mTPijIiHMEnkeiCObQJ2U8XTPAcdEECr
cv4hUcylu+fsQYmsTDUE+LKvUZiQWLWu/E5BVBZ0ozJaXxTwwtrAOiVQAi6Cvbyvbc89tXGGU76o
mJP9dhyxGL7OUOaH0CAKgdDpqGdxhlzFTE94L/Tsk6MVEbsXSVW7CY8Z1MQRZFLARg/gluhN2wbH
sp28uWzyJchoYdbJkq+yQqyfc/EMZQRvOSDkpOapDc3VJrX2EfAHe9q39ta5QSxH14SHHZZah4O+
xbyyDIzOV3f/Si96Tn+V0q1JUiD+XQCxQOWsHgk1f61z9IUfbsFQjQEUdd+QWT6qXEWbXC7b90hh
mS6GZBBkIXTEPH2KNOToi/2F/7wRfP9liaGxnqp9ZsLPGhDRZwmSY6nAhCYuG4U+VBJtNGIGFeev
4f+wSy31v6cjcEUHn/m/AdP1ZlI2NiqYrNxnT9UqXuZn0YaSQBeqd/JqwOb586RyHCkOLRAvlw/A
qEuDza81Cut8hYcygEQEbHaF3CUq18l1sblseYsHyWny8CspCInYkF4GrHu7tHUMh1HHeIRg2KCT
SD+Ug1VY+Xo7wHNG3s5zpBzvvXEGVatFcuAozb+Xa9QtC6JYUxUHLKn7Knwq/4bW5tnvvfw0W2JF
V6z9e7c4sAJzBt59scyzpGFOZ0N+4Cf2dsZ17zN4X8v4SEkWPC5pfbzJJsUt5oN4UA0fLUvOzYL2
+WN0tEUvCpsB3wxvHQZSAqE3yiZetADJ7SoDMp6cocodu9/OlHpxZxymH0SC/uSOHOkdwPT28vdr
IWVQ434qS94CpyeajulH44IGPlEHKuHEGqx1ZCz1vgiQqudlsPxtbdwGxLXF2e4U3FBplRokg7Yr
xJT9a0CaDQvJERYx71bd4VObq0meU9OetxYfj5JVruzoUfVBVBW/NXFhEdaURUYRwGkzlc3jrsq+
xOePkC2aCVTWSFPaTySDtUOcgmPGM3mnLJaqjxIv22YOa7KITfs4SvhArpgZKYST5+DCjjsW7lZ7
DHN6JKV1OOh9BwBZy/ARnR1om/KXCnFNQRHXKOK/6kkVN/F08Kl14lkYsnbAufhWPQ6N/6G5N8ee
IFcCHgB09HlhXvDrg0FeAzkUJugDZyzk9LfSKpHXLp9Zf/PlfuGoRsplleh5ypEkLx6i2wDvskVH
ble0F19UhjzxCbZk2JY+1KRgJvEvwNxgd731obHcwjWBgx93i6BMPnBAYuF3iLyelfJDxU0sBl6t
nlf7JXMScKowYPW0xa5AsqFy/BM60k7Z8rFtnaDknM0sbL0Cgb23CrXd6mx3aB5/msS6BlU7d7Sz
ECEd4iQBj3f5FP+izhC/BXybM45ghWV4Ub5xNG6RTi802rbWQ187Bcc19PYzWVIk3wcTQpNWhQiX
k2wPiE2gLyCSnN0nanzSuBkLfbnqRTb1MNtIogyQQnTMo82yeP02dnCohvC577Uq7NeRzX/iaIWp
7D1JFbpCcpXSHrQdAcq950zRN4jeYBcALx1wHofwozvPBIcfuA1CgrQByY+tP9l7745SJHUpHQaC
VV4z33+4BpaqiUoDlBnt3SwjFbUiwmAnOP3vv2v0Led6Vu2lmoSvIkdoYl430UEC7kCZgLe7gfCG
tCrUgv4iPbSEvu7g6TBinud7kZvGryJ4hccaFwiFXm5s87jsTB8m+v8udEzP1hj2ByJiK28JoDw2
TuQYMHteRnZzoUy+uPStiantmOe7NvHZRArqB2VPqM10yxR8u7Kv2YBY8IYF3kesrOx35OnLc2HE
QdbS/i26J+HtVgPB2LGUGjCGM8tCFRYcnMJ+esY9m7hTCaV0RTRoqtHgRsyJ30hicJ/xdTCd9Jgk
m6iVVyWWIhRcPQNyOdMvNOaSgQjAofZrGSue9A4udVf2I3pq3yvHCF3ejgA7BlH2g/Oyigi1LSVK
YdPddaodB7l+SQ75WPE2cEtSM/9pn91hmcEIGDC/HFSsTwUoZkg7I32+AzVrWEgaBIYhWRsp+Bt0
NHnbF609AHzt8Nflo3uddOArDS21CCIQOOeaoHnn9dbFGiJWQzvpdo0ut3jplTX4N/tIsSQraPQb
GRybl5SLdPdNMR3aPEUEMdgFcw3vbE2p814CR5EEYb/6gResNMiHM4Z8YMY2MwLD8a9flRQ6j5kT
tt7O8IDDMgHwAhZR4tWGScDzEg8EarcmYf94jLlaLWYTvgIJ1yteNMBaqyzedUUr1rtd53itAyxP
BhpxwXWCQnueX3pkxaLMo6uNOpCC4gxm5Wu2wM9q5AatS13tBVN9E8VegqOGCn+s2ti0fE68JnXQ
Jf6TVkR9tPsBSYsjXXCb3iTqr+jJwkKKp8pVi7Z62NhTcTwmlBDdVAntXtSFjbL4/HNI2LvhJ9nV
w22mSV+cDe1wXbfZe31EBSzkmecAVjMdtIDgoAnSTBaXvTGpyEN/rFG6KDLUACBjNhBFk2K+pBKc
vwXFPZcEM1owicBQqr03F/NB0vGaZBACkL1ACLizen8X14KftL94ZJkPKlBd2cxCgqfNZdOsDJH7
9Qvfv8LWfM1PK7Za0fmxfBwhkoZol0J6GGejqVBeb0sNg8ED4vMbrZ9FnRy5hvNR3fKLR0YnCoga
gw8jQjX+epjibe3oRegTMdxoNMsJGspRTRY4lVV3pU2ojxoMUY0sH70ixVCFlDCOJrlS01I0fiNC
9PEoeChOp3z5Q8iSkRfMLNvLhouovl3hchFoDmHWNoeZvIlNNve5gMwWTjR0DJ+5I66da4OTDcE2
PveGgOHfAfZqrdf33rzAo3b0n+PSJHjVML+qtSRnds0o7e5SXQPMF7f6PwnZruGGYpBIGmiHZxBe
wWVW3IaNsCLgx/NvPCJbB0BLQn0O/6DfQl26G3bpM8NxK+TSQpRF7Xyw1PrBDb8BGIeBXuiop/fI
/XLtxfnx5+3drtrZdtzzdwIms+Gu/ZnJtLu9Bl0NHPanCeqq6xt9sXVpP/ax8rKQNmgcVYLdvSs7
oOuJDGZtNB5e33pr+MijDVVfP3HWfGa6cWZ8XJJtX+3ZknsDOB/HvHrM0GB9RX1Djo2HlBWczzFb
TAUWI4L4VQuaMd6FjOvVimV9e09tFg8dAZI0qFk7tXlEc+fk3xrvGbOPdYbbLwP10/rCtHqEu4jb
PbS8kSsRY2SxMz/dwafD+8flWw4L3Kd8XdycHuR2+MGwVChd2Jq/XAIeEOZpc1DpMRPYSWGsBVYr
crvfVhedg7KQFAcqM8Lydwi/BS4vm8yYqpTmPl8v/j2A7CFMUlailWLxbqT537RINGSpt+5dcPYy
ZCT6hhK4EGxBT7l4IHtJB5YgZ3Hvg3ZZ195KQLOKDz8fKG8xJF7KHq3j7cUp+8AVAT+tIX6C3Yp7
59zyTwvPNcmiYICwMpiBN38NRF3/yW+O44EjzTScC08oZtHyWG4CFR+d4f3sMzzFVm3jOw26vbzu
+r8abs2t3ZSEn0fw7HcpyLIMZ51U2oFD7ozeW9cv5T8Be2id8+6eJd2U2H9pQFe95TlpQHk3iaIn
Wp3/k0Zbp2YOTCMmoB6cDQq/NfHN+/8/g583MmLtCZEG82iFDKIyd5hWU3HIyVp9XTmV8tGVq2fS
vsgLPcdb+uBdmh9YJ8YFLW3U6wyu2CaPwWtHN1ARXiDreEsTCoUhBUn/IkJRyceCwzLI3yjaGTOy
D9AyCAcrkQEMJsBXLgTPOTZrWb3K4r9Uz8v0hmh6pY46CuycAgJ6Z40f+wzHneB+xcVsTk1tcFyz
0pGpvmPytLwqbGjkTF3dOx1Un5xu0Kxpf/pzzmBprJzhtV/sZPeXJgdpjr0ArKaRfdxdinCmNTSY
OOt6voyXsbbEFouFvjdHfCJhZZ8mZgJwGm7jS3IYtAn12vdskH+fMTDgkX77OwjpN7YxXy8nkKJO
rw0kggN1/Q5AyWdLAOsEAiWhstOe6+r4nKgYBXePKTTv1cZCDapjMtC9RuM2wl5dpSEUcFaY5Wjx
yeC+Ee29gsfMNWRn5rBQgCjnLCl9OAwYYP36hyg25FeEKRYX8mRL361jdLgCKIJex8iqxXloEACq
BBS+BC/ZAxx/OO02t96b0ukPA3qzvOBR/JEe0hHP5gDAfb31dKYYnYJEAyHSZVZR3nE0DVHl/SYi
8MwIqDnKdJMKoFFA8X87eTY05lv0ULOFGuMaeVNHxZuVmpN2pNHLczuAa1cx2H2iMLNLXeeccxLl
Swl/Dkdiemn4dPlqZL2iPOZI/HN2PHhzehAIeNe4Wzp686zU8n68NniCvWaMulXtKYvuXz9C1nV0
lX44UtkYiJ6t74W6NZmsO7WlxeaWNRipkaaZHKL5xhpw51ESr3w9hHq/WxI0lxX5yCyHJYrk18gb
ByoGGyXg+zCi187X9DIilsBUeLZiFIwLuBjRgHFqrXbOI3BNF1sIMiE6rF9qUka7q387MAgtQRm0
eYnwr1tGWnRNXIF8loWHZpDz9taU5qQlYEvbUoxnOVd7NjYec9x78WE5VMqG03k5JNRtOMb+UHBJ
bweUyXbXUMmIiY00ei2vtaY+6D+c4x9lXIrS/wylNbqixoFfaz2z/54pgrJ5l4kKNnTnwJo/XcZd
a09/3XOzzE9hvXtc5SVoqiOxmlMYhhH2msNfpPEb8ZlQI8iGCgSLQw53x3eLtRR/WacYFxY+m1wW
dVmmbJcCa0kPxSsHQaz1PtaA/uv2etWX9fdmZCO3a4NdrIdPkKjPUK0GCKZ0m61WnffZfpsFCYLz
bsxcptb8XgTAA+EDQXm0f7ZwNrJeawfwJu+6qiDeGxSdjGIuS1ytkO3v0viNuMbgUW21aPzfdov0
txMASgnYbpq6CoIukCv62VfEGUh+inXWx/9d6dssSh5/lLr+PRwKyrrPKQupC2X1jfxB4syUK9+x
XhaL22Aa0omLFoAoCVghV2xk70YZl0YtY4sjRjntio9IE2F7tW+3pHhF/qYOlqIPIWe3qXC7nTGX
O1InsgEBEko+nrpt5o5TjcdXeuTpp5oSu1s/toLbkEq/9GGyLqfD6HIWfJu5sic4oSpm1xfvEh8H
bW3Kj6Th08LrAB5swLyJXA0/PJMSxn69JKNw4NoHGVs96ati37lEVRWmwvxA2qpq4iB28hs/4P2w
87WEK9QQqd1KG5e05+mIlJnY6plMjkMebsj4s1VAavYue8pP5gIISYEoXO9/2INBO28tnF43eNg+
cY63iPiki8Pd9T70rk3dMcJjPoOb6shvxat3aWBt+a5OSGy0wYb0SoslJ9quHt1sI6Fn8a1i1J+6
2smMQBxvFN/AHQKpjXnJ2PZxgI11llHBqSAZMjAGGbEeyKEkFt90xLbjYm3R7pCuRtuUjRMMRoBg
AsX9hRlhDBwSHLFRsyExcpnVj/7lNHLu1VhleXwfFvLxXWYRNc3MyQqU6QLMBKJioMxPVU0sKkcS
27IuLCkoIXDNBHQJu0KZMox1tOYDYJ4aCIF0L5TNJv8gmmo1Gokl8r5MolujeesfX4jjWFNv4qgq
vX/TUu7PXkrfwZarzENyzi0n4woNDEolla+f3WZgddlohAaFYn3jBIcSpFv09rjWObdrVSJCEdQ7
avhEBkrV9euvmnpxp9z1BgK99g+U7gHa/Peyb2dtNTaLvpG6SOp4x6iVX7wYi0j1mVhCVi9uq0Ws
u4IneA3OPHSzZ5MmBYVYJwn+Q4ksL0lerELRbvEtmbwdgc3h1gVPW08ZZln4O+5k0et9kotw/oPI
vr34I3s3099O5HtXttBLXV+O4nTeK46MVOzcfJ+UgwVzHBOsYlFB5tCUyJG+NgQR4juo/fXkqgHR
XJThed19HgJwcmbFLU8mFL51qIUzL/REvcCyartmW0PREUEq5Qmr3dL/AW1Cl/zHq8RW931Ewwl0
RuF3QBE8JtPEWAs+PhMSo7k5fy81fXmGmnDNbILxBH5hsFIaBoeHp7vGUbujHNHQP6E8kXzy26K0
zTZb4qrSsVKB8byfI2sQO45SwLmqNnNcpmLMTsuve+/3k+ez6YuRRPcOpmMz5wK4Py5QDeRToxIl
CdgGa71R/GcvmgnNfKBZqOl1/FMUO+QYQ5Po4Hunyog/Q6FT1AeaTr8PmgFK/hRmGEMM/48UO7Ph
EMYWUR6thIPa5GMdlmyK0WF7glQGUf9bSZaL8R2rhrUDciADtIJaAx6+/68j9pqujzFK7dgnEn+r
gNhmCYOCWOjgx/0/4uGfjhSo/IT9kmPUzLHcUcSjxwiVDLhdjZ67YZM4yPlnQcVYCgnmVtjxnMHq
qmOX40xfZQ6pgnu9X9ykKG55KqGntlAnGsdRvsK7wW1IRx2GWC2SfjvAxWBrcvrZUEy8YGjnI31c
S/VQkx2TjJp+iIXn8ClbjYHcjob/xXaM4b++ShQEFc/ggw3OvWTEItW1VCjjFxtDAyQpi6Eh1LZT
vzG4biycqWyzbVEYRSb1YcDQFJVBRwKVnTCLE3bLVlp4epk3MQ190q+GStkQ5jCpj4g7sXv58zgs
pEWw+w9Jx99zjHQYNu7NObhIkq5DFuz+upgyL9iwybfENqJpQ0QSAPM6TYNdSA03GmL+lpA3aINc
xBi42/dczRwZb0gqZ01rbMcoP47i4/9AdDi4wuy18mSVJJmzc+G4Smr4ebT4+Qv5ntfsiEeNmIb/
9LYiQyVo5HUlemvlNuBdSuGwvXXdFj8OlaOs6sfjhEf6I7CjbMXaWq9kSCrfYxUUnXoVQ368xV9h
69Z7ebmSFk+fvqB3YkmZZZKtscmrR/mgmqJ99OIdvRrSmf+vCAw6u1RRvT6BkUWKYeLJO/+EeFdp
ljkJpx5zUBkfrAydS45ZyXB68YAUcb3P5A33OqcG5gHbksi4A0Bkp8YtqiF3Jt1k15jO+tLFYwA1
8FKg/SN3wXTanjXnfosmeB8wZiH7raz1pLiI2gbwbsHVwnFN9B5WebiOrCa7EmCxFMfUSsxrELpQ
BDRQOa8znl2bsd+sk+XUwR6bFi5qTbY0a2QG/F0t5DPIAf4aANpBpJqVeXKGtGeTjoBZwbDSooXw
XhzOa+hTItOd6E9oYCXbPyNPrwbedbGDmQjx3xlzf9usmmNItV63qjqWaNvvnK4vFj16/NyUSKXz
p9VnOsYu/4LXc8rVxUjKNr1S3gZhfZVOWDeJrKINslTOSWDsa6H9viVgBZD7FtNSxHEvyRBlVbe3
qq3+eoTk6SU12++LmkRcSXHEMJ45Sx7UPjtC5HQbya4JgEeEtrmoFBzrkD444egqFsUX6lse93eJ
56XKh/0tudsfdCcClDpb419nfp0B/7N/H20X4+ll25YDJRXUmmZLPMwKBsFJSs7dznEHtyYLw1Zu
SBhKbE06c1AP5w9hWjLyu9t2tZoR+IzZTFbCpRB6XEeO81koUpKxKjEPeAHZ43oSJIBbSFP8np6M
V87vssgiecyTNvOqTOhhG8sDP88SFOBRi2frBzykbU7KRm8zlesldTeoLPCoDmJKjG++S3q7/Sfc
2Wd4s3Up4TJFEAKjemilBaijbFXFiBH+3JAxfjHIisQCeBpA27AN4WyP6hIYuAw16IRK1RrQFb1m
ybaF7zMFXsQNKgyobX4GsVwdV0u5GDwizSm/+bRd4AuvtaGkuUovmIRf+PxUtl8sKTQmp9rJmTpK
eeu1uH38MgQv+tOca9cOj9qfxHn8nkISWJlFvJyDQuT7N5A63294wlYHM+WHqtH6qhii3tCjrLMR
43/HNrfzM8r+bIokJc4yM9c0zti5+RNiPWSb61JnTQp+D8JjbjaIr4kOGz+IUUUzA+aLbILUV9eV
lOFpG3wb91XgaFm/s/uUJNmEjr4awLjOBlwDJa7O7SW4LhqhszcD0de8aWeUCSSx7QHgKT+csUiz
ychPVtTzE5HIJ1IHSfxPD4Tt3pAk0l8U6940BDW6EBe8MdDrLhqL+xcMEkgmX17WKZyyFBrwnkzu
yJldI76zduwmfFUvIqghG4MzOZfjgPWOi0kZzQSff7QmIPzK/eTxmRt/ssUEz4Xhjqg6UMmxLIIM
r7ysB1g9lODKAniEmyJ9cqQAKGrFfYgUXNoL+VSJxtCHxCWysq07QJJYUh9hMHeUxcK6DQUDTnqX
qdhMYs9nVgftij1UgtKmk4wp+bCMZBpi/sEN8ShAPs/Vp+87AOUG2YWFtpOHkgzNIO9DOZ8AGbyP
GRwFxqOsp6bKI3QShUMUsYwFW35lz7Bg/ptBJPLd81ijKtH+LT1DmBq9RkpEIXsSQIuO+iqggJq/
lW7QmNkJDgQAcl+XpHOUmUVkvVmBkP7jHYMn4ZPTf/Y8efLfrVM3cGonrASftbcyWyP67SIt6X6w
ilqx9Cv7h2Lu4uXX25CEiy6C372v1UE+HzQyKgzoC97MytaKBV8JDyLiakP+jdxHoFfiIyx+IqSU
bPY2arsO4c1bCzWfY3115qOfTmhgxTPzwYKU1cQaHCDt7MM21dMsfTdqTkRxRm+2Qh1/4EprfXtT
kDW4R5rhINa8YMcXJTeoiSCLK/olsFPet8xAAk2SCtnAHeRnfFWjzk+4E3DSAIrNY2ycn28vhTIE
bJasqzE4gNGjCLPLG2gtC4+9LgAsIueZ2snRIJWLkd2GdolcjilWcnwPuQeD8sJOW4fdlKfy+7RF
g0sFslOPCcU9/vwvy+dHopIQ7tI5b6hHCeptodwRvM6qzfaJTSjC8G0e7q8Ibnj/1vkEgytba4Pc
9tkJ2yvnoHepw/+kMGFe+H2oHabxleH1w/3gfGgxuGJXuzk73vmH7YjSFrsQBew5y6OnvkwFIU+X
aho4c/QN2qhjjYFnEoXfuI0M3I7FXQFuVDO9j6dwX/YKcvhgulr610R2q0v5H1fmBszTvgoIFqeY
ZeEAdqYLb3iOdgRUX6Agd3BG15t4LJ+Idedkd3FWbOaVMS/AvQNcPL3QE6YyBhUlkaZLnNYQaMzw
TguJGbdpDd3KYYprAvS03jnz+ve99awuihij46DGFQJPf/WuCKQ3nf97SLFMM+S5xPa7fTOQ9W/i
nVyq6QMaqnmGMg3VSitEx9LiSdK9hv5msoImISJ5wyZwtUYFCbBmYBZ5ZJjyTknfV8FRGNoig7u7
piLDhMDCQo4cn2lz0GzWR1X0QgNOZGqeaMyRN2BZwpmfCyb3pMpk6MBbyZUmZCHmdbj+ZIUvv5ra
n/VMUjv4oEPVXqnCIzf6mOH+GuQz1J4NrfM9+9LhvpVs/VYwG4CJbiYMoDcy6SpR3LcpuJQMAskk
AzS2cSqdm9zCJg3Pf/fuzVg9FQSlW8TZeMLskopVWUNdP/gzqAMfsszjAc9f2SKZ/lig8C2HA5UN
7/yhrzBmkJD5j6+l5YZEV0JL0MjEQy5Oa31oP6AmFPOQRKSlu5QrIRhjl19CJ6Rio3HpAtxkUbKt
HjDLJlwXct49B9UyvkECmpVqqTQz+FT3IyyCnShOEbv2ntDmca3pCjSkI0ag7EzDpOgmxaOrGqlE
BYAys4raoJmGof+zevcSssoBHUBrrf2TpZB+PW1IHr/ir5rdN4XTTqwb+jSTxGI8RZNt+F8O0pzZ
PF50q9ywaUlfVs3Z0qOZpvHWYr+ZLJZJflmXJrXSiMj/g79WWwM/OCbVhXWAgxbxMt69WbJhpGzu
HXqYxOAmERdgYCd5aEG8lGAmvxhUaRCjv610DutVMt2Kaj8PaTosK5E8YwlRu4Myslbz5Z8QLpnt
fd5gHaRbhhxa7SkD6JidOtmZ7LuGsjHQh1nBaO+jjbhVWJ/5p29PxWW+8SMjCbBjesoYlMAGcus8
OOuOIhyvEIubJjPM214IyaqFBEJAZh9K/T5dzqJNNzZiC8sqs1zdPD5dRR7pleyaN5SpYgXYgeh+
DDlmuSeM3XGqIs7IujSHJQunBFEYx7C9kvfekCnDGcZQIwmUknQXAD8kruVyyEpNS73irLVOj0QH
xoiZll+F2ETFwCQofJlaAf9qlcVFiR0rtEr7UCtghe2sd+U+SSVt5dQjKUVoAkAtuPJn+hB9PSnJ
HJkPhZXE1SlnFRKRqtBYxu6nkIiNJ1OdUbV70LYvOwucPOdXQYONtgSYgqQ0cwt8v2M6WBxjZYVr
ifhCyIkCipm0frYLnecIlvcVOBOBDuMaSieWZlzfwN8ldcVhJfzA28lUD2zq6pWRfboe9BIVAJaT
+7tRe7cJpgYjU9iOgCzm7Stj+WoYsMWwPCOEB/vUxrvRC5TEti8ZBEhA+xOMOfTG3IYX+deKcttI
W8vTqatJgFN6FuZy++qArClTpSyjNZ5a41fVM/BSb7sLxtNKe5MvPOZQyTSEsMWXPbyV9mrCGWL9
NSedtvNT99cGr3ZUQsG36kTj2Wj05hiYW2q5igzOg8fMTDiCO37iao48J+PTivTTYFWJztr2Dg83
aTEtKFkS2zgXy19s+AoPvbXYObHGEOov7sGjS+NCmbiLCn3DB592V0MHPI4kLWOlG2lJGQ35vB5j
dxUZ1KQKgOcMV1DwOheA9kZqXJGKTj8Y5lDO48D13ZLVJUYi7/hRFkVP6TbJeBW1sM9nOJZI7F1A
DeqLS42i6aC9ua/wnUsJxR0ih33vt8elQLl0S/y7bAdxfPYZ34lDDnJSAEh3jNspc7LoUfcxcjRG
8nYuHGba9/OwBDgsB0wXsZfvRYqgovJjKFVmAwAV9XjwLg4sXmPfR2eHFEuEcVW+ycIfIUgNq4t0
eOB1O9plsRmlZBLJg/nbmXzOQhqRt6VBef1nodvY899XWgcb8umsrZagoQk8kXqsyB1FWhnl+nW0
/gtDikusCiyg7jrC5ENnXNKmr4P/02Z5UorfHdJ6mcPGWgd6FyHwtfuCeOJ/wtCrXHTHozFgZKSd
To4grROcoAHHGG1BvhWoUhJ4bEEsZsyJkZcHhcnzZyEHaNSkOIWrnXtvXozcnUSSiw+aJaD4PdaK
7HQ/3ejQCjig375HXKToxl6dOL9eUuRPIxXtA9UPJyW5yYoZnhCkaEMpX3I1qPqLlCUXYH5C7SwH
yDjvotoNo06sIYY6RIQBy5MZ6CM8RnYIgNoD2zKULrtITwkOaUcoS/4annlFKQJLsG6Iu0+ZwoHl
Y/oj2qQYODn6du7jFNe8XZ4oduVz8SA08a7m5EgC/fwurPWIZaSZIbleQVyaBCWpa/K45ltgC3c6
egyxOuILz4kLhWuHwVUDKYOL0Gm+tnWm2WEtP2DJyAqL9OECB42tg9GVuSxEEuUMDXQckVqAQnKN
xru5nXWt2oXWRW/smPgTBKlcREc3vAuN0zvu0hr712zngYhaNGbnLQds/g2MAOdMPPiWHM3G3tkC
qR3IDOLND8gsTrz9rUML0ExEAxn2qo7/xhVxko51KgcXFyJ62Tha6GWkXEoaG/LmuxFzkmFKn+Ee
2tAIGGnrUiF+7puzZculpLXgsAxykXNOo6QhyKX9l1syUjy8AOuYejqVeIbwXFF6yHFodUWTUIPk
zab9Uo5W//EGXpn8ZQZe0AQ8zSHzQcnPlw14BCimNygUJ3E1zIEmW+j/X2cXdDA22QX0NOtPjsgW
FFjja3pCiDJ/l6RhMWzbH0VSw1z09LgqL+RDrazMNHCFY0mMRQ+qQFk3ZisIpiLix6wByLPG9Qgr
ZOWYpK6QV8qZzDiu5lAvxFWJ21ybnin0aTYJOX6fybyCVURLYLePxHqYNFI4qB/yiYjX7oetQpTT
QT3Znt97gruttLRnGdUdY2YBwo5A2CyfY3dOnqts7AiYtE/0apwlzXPa2hAzlQGaGw70g3YmKKRe
hu5bSIGPhp9z912TwRGjWRJttYsyc0M7gOEn6G2fBxpR71+IDeHg4jPLPFp4ROj7IghdgOcliXps
A/p1damB4D9nslkmg+k3Gnpobdm4z3OjMVIYOC//iTd8iVLjfDIhGsE5Y63nW9Xo9sUcpgen9MI+
XWA/HEVcK2WE5l0U2hMxuznruXfRjeE3L5Rc+jHZCNBkV+z7PPgpZPpFoxWfhPT5/WAgOFMfn0wy
XpAeUU2WaNcl1ehNdGtDvp1iEsjEIE6XA5qCnX9/GD+IjGrUkA0yWk739ahoX5ZLleQSR/wYaQSk
HHGwXoCZMEk6nxCeBEaytNT/SvPHQPHUVL6oA5ykn8rzEcItzXFBpUW5DH57QYBRXFb1s7Gc2S9U
Igbb5BVLXJD6IY6Wg9tiEbzUUt5T/y8h3dKSIBYQ1tIKjY/IK/8a6CiA2GtMGM0IyL7/WxOHIJ84
amIv41poM/yC4xEoQmvnChUgNRhTfFUOzi9kEWFQhjELX12RDkrduD8nPSNRAK5SbxCz4YyQNccd
a1UwbbS55KsKqTxKK2YTlPyR2OyGTWZnAEfAMJcRrIflo2jF6k76gUXT7xagCXbc9sRjxUNEUTLJ
SkPH5PaYKqs0U4GDRO+DNJb0Buv9V3bgNvCR9gclYtNIuOkMWsGFTbKooqZuxLBM7Sljs+SXsfgM
6E05L9mE1Yx7FrHkjooUpQWqEnozvUWdUtTzbYxFMzSydsMQSTe6Iz5eF+84rK3UJK03iukn9Plc
xsIXKW8M4yjgY9Th0S+TcteluilLzlVa0jA1T/HrpPAhIzFv766BwqKjj12aLhVP1Oico+wkrehI
Do6s8IARp06URHsxLnbrOcc+qjcmM9RqmqXyJSrHNgpefe2bYcfqgZI8SY5rjVnnrLTeLuU1UYlJ
t2U6v8bhwJePpeb8JoXwvB3xyHgT53f+WX437w927/Z6KYdwddohVU1FxA0HqVqeK7rM7mSnWyzp
LwlynTyiJLhoFVCqJFDNGNkbXjwk2OoaxkDQSc4Isz2ncenl5sLLqE7qXXXudgrUVp4V/Y3F28/1
0TwY7qVXC4HBhaeYRdNGk8E3mC3HugAh8QdwTry8ZDGUaTyNvTaUcfOabKikV1mQ4EL1zgot2O5x
XVEnFreDoKI4RBptR0xH4yvWZvIjkQDpwLAMgFOWpWcVrAUCsIFm/R1Wv7zwff8HRBs98tMVJEUx
8IOBP4lthgg4cKIxUmbvRucDraKce6Q1DPNvpH2w8VuCGqy56gguY3q90yXfiJqUBj7ICQjjIym1
/93AS4i7kSLhrdYYaIBJfPdOYBhufwh5jGNiRYtnJH0KkdE/XHfZiRa3TSQnZf38GL8KDnYnxxJP
RodgbH8tLt/gD9N7juc9uQJikPVCiyMQ3VMMlJkpRB2LMErn2BRoz3Kx1eBfEpbmRmQtqU/wp2qO
tZmWjU2Its7CtaH04BkIHCVlEr4cGFVCvrjEZj9O5sbpeQPf0XaqCNfeSsR/nRvvBN72hVOV+gmw
nuGLdyAlZk/+KW1H2XS33emCDjUjCFvqh18OQM8k+1oPpq8jz6YcEnLhH7bHotxw+ctkA4CVcTPl
+OVtEGi5r+3AeEflg03GiuXycxTa11HZw+B+zVPY3fbv6wrESJ8Htqgwi8UUhxNX3rbVqQGadUjW
/dudwpqSavluM132n752tKnSDuyuKFSvTPf8oNQGW7d0p3B6HTcUfrW/Abx+nDXA4JxWCBmUyNNM
/9f5sbfwJK/KdkG7KTrpBH4e1KibwSaKRfCwiWOr/9oGHVj2brAhNNfW+X5tsVXOBpJdXjiMVxob
pC77I/VseRFkX46Ei1LtK7NL+tfOSbspmcwK2GtyeEdYZGmnNz68ZnYYhrLgoftdwWWhWK5tA2m0
OR0Rp8y+mp8C807KwTh7DMKIezfe+Pd+MyQlm8LO2xBF1jZNyRIxU55V964wyWj5voKtIfhDInDt
peyj1EHitmikFWgT3Saa0o7HIFEghxrxdmB+GZkR+by87gxaeIY4hDIlH2XW51EBho2YKlYbyxaA
9zcErlm0Mz00dTqcp/JVk8PhBRPKldlws/hnK1pHizpp8URhZSqDozLNZzCo2DiPEj0Tmha6lUC8
/FtfqbiqhLkd+MmiXtI5CWKT1qNlSTuUh/cGkgptPpMvwiDYJcjsAuM392PdQ2gDX2gfY9ehwQ6F
QW3VDpic1Z/+olQ3QDvObMi4K9gU4HZr03niVwMwp/gHgS80HD2RMgfVSiwvj7Z0zdVIZBIw/6NK
XjkZdSQYW0ZAyP74pRJuHbTdwkiqrqaMzYeA76WWfIDkDLheFXrMvl0m20NPPtfG188qQ4lCSCZQ
34xHA0NmQH585/MQiT5htlN/m502fUb7WpjZ6IDCCXa9rAUlXFs5/oLFjgKvFNcz2kWOvV1FPECw
T93wSO8tu4Z8MSU/8s5u+sPckU785iqjjm4AfCNIxUZOydPY/r6FMxIGt+2VgKzt8EmghgE4be2z
KaPqGyzpEkCIA7r6K3wTXSIfUHb0vUP5vfrWeHFswMFaiDN75XHjJjHDRQTwpbnH54azceYrokH0
qsiObgnvgqKKVskilul3fAz//pwWSR00RZsP5MJs2UvnCvAUpIdaUZOfIJBX47XdshIj4A2gxuPI
iG+/pL/rOiZxmK4saCkbLZ2c1weFZC3RoreUo/33h2XzKRFAOIocnEsN651+gnSH2Z+sBj/bwCTl
TpqwrMB1nrGaxBHs7zweogM/TG277Hk+naerEQS+9pXHoRM8v4nLOb/I+MSKVSgt9VtnVosSiIK4
mO9LuaPvxf0T4QGTHCh1JH2w5Z50W+yb6zlF/VE2Thg0JE17enqD/AJWMz67MeOvty5AaW3oQryh
r+zquzL+6BaAa0nxN4ZO10lDXUiYKvEloT8LfnP/ccO21CXwlQf8UVKHYWsggkA9F+782gO+nhxI
ZzSzUJp2kptwh+7SWcrR8SmGWRWyz3xb9qP6qkPiLCXfpWPAuXINECtpPiyiTqo1q/rQRWpniktp
VOdPvcoYqSazrk3qvjGDhYxuqwh0ODYT6iiZ+MxyYTrT9m21GBodXopDc5W1SVm/EBLxNdc0WFu1
FV+wC92a0AJWevIHQ1U0I7gv+INOnOZ3sEODP29i/UAA7BM5Sl638RnOXR/8wf+fFoSQbeSjjv30
1DGpigheqaJvN14A+y7AkWnTrjtFeJxXqhPCYyem5i3tpCjgZBLjwWBT8ANIS5FHNGF7O8wvUiQO
tQDNaBd0hwDv3mdXH9XdEkGnvnXrTkXHCa7fxrYc+4TF3TZcxSv0mF/934awdNCtPf+DD7V2FyEf
fcl79Gkv9uzTKvFkybLiDxT7U+MySVTYdU5JOZo0wr7vynU7R/Pip/0jE4fT8/abpD/3CG5CtkKX
DBf2tPXSJ/HsUBEFPm3QgyAnTRK4u5WU/IjdV7P2pcGF/E7z7yY3SReZD77CihTNs6Qv5alA6n7p
ljOtdl4S21ptOc3a+m14NkqcPDSQjJA+9CXG2yhD8CAeYjSX1EVlM8gifY/rHVJ2/pCkWD1tTYTU
nuonvEXmQotNwljYGU1d/y3n4D29tLTAB8EhOnh0wo4HsU++ihyeLrhnvxogGr2yghbXlPBPXdy/
XUDM0dzRc2ZR4nxknPlYyeR9b8T+8V9EvqbrJdiPsQdRWS93qJXloKoobBYe4U37cdetHUiA1Y8B
4SLC7ogqgwDcWWj9FxOXBNY+aXI+9v1w8NRicdRTasJ7d6D8Lzlx7f/EaXc0dZ0TCOyRudBxe/4C
Z+61dMyUbaNu36AOUYmf0lbmvqNnbFFGLOrH8VZ1Qf/lgQYkOwUIDAPNhPppZjak1W2WfichWKFj
qEo7sGV4Cf1d+A7rcqfibtghg+uEPvW09MooYV40E+R0h/jBhJrpjxGI3+wXjXXwGQDzGXzN6Fdh
+8y7mSJLzID8t4hxyMPTOG3HO6rRM5VW1brLZb5wnZB6Oh7eOv2fN8G6WasTWD58gnuMEW1hW0VP
MF4QptPXJXY8uhLoRRfL2jX6sff7OHEyduANAMPn4F4g2aO9IfSnksWblTsrtvNsfYF3PO/xLpGm
BArwFYVUtkuTkp1PHXplU9P8kFifLV2xBZniYR82syRyqz1UcFgbGg3fMjntFHqe1+tQC5lGNmKB
v/hqsLijn9+PGDGQKDYpS6C5OkkrpNq+kUEHJB/SWZW4FWN3EQ5EXbU1zoAIouqP1pfKfkQfRNWx
FKNkontGbBptHSHl+4F1YPgJTxTYCivJfHEcfiCfqAy2CSJQwBpKFXKWyRhUenzpBuhr7qIsJh+I
Jjn43IzsMiKjxFEwqCtG0OxiTIJG+pEtUF53dKfJIMEjbk4QuKrDbY0fV/c6tjiT4ZXr/1jviSQ7
39cXOHR4LEal/2T3U84WcGh8dVvzYPOxQaGY/QWNJJJjxAAaJDXePipg/cUkrTL3GaM8ngqLLIfT
osVZJvZ0BarHXp9eB//s1p44zPJYUi4jlNtqBhto86odThBwa4Xp+9iXSfA+1boXtKnnGjIT8Ecc
ftWIrwU4fF5mZ5kME8m+ZyuA1HxhOjjUENyut0UnlyuER4iPkBoi5qWINktYBoFxpmfIJ8Xb2SEW
oJnsHRlC7Eu7e4LXdt2ucRnSeofiwgLdrItyilDhbvJY1Qm0/qeX8Poxzje9Oj4ES1tB2SBc97Hq
oDlkH+Qa6UDTZAdOKWHUMnAZUTRqHCGtHwHsc1JjiGvCFOch+4BeJLemVAPJJ0oLIwNTuoTHr7IQ
Ku6roLDtL008SNDvSQPPVbmYmdeTQRBLUCS/465CAUH83CnYSC+n4Mz+yTtQ4dVurEGSMVoLBCp5
TeY8mPuBZCgb++z2vuw685uFzwkb5VEsPdWUEYYInqBKd+C1k2vyO9dIMUtpEZdxcVwB5LfDUfJ0
NBheaPly3rbEsUggX39UROxyAF1Ajo9jbD2lhD97rvh0RNddHOfISQm3wxgtIHqLExZSYWykUege
nV3b0XM4PnOj7frB1T9qPGUGL9+RNtm1okh/mkgJwDV3wdrog5l+YM/uBGua1hHymGs/P1nUxRdL
60w8Qgrn6UDSJ/v8PNx8gOfez+jsMIIN6WNP6qUYNFW1sVhvnPIqEKTQkjhw2Y0dNmH6JlDl1cY+
y2Y5BY+40PlXAk6eBh+HuSH5Mg4GrshqtwrmT+s4+fqlEtHhgNxHrjEzAjCbTvOu9sDfKFlYGuct
qRuZvYKgm1Vrwcaa1gQHZqPZkRmVmccLQluxnJt1Z6uWgVTmKxcyy1+6RY9OY+fZGc2ghNKs9qom
1JsDGSTr1IRh4lKJwz2cFRANi2s+QKsulW0YKAledaw6hmfDTgdP0oEXwRAdoxIacATXcawE849u
WvjYm3ycZr6/EfH/ddAksQaE3s60sBTH+9vIpzZgyHY75cLdJECtuTjat0IfbQwMTd2Hj1ZT85Ht
bFR/KmAOE4C4Vootllh4fb+uUaWxtEgmM+7mm2QWqW7XfqOqc9FQoJPLXONUkvcylmUbgVyX2AFc
tFUgAgqgI1UUSWfC1a2Qm9y3fqyIfQ88rol/dK7NHTgG8aBoh+1lXfzb0TyUHvXHuohydSDMm0pk
r0Sa/TaZYO6V/q5Hvln3h0tpMzctMvqAkoekIPXES8VGuu90czaX/VGfK9OYTd0rsh+GxONAXJ9f
G9H+jH/7dnkeXE4OphrcVfrkamuWsWfaPuJN586IMIwDUjkY6D7B9HiqcGQLykTlsegp4Amh/Z+9
LQrRFS7fjsi2Fv8WZiSn0p8utUEy+WfwexuTKUD1Pwl23/6gu48TCpxWcGxrCF5ZOL7se/KAT6LB
txHMgvww1uUApoTjrgaJupuOb+JqHtItay37ht2rAHkFA7nRmRkItbqznVaWBLbV4/iHpydB2c9m
CwGusQef87IoyYaCLbSUmayNpubbyXkbtsFOmSdMiX4/PW80oRwpuSVUIT5VrxE3LwQhPrV4YzTG
MSB3AnfPv9I2W33jTyYwqmsf9G0zqEYRO12RFglHE2G7+xOObmK2VX7iCbx0OYEBIlJRrL+4J+L5
5CGqpwbt2mHkmNsJR0rII/uyWz8cL8tP9Wl03GgnAOFFyBiAk+pVzTJsU95LH1UNnSW2dRwziBBk
SWtUmUME0mUO5M+koDMXpyiKSzZEsc1Asb51aUztl0yr0PGStYLJciullzHoN5xWS3Ww+J8SJoiv
lgqwXxgYbw8C153I48JcQHbSN/S88YxRsc9kZVhWCAYw4J2qSPJ4dHK9lBldoNYfnkTWaCy4cINQ
dXGxjBq1FBBWALQR+RMsu4xPINBmvcEuRVPiUNSwRnNwe9GVOC2Fit6o2rcP/jTUa4d/sKGVYWD2
0TG/zEeMs3MJJhjQyh/RTi8BzTX3mKavgZ23EGu/+8RBncRu39BpGb4OGCDLe872lcR02RTGMIq9
x/gTs/xkzVk8NA6UDS2sHr8ylvGkH6vBSZa2tH8yJWaLpFXsUI8afxXTjZCE9hV5dJ9n+MtY/ckX
+pxD+uImgMYtg8WWXkgV9QKYS7RLQurC42IUvWCTjV8GB/vnCBzP1qYKWiVMbkj2ZbxAvTd8vfi5
A8F65xlkZwl0MOWpGEj2HCV4gwEMk63xDk8NHK3W2NleYOlTJ8ekyLen1b6HutMKi24J3TKwcCXi
Gkj5bgPWfMdAk99+oGyk5BUjUG2i9kX8zCN0enrNbrswRdzOgtLwDRuwDgkNbBYf5T3cLcNVg2jn
yh9uhT088iZmI9LT+RDh2KZ3GSY6tf82y0EPlqDK8npUQVJBeVhFp8u3QQJ7LN3Zmj/7bjYiLIt0
fwkLxzkcDuSxutuENLX9vaPb3Pkmvr8pjxBXuujgSMrzpXJSF/x4+M8o6Ais7utEZe9Xg034IWh+
kHWqTe3QJl2ro44iHDJ95NtF0R2TvdeiwYr59tJoNVJvve99Bha1IlvaY1kW8pELK2DHv0Ni+2kh
NiEVX7dQ1mK5F1Drwpz7MvwiY2doNqm5Xl9zl9+BUeVcmtzDK4zBsgqNaXeOFehcUOjsxmiYbRDw
jqR4zCntnJ7iHsZBMGU0Ee15oUqk226e6THT0qUt2g7RHguXcuHyfBuGHRlyM0BSbrwKqyEftIvJ
Rse6VcJhLPlc/2sdKxWy/+obv/64nUPrccW1c8Doe7637ZtAijv057afzEBJ+kVJ0hOcWU1LffQE
1kJTzE8ablb0Q4q0k24Oew/v7qiTc/lt3hJBSrVzZVRlOOEvmSKN0oQlATppZnRoHc5+itHfIBzs
uRb3IpziuX4Iu9nQNnGaCUodvj2CxDt/CydzZDT9isXNzktmT65ipSgUO3bEEhL+y/OyPjvHWmBN
k4fRyj7/sbd1YeD+bbT+0hSB9NsQh/jsIWg9VoV8DY3SfFryVpUvXohfi6d0ey8FKnU3dTaZeqs2
3Fopca+I2qspU11JfkiTv+YqzeE+RWxDBfPdWVhUzyV/mhWLe5bID4ty7TQmH77EWSEalF3qH6vK
ojnIPzn1/cev+haYsjT/nj77MMaw3ohG9rLAIrvyhUa/xg1oszDCNj/6K1baqyxt7qPbksHnk/lB
TovGLfaxQ8HunNejCuThdy79be3mrHScZggcWTxQBHp1DYVDVsEwbsRBwiM2K8uj5WjOwYdOyNRh
wMKJbM0rprTII/ca7dMpuKUI3E5CVREHqBtR5Py/AvmcSFgPTHCMIUlOqCCnSmVDnmw43tpMJSiS
UlSlR8sYMhAKdMJdkDypwfo+HWoU8BVKLli9fzJceCRqP2hXxvVD4IiwtoUnrzzhkv8HSGlce6NR
ej/6Jxkqnve1W9N+h5RZujBIkcUbzUpxjFCeG6D867y78gaay0muKhB3KgnTWEYhRYfGL6cgnuI1
2L3BwdVObCTIlJunFb+c7Ex79XocQm37jfCsAGrGSKkYZRmHcCX9V5ZVHUsKHWRGHP5lJYb8p6FI
lGqdizoXd1oY/siwFXfk5viMvDYq5cKu12VwS7BUy5D6cRtjq2dO3lhYLEzV5LOo4CGHjOJbyWbE
/jI4FsI6+wHtqlHNCE+oTwmhi/rdkiaQelwgVHXwQ9unpwUjx0BPLkF1Q84nDCCS+GwKZ4w5mR3I
CzRhA1AGZHpK+CREwgjPRtHGwPaJGyiHPU10kyVj2hu/GnDBse6XVjysnMXZEdfAB9w0V3NYK+Sz
IN9dPteE2UhAUFn3qyJ5daBtq5G8LE+3CkIOE3vxf3Aj0QvNJBmDH9//kQJ78GLanrWZGxu1OE43
IPXVaweSLnvvyJYRUJdgJRmxOFTvaWq1gFLYYAB659fzbZniMmOu1aXNhwIWp+QG7Yvsctpo5hGz
jVGSdmzGpmJpGxKTyiDPjgrllYHY33ys+jT1tllnsr9aU5Is6Kxby7rv4/1EqORTfo+d69q44ipw
vtl2JWh4hRaSHhLpL1KUHWnMkW5eN8kEe/CUDY06rHfPj7QuFKuDb2oCv5BKCzk14TDYJNL1wky4
UeHQee4zXkBhnQeTCuJ/jmAWoKh8NhQy1WkIGpyZTUd5EcIL1MTfZZEXlFPlPCVyDLXhpLY7rEVC
XNC1tM1F/QLUMBIUOvoRb8HEKsCS/Wor3fU5tWJHMy53ZLQ8aw6X44wvvVB12NN/mu+5BXReQOrt
+jj2HAVwCNQY4a+Xw/PcTzd22ou5otwvi/0cqOPzm6VVUupCRjgXySdJn0UhCJRP184j1mCuuNUD
XA6OerfUC9HLl2+LQj0vtHKkz3TF3oLSQtmD0W0FtNaeYeHeHIgJlrJEXIGZ/2SbY/ZX8I4k4lKV
bBhWgD1KpHM2VeSe7fyw2vaJhkcB60mKTjPVkvAjPNN8mUqSsY2JTwNahu+KPMa+MQon1SxGHeVp
tRGisb+8NL8tCbqk/UfJSpi86kn15cQ4XozhWfT8c6EhUihMeVEO4AgQc0weAGjs+iInnw4qxTve
lk05RWsghd5yvX2tQKdLH3T88dslICBjgYABj1dP0gXtYkhFRDvZDaCtEqPvyR5oU/9+/LSq6Oib
shm+cvud4xjlG/Jn9/8Cwd6rjJDWpGJZVbkym3Mc6N5vWaWGMyG8dRF2Jt39hTVGXbA/0WkFer94
elbmzCO7+xZz4quNr6m5AWvVI6wbBEwXCwxhYjf1S6G6qaI1wQqshdzMdRPSmtFgSdfIj82JL+Ub
p9b+kSzkySo+eCxgjP2/ICL+yjzKVmhMrSDUPTFMFTOx9CENV49liQ5mRFVY+AsZk+xKooNi81kJ
W3YpUnFS60PhI8XTSnkzFbhqLz+WpZjFCeVmD+fJCxR8iqMIcgjB8V+EycpmsLrYGSBsQeYtHhHO
k6asj8Tlv74Ht/VTjWk0Ew0skxry2YxuxL3+dwaRK4AEDwAPff8ZbbvoKoSk+4ZcC3jjM7sIv0HS
a/+H2dmBy37xhUcgO4C3nYjziyW79hXIL9WOf04gADQ8t31Gjf2w29BDPQivpcty5C97FJDU8aA5
xH/WIeo7mdVqx9a/nW8A1xHeaod6i+R+l3g1IwUX+VFIzxrkN9S25Ts+i+W1rF9HNkXCYFnqSyQ1
MzRqhA+gb6vNUEQWkLvQZwj7NeUdRj7zDy4f8Kqm5VG5xcKe4eCxq/KDsU12Vt3mlBZNcY0ckh5K
QHQ+bdGlV0IcQGSWDzhHkLttMpkrVWfx+1FthSmRnLtycFLgaxzaHkZ20TC336ZPLBSB6UTg41We
0oumrpfZqja8n18TQG7M5Lk0jogVDUvx02fRuqtR9i/+6qSUER4SMxm33O74DQ8cnbEcXyF2HlcZ
9/R61VYcU1LByZEfuvUpKtvOSi37sxm75GA1gtUD60B2d55J+61UUzXjK3510TJ5nwyK3WtLl06i
5xHVfRlbSu1D6PVkQMjSaf7bSwOlTgkCuBdDVXK6P3kHBTqXKeJwkLUjHHa7g3tH0UD9dTVBj4Mt
zUhb0/i1WXIZHVg8QzAl+U8sHIE1X6wdhOQEi0n/SA5yQwnBt1WEoxi5SNB8sAXpwwN4EZWsOmy3
481cCZaJYDYXCiUrAVlQt+JbYETYQBECiG34y/phhdMGihhwh7g/I9lEyKbbdM0JNfGKrbIVn3jj
3gMfQwpeT6Lvt5iqdcJrIeCm9x0Amplfd1ZMnFQDKlfLXl73+OVCu/PxxaWZM6FhEGeGpuSnyozi
fuiYeiyjnHn7VpM3vFuf4H/nsSdiaSFB0cjSqjL74cCAR9uhk8KLK8aTcaqecrfcaO+MK75dZMqn
V1OJ+OtZojFgKOVMfyMmj5L3gQN5HvZ3pY5aR4d5qKKr0+eQ1bNEjlcX/l+LiYS7wJ1QuKI/O1uo
a/68haRbz6yFk7PQp6clblHDkXpocRcE8TB1bAgK62r4cchC2SuOvwebdbXPb9NJRASR+01fjCth
+DRcRWMSScBVOn+onIXIpG+hbgfpVKJ1iYOAjp9kSOsSI0vpliuELXR4kmn4ZyToXJmAZsYAoDPL
gVdCzYXGHbXWhOhXphpiNHMRZo8JNEBosb2ZjmHED0yfzZj6etw2XElyKCkKOQreXjbtFOfg1XB4
9yFV5vjN2S01//dw2GZ6Eisy79rjOqedPgp+VeaqpqO9dsjLsbv46vH88YJ1Q7s+cD2pncBMQKfU
OeNrXUgztGGBXa0QMAwPPrhu8iws7T1lqma5t8g463Uu+ngB/qnOjR2Ll2HKVp+P6H+3W9YCBAqk
fHDTHycjzcS7Ortox5Gksn1kEN/WmMdm7y6+UFjJgBW1/m63FNUFPUshOeQD+G2qLwQ7hZ983kTW
XJWPZjzkYTdq+4Uhr0qPGIiXbhbzeA79hyRSLM6XXSf2cnkwRYZe5bpLtBNWPP2c2TDrj1yIIy+p
vsHykdLV5pCvwBfjV/KVIYUjqzzojJgrc+uyYfBALRmQ/xBW3V/ZnXDaKnitSyss0VfRdkrNUzqM
mllZMZTWlsbuCIE6vuXg8H8xT11CrMIqGDfnxnAgzAwfuGbO2BLqoteGYxmpc6C27A7dx+uecvCH
OdpQUI7DL31ErPpk0vRsVdnAswFzZPqvpXKugjZPN7buRuuq2mxhITqT/3oeYJhYwgd18JHHpbFI
ksBd4VlqYB1D9+xcaDbp+Tlioa0mQRTLI23dwC+P3jZvyjJxWFgwmR/6cWox2+mYPr68TifyVwLE
63VV1v5Kmm6H976tya2TFEHG6rZre8K8kEyBx3UVzUJW1/b0J/wgllzxf59YucYX/Kia8zAvnjag
OSbGdqyn5quTO+q8ENZPLPjY72AlDrnONIykoot5hYyjhAX6C2NhUboaxIZBnPs5e+t6buhghxJr
gHV1ysFROlk7tUjvQYpYMK8ZD5D8OlRI4xFVOAntCT7bfGOzChzRow0JXduJqaDEPMqLHJDLh7wl
+JlzS3tHxMJDKmFbPHYXEZX7ofezyBB8VNNYVHm/QnupvzfoPdueBeZyTD2dx06xwS9t0lSNfXhi
vNeYOPQOxP2c0nHCGsioALZllOw2szUYwFB+9fiu3xC/IXK4OrWxThb1mDjmOVsfCr5X9Jw9L1Oh
Q9yAs3BAzoSk9Fyb7g6I445k5ytOSSxxAU2C3uKTowzb+32l3ljijqmA+umjLI/clI8iEJZh2Cor
MN3JApezO6P8TINdceCVuDfW3CjkPivojX0bLQr4qYsUmPXMkP+Gb7mY7AwWcGn/o/opvdHPnNaR
I+72roDtDdoLUEfltvmhh7EqUADpYTddoVn8ynTp/zJ1gbtDdXgdV31jXPK99Y0qsWA9WCF/Tyfo
QBCPZnmxarKrGurtDclaKAcJY2gJ2oobi8xvglOwi1zb+XOgfxZ49H1UNkivFQ/eOba6WDMoVZUQ
D8EDUZLijyhuajHK2Nj+ag5EP8ixmL54NLKGEDmMBPzmZv95rvxxKGjt5gGzRalasU+MPUWOHv+b
GeJmG9GwZK087TW6ZKctrVub9ns1OSmSlxjjd2+ft3OSa32hYlgIyZ2qUkyq0R87CSj0WCvEnsqQ
bgjDSiB9i62CsahDEIVQO0kCP0i83AuvKjJ0wSR6fUUZ65+3JkLCzaxofKFPLPeQ6OfK/84Z0cab
yFdUjUYSQzguWGAKPs6hX5CdV7RP4GaF7c4rjnkbxvlz0z3hA7SQTH0WQHEwaoR72deEs3iK0Awb
LowyWg4B6PD1J4oRAnrg9UG8YadOogPKaZBrSeiW3awOecBlWesJM0ytmLhFdxZakQNbRFJ6mstp
3ppomSvgeRA5TrBdvSHH3RXltJW0W8kI53OJdeZroGCk3dfARvBpuxgmdQDNZRqAnQygiUnBN5Kv
iiBob4LazFLrsukPLFXpBmHQEcuYWAJAQWWKUF/sDtgRUaejYvP8iy6FRxxjXe2WH/Nwn65VkQki
m0ixcnX0ny4yjn3GVV0EEI/pcsdGLp7zxKAC2yKYB0pG1fFYDTT0nnppExjYFZ9C6MNjGSLLc7EL
GFAtrXg1XvG5yMfz6mUxp4JMt1crcG9wE+EB0HBHkSPSUu7Ski18CzJCFEIqgdfwtqn4vvWwZUEL
Zft3smehMHt24W25ZCbhmy3GNvXysU6cswCzQzalU69vnOBo/P+umxog6wb5vG2aATTjakMGi+x7
lCs2VjOhAEQeKYb3OAKbV0DM5xGdzp3FrIxpsrmFcsqXeF3Hu0SZ4Lb4OrqEIlX+dQQsLzVI678+
Ysr0FzpEy0ndcNL4nk6o2IOdrwqTaXqJJX07FUgnGDoYiUhCbsht7M+ZDVyjPtelZllv/PZrFc5y
K0dJkwj4KruPsWwTiBH+t5ra24J7T3nMwMxfUzb5ZYtsUhMhdqHCvLKT12cph1+pQa55PjBopJcl
4jidR6/GYMwUeOHvif0NNJMgNjvNfxGKO4ocMEfoj2qqoxCfzFPJEnr2bf5rE9X5dGSxsQjXKblU
P1/9CuB6Abzl7Qy5VfnDgD4x5raZuQUNfraAijqr6srTgu1izdmesyYAzqeyT8o4IVvak2RMXDR9
KlPYzqitzWHnMVDe1j3WUIvUXDH/Ueel4nXymHyN8oXuJZnnT7fYur0fa+H/k8NnTmZhHheSQtBT
CkbKw+rjo39hUG0vHE8LPaltYtsYTU2GDXoZyQPpkRllJm+U3mLi55Q0nQH1MpH7flz6phPnFze0
GMCrELiEzO7A3mM37B3S4QwyRtTjJ+c7xO5R14wwKY8ICniCyR7u/aGQaq8GNVi4BdxDgsLLahnB
CCh+JKSBxPuPrDBTFIgUxagagSFcLe5QWphswT0vzFIxEMfuEX7Yp0KsKlXjsPwb+v3U95qcRhES
ke+bCxQ0UbFb5nFQJ57FBs7vKDhhB4v0tOZBQNYLnE622WKskzFLjl0tgezN5TH+VU3Zi70Wod9r
G3kauH+gJEid9vr0Zk5Ew+96DpU1jBy1JDWGsRx2VNTbLbYHR4JLY8DXHRLCK7n3TbeV81T0w67f
qfbPGgl6l0hqZsv74/zHxIDwx02CoadlBV8EfH6O5RyENjwoF/QEikY+RuIk1LHpdBH0b4Y0hBQF
ZrbmD6ytVrANUvckNWbDtloWdIBq92Xg7CrMrvps3FN9QgWQCuOFY9eHPLCJSvRw1nZ/gHjgiZP/
baYxx2fwuy+fU/JFDxb9P7ltHCaNgtDHeaoIj/p3u8GbLlMoyDP8shekYQPF6nis3lGl1+m0xSeQ
bR0tRaciAnpaV02gps9Y0UFrm40u15XDHtm3OUsU78w5Cu7UkYrqNE7fheFSUMWceLugsrU/kFg2
0AwbkM4VGSEThaH7GZiQV9tmbYP+xXeaButQfN8EWDBYx18VH5MfCDN0ACxPnFRSfbIFRu/fW719
0NSNX4PymnZ6iY2vfAN968qY+qaGua1yxfcj4PTF+3XAqP9Q6Dfr08mddcyghzBctIU/NNL3Nxwu
Lt2x70pxnS6d5i1IRK7iY4/2XQijxYMTTJvxXqV4htv21k4NTrMK/Oh4sRu6/zkziTXBHYeIXEGf
j6KQcZydFj4I0OWYbi8KXGli1ASN96xCjqtreIX5ZAUOI7z03BVEf/ZmGXS8LUX3evd1s3V0b5+g
q7xHGWW+VVU3EeBxZ/2Ov++lFB2a0cX1Ht4pHP/EOv0RX53lWFeOZgFSdeiRVBKzRLa04HoJnC2d
64d4JzpHP8nqlBfH6+0RXO44e8D6ofqW+5e6B8wpivmMmQBFMtoS9fzlrmmNSorKT4Bo6R9uLnMT
lCmUlojC4U7WFiAHnRMXqpq2WPrehMnxkm0mZQjyjUtLlj4Aess+joNUKwTKDL665wIUrK0B4ESW
18VehB3gC2ByiaQPqLyn/owmsN3Fao23NDaN96CmQqDiYEkCb8WmVIZeZ9BSaRbHuhloaMLcTzdE
3OiS/K0CTB7e/iKAsFxrcYDGSkSa/X/JfVF6/h90hcn40vxtHTNd7QQfkvC3c1n0Sq3POFKnBkjJ
2rL/UG18VqVvlebLvOjvCKvkZCyMAEr/DClC3WIfgUmwcpP+K5PBrw5Nmy6N8ewK5pkyc5dNI0/t
h0NY3b+6RXQnpq5bwGpI5RHvzCDvKnKABlnLM9YxEbL0tUnc2YW4t9ml6yzvsd6DcSnqY0HJOwT8
JRtvW4YEbB5d0fn+6oXb+u3FSPdkCACfqKQQxzsBHmeDxxy0MZDcKm3GmnAbklR8gcuY7uTkXFuU
zwGsbI8hVIZpESgiS9kP3N2CjfFpanzSw/6dqrLW7xTZGNGMt71LzAJjV8mxIJtqZ01VQxMIXUQI
RDGuUO2RfP0lTew/giC+EipjxEn5BovCT4AzBNsiep+PNiVYjPZUM72fQEzA1MHzs9tv7jW3pRSj
q3+ifN8CMeKDhSynA5rkEDLLlxDglCKR5eoVKD2XaTVMIZK18XzfGr0OzeWoOGNqfVUkPC2ltyIH
VRNVjlZihDJYvHPJ0UV15fsbegrvp+M+a3b8MuidLCNy/ORbCiLmpqZmYLrWCAoCM8KkdMifNa7a
Ef5i4d0LWKqASwZQD/5tlHTpbgKBUTPN7qxOTs0P1jYb1P6jmC6hMLYcwuo0CUpKKa9mGRNB2uW/
5kjV8smeteIhXXu8GDpFA6MeiZPw+PIHvxaOU4secCiYVJ/sINo7vJpabfbklSKd+u6bV3wu83EX
jySs7GcQM0VbONS31nVp9JLwepg4bdSXwjVOJLeo8c2cyJdZ1AEgHBOWvNrDYINnQ/0TPjaOHj+s
TepKYOAprSoU1ZHT/g51hAYKMaNlp2q/rR1LNd7hzOhb0yNNEbBoxmRhOnWUZSL4k3fOtsaONBDI
TdTiqDOpAmPnYsMAhi6JRnTJpFXUXR/rSDDSfYACkt4eUYA0d+duh3K2E1L64AvzebDjrLetuMJj
zKmDWyPTE/Ukjk3IHIN9tA53akL2cWu8Am6tnsok2UBFC3NJHXJzRSOGQwuIdJD1vA0ZtW8EpR0Q
xm0L3s/pa0PsF5fShaqEhxfJUhSunRjIl85Ds6wGZvpAaqIuGyxcMgaDxoAd7gG+OsEQtgweuOpI
fpp+LQR7JkHCNSlyj+wac4P2bHymyeiKj/2L+0bJvIziPZ/AZLKOzHD+fiQrr4cyGxfRy2ikgelG
aZCt9kqe+depOUhlpRKm+OuByE+frssg7WCDmsNsvDLeiQF9+tBYJCeRRyxeI47FGiw6PbkIjMiM
+zCbii75L7HP6hJ2tzphKks4zNHjmI7sioOeNOqn/Lwah1LCgFbyfMYCSHYYI3uwEYsme9eFe3St
qCZGFoXExRz1VV/LVXJ83IhYvlWTiN8z4UHclvN0eJbCZ1iCOml6y93HoGnggeYmY+2Z1Ye7rqsJ
OdmIho+Q/lk1KELI1dkmngl0+O6z8BcObQ9LZIXb4g85ydIJW3dDXqkINhGmbzb4tIcPB34Qn20K
CUg+haS45QEq3qGMTX6bPNxhfgD4JdNTJOSBWERn/ynUxbzl7LEK1vlVCpWOTtEDQ88fkn4lKz8x
z2CIWX6iSf5CbeRTvcDsWobisqcxc1+Ipis4TEkM2HXublYIb9Mn/ciKzQAI0BDab50xCaHDiFl8
aGxMXdBlvEZea0Zbj3oqk4e4OQmjld7B5BlygKw9m3wPgvVDmQ+KQ1IKtgZdsvVTOw45/wBeMnY+
Ey6bbtPzHpl76SS7hq2w/eP00cIpeyJL6y8LyRLTS76Q14T2jYfjWyGhfVK7xws9v4Msvk8LFNgw
wfXv9kPstFshq8MoqTvKPRBpd66PCZsfDVtjzKoNbqj7xhM0rv1504BpruW5i3HOwF0zF0AkZ7vC
eFKYvveAbp+6fPdL0YHY8Ia8BuUQqWeI3hY+9LbnMH+gf1c/qyWq8IGVBpqD7WvQurm2ZNOqSk3l
Xuq8uepKdMwWSsPB19PPBchL8yEEm3RozIxGxQJJuge6gLFlv/gP7tBrDeChWdNPJwfRV6gQkdOg
fNBJWrbFdua+IM6DytlgdtMv1Xh+kVuHICORQZLZeYV/rBn+er7BC6IudnNZklIAmS+7zVCsV1W8
eAJvNjre9esiDQD/gVcTKUFUjDVUtRwMEWN4GFMtkgBFkxnc+/jMmXtuj6CJGA8T3w4v0RmrXxv0
fk7bKlubyqo8rJj70v8465ExK9dJ/rPRVbHPhVMzFTWQYcYTSMkiDaD8ZyHVibO+zOnby4l8vbw9
vwowdiHfqxqYjW3juTe3NVwPPDSSCYIrrDVxP0thw2Ng+A2ZByDCZWL53mlhq3QTXHdTbSM/ZIr5
a6lLwvtCPtckpD1Z7iQcGRUjQRvw/ujzDOmVf29/6a18KbSKTVuYdn43Bifv+2zsHtZm8k2SCIhl
TGqEkPz772APH8Uhu2xG18lRZb/rPGt1qzRaR3/8IXtH3Ci0ukn5bj6y2PneMR81EYjXuaAFYxFC
nMV5/YN9MXHmwsJPWj1wd4aeWjMswPsS9S/buFOH3HHlHkuBxb5rf0zUz4W1qEoWkkX/CaCb720N
8qhIVTXbqA1cXuGr8TV4vXhTVE5h9K8ZH426oyo/AaztHoSqi5uis1TWfx/iYbt3sv4RClyqiW6N
EZu7zT3I9YmZeKbePv1iQaOYhsGLWxaiJpXOe0bmXtYk69ES9ELmrXIVQJuIq6V0BYJxVSUQFAXC
wWW6/GlRQAQWcVQlrg2Gjt9JCoqy4Dt+79igcmt/8vJWGzwjPWStfGONCrNhRt0VHoSqrji2QXQc
zU7yj1YdiRqc6K2MGuz9KFSpfqhXT1qMM3Oqz3r/rmGvyA0W5FG1eCwDfXOJTjt/B08eXNtv1iV0
eru4Jh/VcEKkK7XRSFDFNSOcvvlWeFFj6pXUfwY+wgJAwTbHkdEF8gVU4tf2l6XOrFTfJ82oMt62
Nzh64lIjabiEUDLK1PromFNLJK4eKBPgt0XUs8qKdQHQDXSI3xzu82CObn4twhZti906HYHXRi4s
mLJTUMA/bFoffBipaFBxKCtB24z+soGOvV3BdAUH8kK9giZJrpuIIsi0Pvjm1v63PblaZLPJYsQR
ie01wbPc5Iu3U0aMQI2H9o0jyMqVuIlY/L0yDgBNZA+iYIJDit0HiMCkcd/ObQu9jSIceZQNsGPG
wQGVRv0FADJDEa2iybY9KlAxr6UaeKlX6KGCQDQAyV+puOzYigVsvL6Bs/PT+ikd6DHQVcXMK/zs
UsX2oi2KM5aTFu7pFnvSMRQFnzvkMMWoG5ZthQAbfwfWcxW3/Y5ndRYMxLJPL30ypIo/PKbfKR7V
xsYpnsuiowbGoBovN2tqHFCPXFF/R4b9m/+DtB9ctYqXTjCW832HF/5t46H/O5hw8/v80+obRmJV
vWJAjtV0oLR8VCERxLyb/O9O8kJ8nwvikkkjoKGNKj4u1yOiPiUmt5aVSfAQi7yHBjMjJNqU+yUH
iSJxPQK9gPufOFUtLqWuCCawlgyU3yKz37FzIZiUxdgfIfT2KsMJ9dAzfP0vDtCMdr0UWUb6ZaU7
DQK10mRcCaESzhwyiw5rZjm0IyWOZ/FAho3da2VhIIvXIa8LNBiWBt4aaBdr5Xy9KbmwA0k9GIzF
xU3bvlmak3GFzPvYSA8CSLgmuaRrKBHoWO9CirC64OUkNmK0bl2uCMhdVJH7Ci96Ahuo9O2agcPJ
P8faWHR3iFcFY4yaXygl8Kx5KxGKr4VKPOrN8FJpIixfPgle7hkBx5qQUpgU83QLrT5f82K8PpsB
kLElu+RnzqFKgf6ra+F3GjizWmGszzcfL83MHCwpkTrcugySzrgnda3ETF/7j5OqgOx86mRfoPSe
3fQ60xZdeIRwClg09fCjptMu2Vsz3Sklgz6NyB6of/wnrNnItz9mYWXpJYCCMBb6NSUxlCFlI2XD
RLrISOWSPBsRjZ4baZXtnCT612z64On/71v7uszYpHEvtG0ekevifVL5TCT/32dA1/8lT3yZ8Vxl
t2LNJ7+9ZCr1GMl6mpytL+VPIA1f6adtNI5MH3jfObGJOtHgyX6NTId3+6PQsvt7T20vL5pnAwjV
tVNC8skpmwh/qdw7QbN7y4mEYuklfwr1gMJKEng5nu12yRoqS88nsDw3pp9JPphX8ww556rZArdd
9NDpZAbRLOZ51WdtrkLfIHgDA6WdAa+RnmCCj83BFLbKcpIvDcuJ8w+KD4B+lPWTWd4nrL6lZVYG
99TSW8CWSDknR5h6xQcomvMMsVGyKnHlJByiNFXuXGwxxXYRLCfAH7pDiTdKuw1McIc04KSYrGM5
kpfFWdu0D0Uish/yzBBPgoYtsZgg7pz+sbACzwtGxel6vc4XOJFG/ecKIpbCLqqAtHUekH6t+1GS
VvrGRr200pPJzHEhjFQFmeLdNtJnjoha7BMO3QxjINu/wwvcYU9/sellA/q4db1F9AlQj0uHw70E
FJpHT47LeQ3X8+teE6JVxVYc1/gtg5JbQz15GW26kpcxk20eYL5Ikh5yjC72wUyVyAZjc3u+6RgZ
ukI3MVWUM6mN8TbvTn0zXD8l1q02jS4CNZN1Q2xzkVHJKswblzFIcL5GzgZd92s5k2p5LF8a3mGg
vABYI75Cr9oexzDRA4PuQ3CeGn3wdWdo5ThzMFwiZX6BUSTzBBY0QV10PDACj+S/LvR0mSiBxvJM
HxkoJ8qwSgVhjZr+V2QvOyP1A/kdjOpD3AUUMoW3sHjaCryrph9yosY/CCFr1NYkTvdM/lWfom3i
SYqv/RjcSGaK/woMUOpeGtmIZLI6eDRpsnhMmOmLapUMkyHse0+lwzyddOi4rHzpxW1q24g6wT1a
xtf2gNMoPJ9UtMVnGkCedsEkFMyxf3hMx/mJjmpceFRvioaQTv2NqY4jpbZewHmbMHyinBP8xJej
IYlOu+ftCTpkebvotSUK8LJOflyPFq1fXMKZknMarNivNn2m4b0KOlFHvisrLr/BAreXpe3g0H46
1UQl9a1CtgqyCsJL+tT0wHiWh9+oQ0OYFlkNxMvrX2wvyZs+cMHEiZ2QL984OKuGXoqBxWlgNp3c
ySO5uVno+abVgIB7Gr3jgIwNMhTm8Cr/GK+E/brG+44fqsf7DsrE6Hkk06/qkhpzNDGnKaO4m6y8
k/lMnyGCWcJOWQQWg5SM+rCiu83fJYGzo3vNoVqDyhmsfxRCIDJigu45HHbrKTYSEHaaec2pukQQ
Xm6UG0BfN80vCyh9ZHNqYEd7fLeYjDv65/kYrW4/QCc9+Pg9l9VD2ibSAT7BZjJkFCN+a00CCgP4
D/i3SnCL1+APPoKDrKphoecviemsgZy0e5aj0l3nNljPmmWyhhzOIVlarFxaaLU5wN5LXvYZtdbx
aM8F0kRidulN2i+rmZD26glSWXav8k+vg1DXDmKgkxpru8PKKSPUu/sPM7gCO7KFyp2Cw4H2q4Xc
IwaY66/4uxH9Gph/w7NzzsuVS8P+MTHQAXuyoMQ/+yH0GkrWtuM/oqtT0EyS+dWg+3uDwroyfrSz
pJixhYWzcsWlmgQNNNrZqrZsAj9i0zREZS1p+T9AkyI2enywMlTWyR6E2VDVpTjKqAaZW1laJ9wJ
P4EKx6UOxTFiYTTwo4Sz8zI52nrLot5pG+cqLTDfc1g6ugi4j48EeSYUDPBipRUpyLlpl9MCI3rl
f1tQlKybPzejkt86s9sBXODiGIcY1DZTia4upE+OJeVcjBCnM6aIQ4tMrcLYcIQfVFwhjjZx1fQF
Yb5KCmrtygidWRJNP9bM/9ixdz3EROOVpYbb/K9GHmbG5CfgUmznCLPzYOCxFo1O4bEv+JSxkdrX
v5RvUplGHqakgUf47NrftbuLTm6FFt6kupT9Wh4jVuwrX3F1mJin4bTn6yUSqfZHTd4Pw+wSmy2i
ItaPuAGIorerskKGZmYdJJcTRzJXPfaXcTCk1RGlGRtlXqRIfto2kkpeR1nsBNrqwxCanZ3o8MgJ
zoJeKDci25/MpJ/W+mjkUsBPnn7ux0LkJQYpsvi4IqnGIVW5Kfkcfs6aZVHG7WVp33JvinGqdrfH
Q+RcndBeU82meAqwNyIpnDxZpTg5GMEm5+bifpcSmBVuLSFYicx4xAZD0qVZuwE24CJDi1IdBHDc
4qyHkayrpL0t8GTeomeHguCDwlzSgn9nItkhcYcr1P/X04Okj576eufwS/HJ0zLE0wsi/zhXy9gI
i2gbfLDfZP3khYb/SDvrnXbb5xqU+Q8gggKBV6LRAJi1ELTI+L819rB3XsLJLYw96t2rW4STxs0Z
Bek+Y1FBQR7r6sob4pv0z80bU+eqtE6mu2H6S9SJj8aA1gOx7a+Tiu6D4CwCNxLJgeMGnU+gv/BC
qjxlclbJ6fZ1HcSTQLPrYKt7h9m+VZ1ktqWoGZ6jH0Q3w5ukVplE3bwsjG8/wlxoDOUJNGfYlYSK
690TGUeS6S9yQeGzVxOXWXoJ1brhCuaXeBnwApPCNpQ/GNfTD0983GMFfn15TwtdezbJEuQXZnNT
uyKbMGou2RWHpKArZsKuMy2mMUID/e7dEqq/iamZW06R5iS4vE3DrdWLhIva8aBMKOk3rSS21O80
4DA7CK/EnDSDFVLgQ2CyOtA90+Z7nf0VWZiNRti21HFiqgPW/LKHBWoiSa4PJGazSGeZos90p58g
dWmR7yPwlRTn4z/mDmi+b3Emg8HNY8HZPX2r7X4YI/q6TueL9xJe5iJmwP7ZXvMuYHKJopycjVcw
eOFleHMX+cIEKW5lwVyjvL6KnByoleFjDPwL7ADi93jLUwquFEIJFIpMhsi+b0jjAe4so9EFUlfn
1zGO2Ed6A8XdntCB3DtttKQkCpPRbtbdaKtS9ela200/EYOk3lKPidiOIEiWFyPna1W0gQsFvCrP
ZjPpPB5RxI1VeFel7vOG+C4FTDycsquBgmv7DH+uFSmgH7LTjdMyB0iVkcrAKHF+/vPRK8y3i9AZ
Cpzo/HJqmyek0ipBkBRdKG5XEk7tWgK9fJ9w4pnToXA4WA8VwM7dLShNkkjZJt9MDjSvT2frx/ap
F05tc/Nm/eBoncsRh85usxePwdWmdykEvsUv1PQesMy41wV3gAlC8UbxIRKYb4bP1i8SoQzC9pr0
AzwzTg4s44NcvS3C7UeaZRG8s1ACl9MMXWRzBGC8OAapK0ZC3DWk2rP+t8S4wBa3UeF3gNHA56Vj
ckucxnFr3WNtRNIbLe+1LkYoDKRp+P6FmcKKWKb5WR/fK7Zd3B0dOv3UXByebLCpRywDk1ohPMzo
qa6uvOKGHBKuVBmK6ROoQIZkJMp6vp6oq3bILJ1/R/J9aO5wFntDfiPWrplq40v9R8izF1d0zst3
m1XXdBWO19lPbZlA+phZvi6mZHhLBy4pG9CSdnzmlgeLU/Rlmwz50PILRQEenP+2Et3ephBY53Sx
+nEyg2f62x7piVkbhacirKSRC64du3LOXxjmywx5QjD8N2eSu10Uqr978+L+4oKGhUzrW6JZsXwQ
9ADl707bq6cgl10hVV8g3UGvsy51aVfEpP6omNZEPQXzER0UCVcagUudeMY/TBKwjjiDc4DYdPeM
VyC6teCBGiHBKb1+m4YR3E/cI4LlHprKifM76WRn4nQWnv/pkoeFW6eAuKLr8YwgJ2dVUvfwks7E
Kp2tZ9J/qUCrF9/wIC0flh4XTq6zuAm2zeUeFVEPP6U+3ik7ts9CnBKMYCtXwjRdaMtBXhL4IPav
FyM1N9NBdj0n2FBroD9PV7Xlw8q9nEpBfNYeMc+VLSiwNY+ROqE+I+YSNY8mo13N6sEwkUIcWoP/
UkuthUk6YbbgEia6kl+lENhot6c6Md5EqXoERgvAwESTaWOyHBSBQKv3wDcd47Hjr3AKKF6Pg0vF
yhE+eMfjHawpXYpg5MzgFUiU0gjDt0Oum5fm+OfTA1HR/Cuyb96B67j2OeJ4a1GMlyau32GfKErG
stbvCaliUfW8pqo16CKX33ge+PWLhRN9fy/ykz2WphXlDAmxTQTIE7GKJFXINhwaZ8ryGvmhgv/Z
AZN2737Kq07teN9+PX9OlSeRjpveRe7DELtmoJdChBy55q7XxN4NMrFKfBmJbsqjzwcMuRCYFeCe
8UfxOglNvfIVpsdcSs8oyNUwjWdOspMqUk3snVtWjO3JrGjksp+MrPAu9yE4eWKP39EIRB0IB7ke
/ifcFvvO2CeJK/emCqEgwDhTuWfQ2l3xklb475VTEOHSH6bVK0sO9Ni2iIjGaWTsusRALrBfVl34
4uPGIVbCVHcX3ntxz3oTCop5HNryWiq2RokqbPfgaa5O4o5uwI6ehzQGp+M1QhOVJxAf/aGBajcz
+xh3CNc6iVPsB6ETchDFhjF3KMnpeSFLTMay0QN3A4WN2P5JP/JKdITjG8MfXF1+d+gx/y1N5YwB
FZo1yaunGtLFRB+ubIV0SdW4ALrJf8WqcnpG/+5KWT1HaTgM5dmuYjxLHHNz6U1AHEiC79Y0/s8E
5PSHDV+YmCR7RulbXNlUWRoYjdMxKRRGu0Ypy2QSSPVa++Hnv9J43r3wW5XVr0Lb9zV6o2+lR025
sRelkPKbtLuuvbN+1G9an1NCE+s34tUf7TuJowMN2Ib3kgoc0LAwYHXGiZZoXsw+GpEbIT5uNHjS
rsIynfCrXsapbzZRNA3yGGFfzWqHHN3z4P6ueCQlzUpcW31wEKXHNQAqOPGUZiaYQPjT7n0Lmrwx
361Gd2Er4dyJKzhFmPyPael7cBpWZxtUz73Hsi1i/1H35LHuA8SmI4QniV55M4lbOYOLlB28UiEu
SDY3zw3sBl0dtaS+IX1WdNhF6lkBu7dAj3WJi8FAqTolbYAcuZwaiYz3vcQLJbU+7rtquTViwG1k
Q47e0oG+aVNV8/aHb7Vzzswv0BvfnSj/KMcwM5HGbotYJrZR3xYgaIaNqdbK8rsof87oPUd5b9QG
mmpcvE962w26sOCb5xP1wUsO1mtNiy8Fz+7WhNrhtkWHWonNqgcJfttRVizYcCJj7HAfqr3XPnDg
U2F0znK/hnhBfPBx/0fFaSdjbxHkLZeF0AFKp0VMlBltyz9z2dO2cSJI168YKvA0e8f8KgZs6/li
QrO7y3nW8WEZkkFny/tlWb3cvpCj5BSMMQpjbcOqp8hD7EHqjICjYlt55xyku2TylBsODYyhf5DS
Gh76/c0XCjnq7fsUM1xYnAJxUyaNBKxZRleAjJdUrylAcMNkEFVYTJ1fKc+7KpnkQASpn94gt+6M
CW82cdGcWRcZDU+P4q0oCIXiTRwMEvKRI4kDcjGqw5L1EC7HbeXuJ87JaauhVa6m8cc42ugHVg+I
lNYfUkfUgojVDonSdSTjOrtBSH4XRY5HctMbFa+CH/sz9o3LuRhEBfIQDp4ctbwXY0az/7AaLWiv
mk7Lygbejsg3+0/o07pAW8UTyCH99A0kP5MKXzv4PaHR7O+d3KD0duWiMuptOo12p5aT9Es0DGMj
vMIa0hCRtTNoxOMDJsTrSDcZyxSIvbINUUwiqE2q9yP+d/AheoZXsntFse8M16L+Q9YaZP2+MwyI
QomG5EgyYnUnfZ7AI4aXXKbCl6yyrFh/P7vyzhHSwPQ23+qyDKHSTGr8Av3tXgdSZrovyngTADbr
wgorNcaX/K6iLLdhUJUxH9cjkBj26WH54ygAb+NKI1VFkYOOSV3B1ATCWT6zgY1wyJkjogBXx1jo
TUd6aECo9Dus3cDtnoPmuJLTiiUoCqvCb+Y+5p8eWCwy1kxY9RGULGnpZZ1WN4+TRBH9oRXqgw79
+OnCxWWT19F1siNc5VP1Ak1I59OtKqt2Au3yLcKRgNtvIKjcjl24rm6kNyth8v6j1G1yYG+60aym
X8Wi2xXfkiHakxBqN7+dE1hOEL2R6KPT5ummc58aIkAQWY6diE4EO0MNaz2DUzVqLEU0IFWngwKD
dWYYFVlgkmQkGSQDbIY5tpoTQ3qvFHlprNFf6mcaDZm70R9G6IXURUTwkTg9ClZP/Jmq34gotg9c
JW9VAlWAhdhPpe+Cir7oZVLhwbtg4qiPI+kJxHW7Zp/bLvQL0mc6tDUw+wJCmJXeXCccTrTRkCil
DrBKK9ssiODPGVWJ3oUhuMwV5jZk1/qUL8hVMw4HXqyB86NPS5jWQp97/9deioXaEPXRLK+Ic2ER
EIww27nvY50aQlXkzacqfvRAViBHlZ/44sL2CyYUnypdE5aeEGJsEfJHUJHKqpKrZmU9XDOmdlNH
EDjS6KpFN4jXQFIVYSB1XxwikUZOL2hcA0ncUp+/DC4iT40oDIZXPm8ESLVslo2JJmBgd0skiXp3
PAacZJKxtRtp7CuhBJq3iZ+Ok4t1kXCN8mS8z1z1qFTd1Ye/WhXGipIpWErnKLojcd+vH1nDORcj
DlV0wH+t+LrS/y88/lUpHy+F/Fk5lxSvJaT9EZTC4Cd9r92xEvdsDQhbTvrMIbwVVn+MSFVEM2Ea
1WVFJh0sxOGkKLK2XfNwU4MyyFBmHin3lqj9UZ+ogMj6nwgIb261q/cB8MIwWEw2/6x6EZ/NsGjJ
xY13tAjYkOmZXv6SyPo/2ZSGEs3KP/1ICqN7R8qOuyJA9Tc6WxI7984/pM1LWD7VKkh4P5Rcm5mQ
v4QsTvI2QCBJBpECw07oUgkLO2iAz1HAL+ea1W5UWCAwPD3PGugsKezEoCKXQooXDHeagkYWBpfT
NsMIoJZh9zIoVvrA8cSpsTsTCx8nHxjywgnNrcuLJDz5qlE6zQ1H70Yt76dgcobSAu8yV4noiHYJ
37KF49CwaIB9kZWml/PokuMWFTSvY9bjUSJebwjCgOq9xF5fgdCAMrrHoq+wbVwybtgh7zlXmNkm
sTTsLopzua0onev7trT1c/CRkrFLF33wWKArfdW049JYnSrwMNupu7Bf3yBomXoc3HLl7ZG0HxGw
DKs5xdmroaWLDAKun41oljqBZxTMJBsK6vhFUNeZ/EqgzKlqbbrUDOEZMkqisiC9ZgAeAmYqzXPD
LJifPPd84vjqgRZb9FEEKingfKa9M2QwtMMorRjRwWqJrQgfYaUwHj+eKmjmA3F+TNScIZe0K9zn
YjVhiq0k3cT+CnEvGT86LSWlodEYEAdgjy07Gl8zJYZMBgsU36OYMoKTH1UpZNFApnyK7l7qMu2r
F3hIMvq1BUg44UT39Alcvh8pTYnOVKgFs4MjWqIwnIWjrTyD9MkqkqtJoFD6pBeNbK6kfsqkX4QS
hBrTJm6CPKjfQ+UFbx8aLYD6gJm6MWC5UoXLegarxkLbdCCTY4ku48fA4DwUwoZs56BwtYuAc7HY
ndkb+l5wF6KNE2SBSc97hQL0SJatS/YhuBe758X60tNM9DJeB45pb3z0NUl5Bqv5lpPpjRLHIdbm
yn6HXaK0ULK2Mrpj+RVcb1fxnbmUsMHNyI2pxN1X9vNpgWX9HiQbCYoWPHl95FIcGwZrkuWVNM5U
8BHSySLNYyfX7IYLMDkSTK0ktZUH3LLxflbS3aFYHPrp1yCukSaem+Wn4N1m2Xfn4BpV7/W8FNnQ
I0vEsiFe4PaX9yNWYFCTpJca3GywV3c0k/ijtbQExVQp/txB4tYSq9dB/zmieJ/1yTi4n2q+e6nM
nC7w2t6EGMbM7cr1GGUc+hCB92uuHMmUAEEVrWmfKbgqUlQYAUDJzc1V3iL3tMhsJwesY7RuOTfU
VbyZn/W6Po4Tiefyei2vTjxdFiQHc6Xijv1fUi8UsCtYpk60CwClB7y77AwzVMLKa2CKkkWrdXOy
GO891iLoTmG73Q/tzFIC1iiUA7fGdoum8G8kbhar9WUFZn1yejZ40mNCgiYz55DbyD1RQTRU7P/7
VMrB7p7GkOVWUAmk0zuS2u9zqiUp/TsBqALl6dsqiY7s2/W9E5AjM8ILVKXYwHBehh6gZU96mNbm
j7n96Au71oPsl9br6sFBBWLdbs9b17es7UFjxnMbMNqcrWYcfXGMCheSFpi1IlUSMBy2ud2BAROJ
oK9GFp1sJ0X3RMJHfGj95qDwOxaUTVfsjOwRbRoydqW/AXQJa7Z9/GkSOs4Vf1ixgCEuITg6vpk0
CYmuzk1/FQ7zWNXtU39LtX9niZdt7T5M2y/q9agqxIhuBrbNAcmBtb0z9DXVeBO0QvfJbxtM7A0e
/uhEU8mnSWKJSOZkDFdAHOvYASdeR5DE7YTyc74R3S7zxEHld8YqXIBWuj8DCz/IzRksRngqoxWU
5wQKLZCLV5Wrsivw8SkTlEXO2VaS5Tsb6EQYOJyXKnwANTkWqS6gEfu/2UUelw8oEGurwTSkEHZ2
6l95GIcGfKaHZ2hqA3W5vlGUucun1PgRVPrkhcCWxgCXBI3EdNPjy4FzOCOeg4w/DzYpW/chfmoK
DY9KsmVjOuGm+jqUB0VNx4whZZKcSiB+UvlTxPbPXr3l6G2k2jJaeMzGzDw1S8m1eIUbbz8ar72q
HDTI5h8hUgv4anLxYSbgHbN+kw5V56NuZEL4QwI5QwesgGGthJONigiR7wUtE1gbtICIBns5Y1sk
viwYo1Ct/wmkkgvpKpo7wPbuOraRY9tzZoCF3pV2hxNoH9TJqXSiDhAf6duAm43T5cY5hIUpcACU
nxWOV6p4a0CYyxfQbJeyYUtBTpdjSluyszN4UINgGOYxtogHr+3wq8td5C1T7oPiV10aXowwKALm
Zy61+VGYBGYMG8ZPLju9wqFDA1Hsz6OJVwWyLILnmF87ioJLMhPwaymb403QzwXFFQkFKq4KhqF9
k2WFzZxxNaRibxP3UHvNj5TBLW5yE5bN/VuIbYur7mebvAWmRC1eYp85r1KZp9mSo0E4DU/P+30M
NXe4EAOsgp+8B3cNoxT9y6JXAB597V6c+lkSJqasmjPfIyqBgSv8lg6zB8AetB6IeHig82Hd6mWH
IV30x/DbX1VTBp4PUlLiJIQBdc8bXj3NLVuvst7wfuYlKlesaoPm8hPGn4VOs8rCvohOFzLC+DEm
WmeGxqRvRjBpx5fvW86rRskhgB4f+phB3ZQMgAlshT+3wnsVMnQbyt+6F3BKZWzIajISTitlXr3r
ACvXHW/xum5sWUO+muLxAMqbuPnDTxah3b1ow+weBB0ZgnJHR2QGpkUEuDlx/vRx2MYFwzLnKAG8
ln9BmYPPN+VIYIxXwIKpu8n+jnmIYC2nESeEMwySsefo6FkTXvNcrVeQsO1Uxa3UnmWBRuodG9yj
h+tnHqzHM2xRGjknnCF8sIxoqxfgxLPmFGLHiX2c1wqK/ulrQ1uDJNJricE8eEw2+TF8hy0dm+RE
eB56Yy+F8Aj90OsR0+pK3XDV9xiViJygkbcDAteq2FVtI8ead0zqdJJHSFfQ80hurCdaZxNB53MB
e6uw6KNi+AWUe+UQAuT37HOjhicZFYD4QSg/lGlj3vtUxKSztSC92BSiCBS1Ms/1C7MLaSA4zcfo
I0UQbCV/SYUioizHVCtulsdKiaY0k61e75Iz4DffoV1NQLYV+EHafyAduVpARJAeqauf3YDKgoZ6
ldvBA8IuYED6UzoTiALIkAR+CBaYxq5v1m6iUrcBZHMbvFtG/sDtBpPzFbzaL601/ZAbeHzOGeUN
4v/INQ0SYl8mr0Gkt3mgce9fkPSZZLHTsdkECY3F98yF+rLTjKJlvoqkMlbTfqOnxp3mK4yDTr/1
/YFKvRU5IQA98r3cm5q2LGTlAqB05RlnAcYokMqBFe33zFksBWegLBXWXeIepk4uH/hGrWyuU6Ud
7RMaUj91kHqTEAVarTOWWwIFwK0oeAgvVjjizc52/5tFaSvZhHV6GWARlIIRbmxW7CFvl/rNX05t
qZqnmqOctvchin3OqgBA7c5YDbJhdzitV3bUL3GQnFOuQtIcJfhv+oq6ZruQ2avEhWvJ681fLDq6
yQ==
`protect end_protected
